module tt_um_froith_goldcrest (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire clknet_leaf_0_clk;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire net1980;
 wire _13209_;
 wire _13210_;
 wire \top_ihp.gpio_o_1 ;
 wire \top_ihp.gpio_o_2 ;
 wire \top_ihp.gpio_o_3 ;
 wire \top_ihp.gpio_o_4 ;
 wire \top_ihp.oisc.decoder.decoded[0] ;
 wire \top_ihp.oisc.decoder.decoded[10] ;
 wire \top_ihp.oisc.decoder.decoded[11] ;
 wire \top_ihp.oisc.decoder.decoded[12] ;
 wire \top_ihp.oisc.decoder.decoded[13] ;
 wire \top_ihp.oisc.decoder.decoded[14] ;
 wire \top_ihp.oisc.decoder.decoded[15] ;
 wire \top_ihp.oisc.decoder.decoded[1] ;
 wire \top_ihp.oisc.decoder.decoded[2] ;
 wire \top_ihp.oisc.decoder.decoded[3] ;
 wire \top_ihp.oisc.decoder.decoded[4] ;
 wire \top_ihp.oisc.decoder.decoded[5] ;
 wire \top_ihp.oisc.decoder.decoded[6] ;
 wire \top_ihp.oisc.decoder.decoded[7] ;
 wire \top_ihp.oisc.decoder.instruction[10] ;
 wire \top_ihp.oisc.decoder.instruction[11] ;
 wire \top_ihp.oisc.decoder.instruction[12] ;
 wire \top_ihp.oisc.decoder.instruction[13] ;
 wire \top_ihp.oisc.decoder.instruction[14] ;
 wire \top_ihp.oisc.decoder.instruction[15] ;
 wire \top_ihp.oisc.decoder.instruction[16] ;
 wire \top_ihp.oisc.decoder.instruction[17] ;
 wire \top_ihp.oisc.decoder.instruction[18] ;
 wire \top_ihp.oisc.decoder.instruction[19] ;
 wire \top_ihp.oisc.decoder.instruction[20] ;
 wire \top_ihp.oisc.decoder.instruction[21] ;
 wire \top_ihp.oisc.decoder.instruction[22] ;
 wire \top_ihp.oisc.decoder.instruction[23] ;
 wire \top_ihp.oisc.decoder.instruction[24] ;
 wire \top_ihp.oisc.decoder.instruction[25] ;
 wire \top_ihp.oisc.decoder.instruction[26] ;
 wire \top_ihp.oisc.decoder.instruction[27] ;
 wire \top_ihp.oisc.decoder.instruction[28] ;
 wire \top_ihp.oisc.decoder.instruction[29] ;
 wire \top_ihp.oisc.decoder.instruction[30] ;
 wire \top_ihp.oisc.decoder.instruction[31] ;
 wire \top_ihp.oisc.decoder.instruction[7] ;
 wire \top_ihp.oisc.decoder.instruction[8] ;
 wire \top_ihp.oisc.decoder.instruction[9] ;
 wire \top_ihp.oisc.mem_addr_lowbits[0] ;
 wire \top_ihp.oisc.mem_addr_lowbits[1] ;
 wire \top_ihp.oisc.micro_op[0] ;
 wire \top_ihp.oisc.micro_op[10] ;
 wire \top_ihp.oisc.micro_op[11] ;
 wire \top_ihp.oisc.micro_op[12] ;
 wire \top_ihp.oisc.micro_op[13] ;
 wire \top_ihp.oisc.micro_op[14] ;
 wire \top_ihp.oisc.micro_op[15] ;
 wire \top_ihp.oisc.micro_op[1] ;
 wire \top_ihp.oisc.micro_op[2] ;
 wire \top_ihp.oisc.micro_op[3] ;
 wire \top_ihp.oisc.micro_op[4] ;
 wire \top_ihp.oisc.micro_op[5] ;
 wire \top_ihp.oisc.micro_op[8] ;
 wire \top_ihp.oisc.micro_op[9] ;
 wire \top_ihp.oisc.micro_pc[0] ;
 wire \top_ihp.oisc.micro_pc[1] ;
 wire \top_ihp.oisc.micro_pc[2] ;
 wire \top_ihp.oisc.micro_pc[3] ;
 wire \top_ihp.oisc.micro_pc[4] ;
 wire \top_ihp.oisc.micro_pc[5] ;
 wire \top_ihp.oisc.micro_pc[6] ;
 wire \top_ihp.oisc.micro_pc[7] ;
 wire \top_ihp.oisc.micro_res_addr[0] ;
 wire \top_ihp.oisc.micro_res_addr[1] ;
 wire \top_ihp.oisc.micro_res_addr[2] ;
 wire \top_ihp.oisc.micro_res_addr[3] ;
 wire \top_ihp.oisc.micro_state[0] ;
 wire \top_ihp.oisc.micro_state[1] ;
 wire \top_ihp.oisc.micro_state[2] ;
 wire \top_ihp.oisc.op_a[0] ;
 wire \top_ihp.oisc.op_a[10] ;
 wire \top_ihp.oisc.op_a[11] ;
 wire \top_ihp.oisc.op_a[12] ;
 wire \top_ihp.oisc.op_a[13] ;
 wire \top_ihp.oisc.op_a[14] ;
 wire \top_ihp.oisc.op_a[15] ;
 wire \top_ihp.oisc.op_a[16] ;
 wire \top_ihp.oisc.op_a[17] ;
 wire \top_ihp.oisc.op_a[18] ;
 wire \top_ihp.oisc.op_a[19] ;
 wire \top_ihp.oisc.op_a[1] ;
 wire \top_ihp.oisc.op_a[20] ;
 wire \top_ihp.oisc.op_a[21] ;
 wire \top_ihp.oisc.op_a[22] ;
 wire \top_ihp.oisc.op_a[23] ;
 wire \top_ihp.oisc.op_a[24] ;
 wire \top_ihp.oisc.op_a[25] ;
 wire \top_ihp.oisc.op_a[26] ;
 wire \top_ihp.oisc.op_a[27] ;
 wire \top_ihp.oisc.op_a[28] ;
 wire \top_ihp.oisc.op_a[29] ;
 wire \top_ihp.oisc.op_a[2] ;
 wire \top_ihp.oisc.op_a[30] ;
 wire \top_ihp.oisc.op_a[31] ;
 wire \top_ihp.oisc.op_a[3] ;
 wire \top_ihp.oisc.op_a[4] ;
 wire \top_ihp.oisc.op_a[5] ;
 wire \top_ihp.oisc.op_a[6] ;
 wire \top_ihp.oisc.op_a[7] ;
 wire \top_ihp.oisc.op_a[8] ;
 wire \top_ihp.oisc.op_a[9] ;
 wire \top_ihp.oisc.op_b[0] ;
 wire \top_ihp.oisc.op_b[10] ;
 wire \top_ihp.oisc.op_b[11] ;
 wire \top_ihp.oisc.op_b[12] ;
 wire \top_ihp.oisc.op_b[13] ;
 wire \top_ihp.oisc.op_b[14] ;
 wire \top_ihp.oisc.op_b[15] ;
 wire \top_ihp.oisc.op_b[16] ;
 wire \top_ihp.oisc.op_b[17] ;
 wire \top_ihp.oisc.op_b[18] ;
 wire \top_ihp.oisc.op_b[19] ;
 wire \top_ihp.oisc.op_b[1] ;
 wire \top_ihp.oisc.op_b[20] ;
 wire \top_ihp.oisc.op_b[21] ;
 wire \top_ihp.oisc.op_b[22] ;
 wire \top_ihp.oisc.op_b[23] ;
 wire \top_ihp.oisc.op_b[24] ;
 wire \top_ihp.oisc.op_b[25] ;
 wire \top_ihp.oisc.op_b[26] ;
 wire \top_ihp.oisc.op_b[27] ;
 wire \top_ihp.oisc.op_b[28] ;
 wire \top_ihp.oisc.op_b[29] ;
 wire \top_ihp.oisc.op_b[2] ;
 wire \top_ihp.oisc.op_b[30] ;
 wire \top_ihp.oisc.op_b[31] ;
 wire \top_ihp.oisc.op_b[3] ;
 wire \top_ihp.oisc.op_b[4] ;
 wire \top_ihp.oisc.op_b[5] ;
 wire \top_ihp.oisc.op_b[6] ;
 wire \top_ihp.oisc.op_b[7] ;
 wire \top_ihp.oisc.op_b[8] ;
 wire \top_ihp.oisc.op_b[9] ;
 wire \top_ihp.oisc.reg_rb[0] ;
 wire \top_ihp.oisc.reg_rb[1] ;
 wire \top_ihp.oisc.reg_rb[2] ;
 wire \top_ihp.oisc.reg_rb[3] ;
 wire \top_ihp.oisc.regs[0][0] ;
 wire \top_ihp.oisc.regs[0][10] ;
 wire \top_ihp.oisc.regs[0][11] ;
 wire \top_ihp.oisc.regs[0][12] ;
 wire \top_ihp.oisc.regs[0][13] ;
 wire \top_ihp.oisc.regs[0][14] ;
 wire \top_ihp.oisc.regs[0][15] ;
 wire \top_ihp.oisc.regs[0][16] ;
 wire \top_ihp.oisc.regs[0][17] ;
 wire \top_ihp.oisc.regs[0][18] ;
 wire \top_ihp.oisc.regs[0][19] ;
 wire \top_ihp.oisc.regs[0][1] ;
 wire \top_ihp.oisc.regs[0][20] ;
 wire \top_ihp.oisc.regs[0][21] ;
 wire \top_ihp.oisc.regs[0][22] ;
 wire \top_ihp.oisc.regs[0][23] ;
 wire \top_ihp.oisc.regs[0][24] ;
 wire \top_ihp.oisc.regs[0][25] ;
 wire \top_ihp.oisc.regs[0][26] ;
 wire \top_ihp.oisc.regs[0][27] ;
 wire \top_ihp.oisc.regs[0][28] ;
 wire \top_ihp.oisc.regs[0][29] ;
 wire \top_ihp.oisc.regs[0][2] ;
 wire \top_ihp.oisc.regs[0][30] ;
 wire \top_ihp.oisc.regs[0][31] ;
 wire \top_ihp.oisc.regs[0][3] ;
 wire \top_ihp.oisc.regs[0][4] ;
 wire \top_ihp.oisc.regs[0][5] ;
 wire \top_ihp.oisc.regs[0][6] ;
 wire \top_ihp.oisc.regs[0][7] ;
 wire \top_ihp.oisc.regs[0][8] ;
 wire \top_ihp.oisc.regs[0][9] ;
 wire \top_ihp.oisc.regs[10][0] ;
 wire \top_ihp.oisc.regs[10][10] ;
 wire \top_ihp.oisc.regs[10][11] ;
 wire \top_ihp.oisc.regs[10][12] ;
 wire \top_ihp.oisc.regs[10][13] ;
 wire \top_ihp.oisc.regs[10][14] ;
 wire \top_ihp.oisc.regs[10][15] ;
 wire \top_ihp.oisc.regs[10][16] ;
 wire \top_ihp.oisc.regs[10][17] ;
 wire \top_ihp.oisc.regs[10][18] ;
 wire \top_ihp.oisc.regs[10][19] ;
 wire \top_ihp.oisc.regs[10][1] ;
 wire \top_ihp.oisc.regs[10][20] ;
 wire \top_ihp.oisc.regs[10][21] ;
 wire \top_ihp.oisc.regs[10][22] ;
 wire \top_ihp.oisc.regs[10][23] ;
 wire \top_ihp.oisc.regs[10][24] ;
 wire \top_ihp.oisc.regs[10][25] ;
 wire \top_ihp.oisc.regs[10][26] ;
 wire \top_ihp.oisc.regs[10][27] ;
 wire \top_ihp.oisc.regs[10][28] ;
 wire \top_ihp.oisc.regs[10][29] ;
 wire \top_ihp.oisc.regs[10][2] ;
 wire \top_ihp.oisc.regs[10][30] ;
 wire \top_ihp.oisc.regs[10][31] ;
 wire \top_ihp.oisc.regs[10][3] ;
 wire \top_ihp.oisc.regs[10][4] ;
 wire \top_ihp.oisc.regs[10][5] ;
 wire \top_ihp.oisc.regs[10][6] ;
 wire \top_ihp.oisc.regs[10][7] ;
 wire \top_ihp.oisc.regs[10][8] ;
 wire \top_ihp.oisc.regs[10][9] ;
 wire \top_ihp.oisc.regs[11][0] ;
 wire \top_ihp.oisc.regs[11][10] ;
 wire \top_ihp.oisc.regs[11][11] ;
 wire \top_ihp.oisc.regs[11][12] ;
 wire \top_ihp.oisc.regs[11][13] ;
 wire \top_ihp.oisc.regs[11][14] ;
 wire \top_ihp.oisc.regs[11][15] ;
 wire \top_ihp.oisc.regs[11][16] ;
 wire \top_ihp.oisc.regs[11][17] ;
 wire \top_ihp.oisc.regs[11][18] ;
 wire \top_ihp.oisc.regs[11][19] ;
 wire \top_ihp.oisc.regs[11][1] ;
 wire \top_ihp.oisc.regs[11][20] ;
 wire \top_ihp.oisc.regs[11][21] ;
 wire \top_ihp.oisc.regs[11][22] ;
 wire \top_ihp.oisc.regs[11][23] ;
 wire \top_ihp.oisc.regs[11][24] ;
 wire \top_ihp.oisc.regs[11][25] ;
 wire \top_ihp.oisc.regs[11][26] ;
 wire \top_ihp.oisc.regs[11][27] ;
 wire \top_ihp.oisc.regs[11][28] ;
 wire \top_ihp.oisc.regs[11][29] ;
 wire \top_ihp.oisc.regs[11][2] ;
 wire \top_ihp.oisc.regs[11][30] ;
 wire \top_ihp.oisc.regs[11][31] ;
 wire \top_ihp.oisc.regs[11][3] ;
 wire \top_ihp.oisc.regs[11][4] ;
 wire \top_ihp.oisc.regs[11][5] ;
 wire \top_ihp.oisc.regs[11][6] ;
 wire \top_ihp.oisc.regs[11][7] ;
 wire \top_ihp.oisc.regs[11][8] ;
 wire \top_ihp.oisc.regs[11][9] ;
 wire \top_ihp.oisc.regs[12][0] ;
 wire \top_ihp.oisc.regs[12][10] ;
 wire \top_ihp.oisc.regs[12][11] ;
 wire \top_ihp.oisc.regs[12][12] ;
 wire \top_ihp.oisc.regs[12][13] ;
 wire \top_ihp.oisc.regs[12][14] ;
 wire \top_ihp.oisc.regs[12][15] ;
 wire \top_ihp.oisc.regs[12][16] ;
 wire \top_ihp.oisc.regs[12][17] ;
 wire \top_ihp.oisc.regs[12][18] ;
 wire \top_ihp.oisc.regs[12][19] ;
 wire \top_ihp.oisc.regs[12][1] ;
 wire \top_ihp.oisc.regs[12][20] ;
 wire \top_ihp.oisc.regs[12][21] ;
 wire \top_ihp.oisc.regs[12][22] ;
 wire \top_ihp.oisc.regs[12][23] ;
 wire \top_ihp.oisc.regs[12][24] ;
 wire \top_ihp.oisc.regs[12][25] ;
 wire \top_ihp.oisc.regs[12][26] ;
 wire \top_ihp.oisc.regs[12][27] ;
 wire \top_ihp.oisc.regs[12][28] ;
 wire \top_ihp.oisc.regs[12][29] ;
 wire \top_ihp.oisc.regs[12][2] ;
 wire \top_ihp.oisc.regs[12][30] ;
 wire \top_ihp.oisc.regs[12][31] ;
 wire \top_ihp.oisc.regs[12][3] ;
 wire \top_ihp.oisc.regs[12][4] ;
 wire \top_ihp.oisc.regs[12][5] ;
 wire \top_ihp.oisc.regs[12][6] ;
 wire \top_ihp.oisc.regs[12][7] ;
 wire \top_ihp.oisc.regs[12][8] ;
 wire \top_ihp.oisc.regs[12][9] ;
 wire \top_ihp.oisc.regs[13][0] ;
 wire \top_ihp.oisc.regs[13][10] ;
 wire \top_ihp.oisc.regs[13][11] ;
 wire \top_ihp.oisc.regs[13][12] ;
 wire \top_ihp.oisc.regs[13][13] ;
 wire \top_ihp.oisc.regs[13][14] ;
 wire \top_ihp.oisc.regs[13][15] ;
 wire \top_ihp.oisc.regs[13][16] ;
 wire \top_ihp.oisc.regs[13][17] ;
 wire \top_ihp.oisc.regs[13][18] ;
 wire \top_ihp.oisc.regs[13][19] ;
 wire \top_ihp.oisc.regs[13][1] ;
 wire \top_ihp.oisc.regs[13][20] ;
 wire \top_ihp.oisc.regs[13][21] ;
 wire \top_ihp.oisc.regs[13][22] ;
 wire \top_ihp.oisc.regs[13][23] ;
 wire \top_ihp.oisc.regs[13][24] ;
 wire \top_ihp.oisc.regs[13][25] ;
 wire \top_ihp.oisc.regs[13][26] ;
 wire \top_ihp.oisc.regs[13][27] ;
 wire \top_ihp.oisc.regs[13][28] ;
 wire \top_ihp.oisc.regs[13][29] ;
 wire \top_ihp.oisc.regs[13][2] ;
 wire \top_ihp.oisc.regs[13][30] ;
 wire \top_ihp.oisc.regs[13][31] ;
 wire \top_ihp.oisc.regs[13][3] ;
 wire \top_ihp.oisc.regs[13][4] ;
 wire \top_ihp.oisc.regs[13][5] ;
 wire \top_ihp.oisc.regs[13][6] ;
 wire \top_ihp.oisc.regs[13][7] ;
 wire \top_ihp.oisc.regs[13][8] ;
 wire \top_ihp.oisc.regs[13][9] ;
 wire \top_ihp.oisc.regs[14][0] ;
 wire \top_ihp.oisc.regs[14][10] ;
 wire \top_ihp.oisc.regs[14][11] ;
 wire \top_ihp.oisc.regs[14][12] ;
 wire \top_ihp.oisc.regs[14][13] ;
 wire \top_ihp.oisc.regs[14][14] ;
 wire \top_ihp.oisc.regs[14][15] ;
 wire \top_ihp.oisc.regs[14][16] ;
 wire \top_ihp.oisc.regs[14][17] ;
 wire \top_ihp.oisc.regs[14][18] ;
 wire \top_ihp.oisc.regs[14][19] ;
 wire \top_ihp.oisc.regs[14][1] ;
 wire \top_ihp.oisc.regs[14][20] ;
 wire \top_ihp.oisc.regs[14][21] ;
 wire \top_ihp.oisc.regs[14][22] ;
 wire \top_ihp.oisc.regs[14][23] ;
 wire \top_ihp.oisc.regs[14][24] ;
 wire \top_ihp.oisc.regs[14][25] ;
 wire \top_ihp.oisc.regs[14][26] ;
 wire \top_ihp.oisc.regs[14][27] ;
 wire \top_ihp.oisc.regs[14][28] ;
 wire \top_ihp.oisc.regs[14][29] ;
 wire \top_ihp.oisc.regs[14][2] ;
 wire \top_ihp.oisc.regs[14][30] ;
 wire \top_ihp.oisc.regs[14][31] ;
 wire \top_ihp.oisc.regs[14][3] ;
 wire \top_ihp.oisc.regs[14][4] ;
 wire \top_ihp.oisc.regs[14][5] ;
 wire \top_ihp.oisc.regs[14][6] ;
 wire \top_ihp.oisc.regs[14][7] ;
 wire \top_ihp.oisc.regs[14][8] ;
 wire \top_ihp.oisc.regs[14][9] ;
 wire \top_ihp.oisc.regs[15][0] ;
 wire \top_ihp.oisc.regs[15][10] ;
 wire \top_ihp.oisc.regs[15][11] ;
 wire \top_ihp.oisc.regs[15][12] ;
 wire \top_ihp.oisc.regs[15][13] ;
 wire \top_ihp.oisc.regs[15][14] ;
 wire \top_ihp.oisc.regs[15][15] ;
 wire \top_ihp.oisc.regs[15][16] ;
 wire \top_ihp.oisc.regs[15][17] ;
 wire \top_ihp.oisc.regs[15][18] ;
 wire \top_ihp.oisc.regs[15][19] ;
 wire \top_ihp.oisc.regs[15][1] ;
 wire \top_ihp.oisc.regs[15][20] ;
 wire \top_ihp.oisc.regs[15][21] ;
 wire \top_ihp.oisc.regs[15][22] ;
 wire \top_ihp.oisc.regs[15][23] ;
 wire \top_ihp.oisc.regs[15][24] ;
 wire \top_ihp.oisc.regs[15][25] ;
 wire \top_ihp.oisc.regs[15][26] ;
 wire \top_ihp.oisc.regs[15][27] ;
 wire \top_ihp.oisc.regs[15][28] ;
 wire \top_ihp.oisc.regs[15][29] ;
 wire \top_ihp.oisc.regs[15][2] ;
 wire \top_ihp.oisc.regs[15][30] ;
 wire \top_ihp.oisc.regs[15][31] ;
 wire \top_ihp.oisc.regs[15][3] ;
 wire \top_ihp.oisc.regs[15][4] ;
 wire \top_ihp.oisc.regs[15][5] ;
 wire \top_ihp.oisc.regs[15][6] ;
 wire \top_ihp.oisc.regs[15][7] ;
 wire \top_ihp.oisc.regs[15][8] ;
 wire \top_ihp.oisc.regs[15][9] ;
 wire \top_ihp.oisc.regs[16][0] ;
 wire \top_ihp.oisc.regs[16][10] ;
 wire \top_ihp.oisc.regs[16][11] ;
 wire \top_ihp.oisc.regs[16][12] ;
 wire \top_ihp.oisc.regs[16][13] ;
 wire \top_ihp.oisc.regs[16][14] ;
 wire \top_ihp.oisc.regs[16][15] ;
 wire \top_ihp.oisc.regs[16][16] ;
 wire \top_ihp.oisc.regs[16][17] ;
 wire \top_ihp.oisc.regs[16][18] ;
 wire \top_ihp.oisc.regs[16][19] ;
 wire \top_ihp.oisc.regs[16][1] ;
 wire \top_ihp.oisc.regs[16][20] ;
 wire \top_ihp.oisc.regs[16][21] ;
 wire \top_ihp.oisc.regs[16][22] ;
 wire \top_ihp.oisc.regs[16][23] ;
 wire \top_ihp.oisc.regs[16][24] ;
 wire \top_ihp.oisc.regs[16][25] ;
 wire \top_ihp.oisc.regs[16][26] ;
 wire \top_ihp.oisc.regs[16][27] ;
 wire \top_ihp.oisc.regs[16][28] ;
 wire \top_ihp.oisc.regs[16][29] ;
 wire \top_ihp.oisc.regs[16][2] ;
 wire \top_ihp.oisc.regs[16][30] ;
 wire \top_ihp.oisc.regs[16][31] ;
 wire \top_ihp.oisc.regs[16][3] ;
 wire \top_ihp.oisc.regs[16][4] ;
 wire \top_ihp.oisc.regs[16][5] ;
 wire \top_ihp.oisc.regs[16][6] ;
 wire \top_ihp.oisc.regs[16][7] ;
 wire \top_ihp.oisc.regs[16][8] ;
 wire \top_ihp.oisc.regs[16][9] ;
 wire \top_ihp.oisc.regs[17][0] ;
 wire \top_ihp.oisc.regs[17][10] ;
 wire \top_ihp.oisc.regs[17][11] ;
 wire \top_ihp.oisc.regs[17][12] ;
 wire \top_ihp.oisc.regs[17][13] ;
 wire \top_ihp.oisc.regs[17][14] ;
 wire \top_ihp.oisc.regs[17][15] ;
 wire \top_ihp.oisc.regs[17][16] ;
 wire \top_ihp.oisc.regs[17][17] ;
 wire \top_ihp.oisc.regs[17][18] ;
 wire \top_ihp.oisc.regs[17][19] ;
 wire \top_ihp.oisc.regs[17][1] ;
 wire \top_ihp.oisc.regs[17][20] ;
 wire \top_ihp.oisc.regs[17][21] ;
 wire \top_ihp.oisc.regs[17][22] ;
 wire \top_ihp.oisc.regs[17][23] ;
 wire \top_ihp.oisc.regs[17][24] ;
 wire \top_ihp.oisc.regs[17][25] ;
 wire \top_ihp.oisc.regs[17][26] ;
 wire \top_ihp.oisc.regs[17][27] ;
 wire \top_ihp.oisc.regs[17][28] ;
 wire \top_ihp.oisc.regs[17][29] ;
 wire \top_ihp.oisc.regs[17][2] ;
 wire \top_ihp.oisc.regs[17][30] ;
 wire \top_ihp.oisc.regs[17][31] ;
 wire \top_ihp.oisc.regs[17][3] ;
 wire \top_ihp.oisc.regs[17][4] ;
 wire \top_ihp.oisc.regs[17][5] ;
 wire \top_ihp.oisc.regs[17][6] ;
 wire \top_ihp.oisc.regs[17][7] ;
 wire \top_ihp.oisc.regs[17][8] ;
 wire \top_ihp.oisc.regs[17][9] ;
 wire \top_ihp.oisc.regs[18][0] ;
 wire \top_ihp.oisc.regs[18][10] ;
 wire \top_ihp.oisc.regs[18][11] ;
 wire \top_ihp.oisc.regs[18][12] ;
 wire \top_ihp.oisc.regs[18][13] ;
 wire \top_ihp.oisc.regs[18][14] ;
 wire \top_ihp.oisc.regs[18][15] ;
 wire \top_ihp.oisc.regs[18][16] ;
 wire \top_ihp.oisc.regs[18][17] ;
 wire \top_ihp.oisc.regs[18][18] ;
 wire \top_ihp.oisc.regs[18][19] ;
 wire \top_ihp.oisc.regs[18][1] ;
 wire \top_ihp.oisc.regs[18][20] ;
 wire \top_ihp.oisc.regs[18][21] ;
 wire \top_ihp.oisc.regs[18][22] ;
 wire \top_ihp.oisc.regs[18][23] ;
 wire \top_ihp.oisc.regs[18][24] ;
 wire \top_ihp.oisc.regs[18][25] ;
 wire \top_ihp.oisc.regs[18][26] ;
 wire \top_ihp.oisc.regs[18][27] ;
 wire \top_ihp.oisc.regs[18][28] ;
 wire \top_ihp.oisc.regs[18][29] ;
 wire \top_ihp.oisc.regs[18][2] ;
 wire \top_ihp.oisc.regs[18][30] ;
 wire \top_ihp.oisc.regs[18][31] ;
 wire \top_ihp.oisc.regs[18][3] ;
 wire \top_ihp.oisc.regs[18][4] ;
 wire \top_ihp.oisc.regs[18][5] ;
 wire \top_ihp.oisc.regs[18][6] ;
 wire \top_ihp.oisc.regs[18][7] ;
 wire \top_ihp.oisc.regs[18][8] ;
 wire \top_ihp.oisc.regs[18][9] ;
 wire \top_ihp.oisc.regs[19][0] ;
 wire \top_ihp.oisc.regs[19][10] ;
 wire \top_ihp.oisc.regs[19][11] ;
 wire \top_ihp.oisc.regs[19][12] ;
 wire \top_ihp.oisc.regs[19][13] ;
 wire \top_ihp.oisc.regs[19][14] ;
 wire \top_ihp.oisc.regs[19][15] ;
 wire \top_ihp.oisc.regs[19][16] ;
 wire \top_ihp.oisc.regs[19][17] ;
 wire \top_ihp.oisc.regs[19][18] ;
 wire \top_ihp.oisc.regs[19][19] ;
 wire \top_ihp.oisc.regs[19][1] ;
 wire \top_ihp.oisc.regs[19][20] ;
 wire \top_ihp.oisc.regs[19][21] ;
 wire \top_ihp.oisc.regs[19][22] ;
 wire \top_ihp.oisc.regs[19][23] ;
 wire \top_ihp.oisc.regs[19][24] ;
 wire \top_ihp.oisc.regs[19][25] ;
 wire \top_ihp.oisc.regs[19][26] ;
 wire \top_ihp.oisc.regs[19][27] ;
 wire \top_ihp.oisc.regs[19][28] ;
 wire \top_ihp.oisc.regs[19][29] ;
 wire \top_ihp.oisc.regs[19][2] ;
 wire \top_ihp.oisc.regs[19][30] ;
 wire \top_ihp.oisc.regs[19][31] ;
 wire \top_ihp.oisc.regs[19][3] ;
 wire \top_ihp.oisc.regs[19][4] ;
 wire \top_ihp.oisc.regs[19][5] ;
 wire \top_ihp.oisc.regs[19][6] ;
 wire \top_ihp.oisc.regs[19][7] ;
 wire \top_ihp.oisc.regs[19][8] ;
 wire \top_ihp.oisc.regs[19][9] ;
 wire \top_ihp.oisc.regs[1][0] ;
 wire \top_ihp.oisc.regs[1][10] ;
 wire \top_ihp.oisc.regs[1][11] ;
 wire \top_ihp.oisc.regs[1][12] ;
 wire \top_ihp.oisc.regs[1][13] ;
 wire \top_ihp.oisc.regs[1][14] ;
 wire \top_ihp.oisc.regs[1][15] ;
 wire \top_ihp.oisc.regs[1][16] ;
 wire \top_ihp.oisc.regs[1][17] ;
 wire \top_ihp.oisc.regs[1][18] ;
 wire \top_ihp.oisc.regs[1][19] ;
 wire \top_ihp.oisc.regs[1][1] ;
 wire \top_ihp.oisc.regs[1][20] ;
 wire \top_ihp.oisc.regs[1][21] ;
 wire \top_ihp.oisc.regs[1][22] ;
 wire \top_ihp.oisc.regs[1][23] ;
 wire \top_ihp.oisc.regs[1][24] ;
 wire \top_ihp.oisc.regs[1][25] ;
 wire \top_ihp.oisc.regs[1][26] ;
 wire \top_ihp.oisc.regs[1][27] ;
 wire \top_ihp.oisc.regs[1][28] ;
 wire \top_ihp.oisc.regs[1][29] ;
 wire \top_ihp.oisc.regs[1][2] ;
 wire \top_ihp.oisc.regs[1][30] ;
 wire \top_ihp.oisc.regs[1][31] ;
 wire \top_ihp.oisc.regs[1][3] ;
 wire \top_ihp.oisc.regs[1][4] ;
 wire \top_ihp.oisc.regs[1][5] ;
 wire \top_ihp.oisc.regs[1][6] ;
 wire \top_ihp.oisc.regs[1][7] ;
 wire \top_ihp.oisc.regs[1][8] ;
 wire \top_ihp.oisc.regs[1][9] ;
 wire \top_ihp.oisc.regs[20][0] ;
 wire \top_ihp.oisc.regs[20][10] ;
 wire \top_ihp.oisc.regs[20][11] ;
 wire \top_ihp.oisc.regs[20][12] ;
 wire \top_ihp.oisc.regs[20][13] ;
 wire \top_ihp.oisc.regs[20][14] ;
 wire \top_ihp.oisc.regs[20][15] ;
 wire \top_ihp.oisc.regs[20][16] ;
 wire \top_ihp.oisc.regs[20][17] ;
 wire \top_ihp.oisc.regs[20][18] ;
 wire \top_ihp.oisc.regs[20][19] ;
 wire \top_ihp.oisc.regs[20][1] ;
 wire \top_ihp.oisc.regs[20][20] ;
 wire \top_ihp.oisc.regs[20][21] ;
 wire \top_ihp.oisc.regs[20][22] ;
 wire \top_ihp.oisc.regs[20][23] ;
 wire \top_ihp.oisc.regs[20][24] ;
 wire \top_ihp.oisc.regs[20][25] ;
 wire \top_ihp.oisc.regs[20][26] ;
 wire \top_ihp.oisc.regs[20][27] ;
 wire \top_ihp.oisc.regs[20][28] ;
 wire \top_ihp.oisc.regs[20][29] ;
 wire \top_ihp.oisc.regs[20][2] ;
 wire \top_ihp.oisc.regs[20][30] ;
 wire \top_ihp.oisc.regs[20][31] ;
 wire \top_ihp.oisc.regs[20][3] ;
 wire \top_ihp.oisc.regs[20][4] ;
 wire \top_ihp.oisc.regs[20][5] ;
 wire \top_ihp.oisc.regs[20][6] ;
 wire \top_ihp.oisc.regs[20][7] ;
 wire \top_ihp.oisc.regs[20][8] ;
 wire \top_ihp.oisc.regs[20][9] ;
 wire \top_ihp.oisc.regs[21][0] ;
 wire \top_ihp.oisc.regs[21][10] ;
 wire \top_ihp.oisc.regs[21][11] ;
 wire \top_ihp.oisc.regs[21][12] ;
 wire \top_ihp.oisc.regs[21][13] ;
 wire \top_ihp.oisc.regs[21][14] ;
 wire \top_ihp.oisc.regs[21][15] ;
 wire \top_ihp.oisc.regs[21][16] ;
 wire \top_ihp.oisc.regs[21][17] ;
 wire \top_ihp.oisc.regs[21][18] ;
 wire \top_ihp.oisc.regs[21][19] ;
 wire \top_ihp.oisc.regs[21][1] ;
 wire \top_ihp.oisc.regs[21][20] ;
 wire \top_ihp.oisc.regs[21][21] ;
 wire \top_ihp.oisc.regs[21][22] ;
 wire \top_ihp.oisc.regs[21][23] ;
 wire \top_ihp.oisc.regs[21][24] ;
 wire \top_ihp.oisc.regs[21][25] ;
 wire \top_ihp.oisc.regs[21][26] ;
 wire \top_ihp.oisc.regs[21][27] ;
 wire \top_ihp.oisc.regs[21][28] ;
 wire \top_ihp.oisc.regs[21][29] ;
 wire \top_ihp.oisc.regs[21][2] ;
 wire \top_ihp.oisc.regs[21][30] ;
 wire \top_ihp.oisc.regs[21][31] ;
 wire \top_ihp.oisc.regs[21][3] ;
 wire \top_ihp.oisc.regs[21][4] ;
 wire \top_ihp.oisc.regs[21][5] ;
 wire \top_ihp.oisc.regs[21][6] ;
 wire \top_ihp.oisc.regs[21][7] ;
 wire \top_ihp.oisc.regs[21][8] ;
 wire \top_ihp.oisc.regs[21][9] ;
 wire \top_ihp.oisc.regs[22][0] ;
 wire \top_ihp.oisc.regs[22][10] ;
 wire \top_ihp.oisc.regs[22][11] ;
 wire \top_ihp.oisc.regs[22][12] ;
 wire \top_ihp.oisc.regs[22][13] ;
 wire \top_ihp.oisc.regs[22][14] ;
 wire \top_ihp.oisc.regs[22][15] ;
 wire \top_ihp.oisc.regs[22][16] ;
 wire \top_ihp.oisc.regs[22][17] ;
 wire \top_ihp.oisc.regs[22][18] ;
 wire \top_ihp.oisc.regs[22][19] ;
 wire \top_ihp.oisc.regs[22][1] ;
 wire \top_ihp.oisc.regs[22][20] ;
 wire \top_ihp.oisc.regs[22][21] ;
 wire \top_ihp.oisc.regs[22][22] ;
 wire \top_ihp.oisc.regs[22][23] ;
 wire \top_ihp.oisc.regs[22][24] ;
 wire \top_ihp.oisc.regs[22][25] ;
 wire \top_ihp.oisc.regs[22][26] ;
 wire \top_ihp.oisc.regs[22][27] ;
 wire \top_ihp.oisc.regs[22][28] ;
 wire \top_ihp.oisc.regs[22][29] ;
 wire \top_ihp.oisc.regs[22][2] ;
 wire \top_ihp.oisc.regs[22][30] ;
 wire \top_ihp.oisc.regs[22][31] ;
 wire \top_ihp.oisc.regs[22][3] ;
 wire \top_ihp.oisc.regs[22][4] ;
 wire \top_ihp.oisc.regs[22][5] ;
 wire \top_ihp.oisc.regs[22][6] ;
 wire \top_ihp.oisc.regs[22][7] ;
 wire \top_ihp.oisc.regs[22][8] ;
 wire \top_ihp.oisc.regs[22][9] ;
 wire \top_ihp.oisc.regs[23][0] ;
 wire \top_ihp.oisc.regs[23][10] ;
 wire \top_ihp.oisc.regs[23][11] ;
 wire \top_ihp.oisc.regs[23][12] ;
 wire \top_ihp.oisc.regs[23][13] ;
 wire \top_ihp.oisc.regs[23][14] ;
 wire \top_ihp.oisc.regs[23][15] ;
 wire \top_ihp.oisc.regs[23][16] ;
 wire \top_ihp.oisc.regs[23][17] ;
 wire \top_ihp.oisc.regs[23][18] ;
 wire \top_ihp.oisc.regs[23][19] ;
 wire \top_ihp.oisc.regs[23][1] ;
 wire \top_ihp.oisc.regs[23][20] ;
 wire \top_ihp.oisc.regs[23][21] ;
 wire \top_ihp.oisc.regs[23][22] ;
 wire \top_ihp.oisc.regs[23][23] ;
 wire \top_ihp.oisc.regs[23][24] ;
 wire \top_ihp.oisc.regs[23][25] ;
 wire \top_ihp.oisc.regs[23][26] ;
 wire \top_ihp.oisc.regs[23][27] ;
 wire \top_ihp.oisc.regs[23][28] ;
 wire \top_ihp.oisc.regs[23][29] ;
 wire \top_ihp.oisc.regs[23][2] ;
 wire \top_ihp.oisc.regs[23][30] ;
 wire \top_ihp.oisc.regs[23][31] ;
 wire \top_ihp.oisc.regs[23][3] ;
 wire \top_ihp.oisc.regs[23][4] ;
 wire \top_ihp.oisc.regs[23][5] ;
 wire \top_ihp.oisc.regs[23][6] ;
 wire \top_ihp.oisc.regs[23][7] ;
 wire \top_ihp.oisc.regs[23][8] ;
 wire \top_ihp.oisc.regs[23][9] ;
 wire \top_ihp.oisc.regs[24][0] ;
 wire \top_ihp.oisc.regs[24][10] ;
 wire \top_ihp.oisc.regs[24][11] ;
 wire \top_ihp.oisc.regs[24][12] ;
 wire \top_ihp.oisc.regs[24][13] ;
 wire \top_ihp.oisc.regs[24][14] ;
 wire \top_ihp.oisc.regs[24][15] ;
 wire \top_ihp.oisc.regs[24][16] ;
 wire \top_ihp.oisc.regs[24][17] ;
 wire \top_ihp.oisc.regs[24][18] ;
 wire \top_ihp.oisc.regs[24][19] ;
 wire \top_ihp.oisc.regs[24][1] ;
 wire \top_ihp.oisc.regs[24][20] ;
 wire \top_ihp.oisc.regs[24][21] ;
 wire \top_ihp.oisc.regs[24][22] ;
 wire \top_ihp.oisc.regs[24][23] ;
 wire \top_ihp.oisc.regs[24][24] ;
 wire \top_ihp.oisc.regs[24][25] ;
 wire \top_ihp.oisc.regs[24][26] ;
 wire \top_ihp.oisc.regs[24][27] ;
 wire \top_ihp.oisc.regs[24][28] ;
 wire \top_ihp.oisc.regs[24][29] ;
 wire \top_ihp.oisc.regs[24][2] ;
 wire \top_ihp.oisc.regs[24][30] ;
 wire \top_ihp.oisc.regs[24][31] ;
 wire \top_ihp.oisc.regs[24][3] ;
 wire \top_ihp.oisc.regs[24][4] ;
 wire \top_ihp.oisc.regs[24][5] ;
 wire \top_ihp.oisc.regs[24][6] ;
 wire \top_ihp.oisc.regs[24][7] ;
 wire \top_ihp.oisc.regs[24][8] ;
 wire \top_ihp.oisc.regs[24][9] ;
 wire \top_ihp.oisc.regs[25][0] ;
 wire \top_ihp.oisc.regs[25][10] ;
 wire \top_ihp.oisc.regs[25][11] ;
 wire \top_ihp.oisc.regs[25][12] ;
 wire \top_ihp.oisc.regs[25][13] ;
 wire \top_ihp.oisc.regs[25][14] ;
 wire \top_ihp.oisc.regs[25][15] ;
 wire \top_ihp.oisc.regs[25][16] ;
 wire \top_ihp.oisc.regs[25][17] ;
 wire \top_ihp.oisc.regs[25][18] ;
 wire \top_ihp.oisc.regs[25][19] ;
 wire \top_ihp.oisc.regs[25][1] ;
 wire \top_ihp.oisc.regs[25][20] ;
 wire \top_ihp.oisc.regs[25][21] ;
 wire \top_ihp.oisc.regs[25][22] ;
 wire \top_ihp.oisc.regs[25][23] ;
 wire \top_ihp.oisc.regs[25][24] ;
 wire \top_ihp.oisc.regs[25][25] ;
 wire \top_ihp.oisc.regs[25][26] ;
 wire \top_ihp.oisc.regs[25][27] ;
 wire \top_ihp.oisc.regs[25][28] ;
 wire \top_ihp.oisc.regs[25][29] ;
 wire \top_ihp.oisc.regs[25][2] ;
 wire \top_ihp.oisc.regs[25][30] ;
 wire \top_ihp.oisc.regs[25][31] ;
 wire \top_ihp.oisc.regs[25][3] ;
 wire \top_ihp.oisc.regs[25][4] ;
 wire \top_ihp.oisc.regs[25][5] ;
 wire \top_ihp.oisc.regs[25][6] ;
 wire \top_ihp.oisc.regs[25][7] ;
 wire \top_ihp.oisc.regs[25][8] ;
 wire \top_ihp.oisc.regs[25][9] ;
 wire \top_ihp.oisc.regs[26][0] ;
 wire \top_ihp.oisc.regs[26][10] ;
 wire \top_ihp.oisc.regs[26][11] ;
 wire \top_ihp.oisc.regs[26][12] ;
 wire \top_ihp.oisc.regs[26][13] ;
 wire \top_ihp.oisc.regs[26][14] ;
 wire \top_ihp.oisc.regs[26][15] ;
 wire \top_ihp.oisc.regs[26][16] ;
 wire \top_ihp.oisc.regs[26][17] ;
 wire \top_ihp.oisc.regs[26][18] ;
 wire \top_ihp.oisc.regs[26][19] ;
 wire \top_ihp.oisc.regs[26][1] ;
 wire \top_ihp.oisc.regs[26][20] ;
 wire \top_ihp.oisc.regs[26][21] ;
 wire \top_ihp.oisc.regs[26][22] ;
 wire \top_ihp.oisc.regs[26][23] ;
 wire \top_ihp.oisc.regs[26][24] ;
 wire \top_ihp.oisc.regs[26][25] ;
 wire \top_ihp.oisc.regs[26][26] ;
 wire \top_ihp.oisc.regs[26][27] ;
 wire \top_ihp.oisc.regs[26][28] ;
 wire \top_ihp.oisc.regs[26][29] ;
 wire \top_ihp.oisc.regs[26][2] ;
 wire \top_ihp.oisc.regs[26][30] ;
 wire \top_ihp.oisc.regs[26][31] ;
 wire \top_ihp.oisc.regs[26][3] ;
 wire \top_ihp.oisc.regs[26][4] ;
 wire \top_ihp.oisc.regs[26][5] ;
 wire \top_ihp.oisc.regs[26][6] ;
 wire \top_ihp.oisc.regs[26][7] ;
 wire \top_ihp.oisc.regs[26][8] ;
 wire \top_ihp.oisc.regs[26][9] ;
 wire \top_ihp.oisc.regs[27][0] ;
 wire \top_ihp.oisc.regs[27][10] ;
 wire \top_ihp.oisc.regs[27][11] ;
 wire \top_ihp.oisc.regs[27][12] ;
 wire \top_ihp.oisc.regs[27][13] ;
 wire \top_ihp.oisc.regs[27][14] ;
 wire \top_ihp.oisc.regs[27][15] ;
 wire \top_ihp.oisc.regs[27][16] ;
 wire \top_ihp.oisc.regs[27][17] ;
 wire \top_ihp.oisc.regs[27][18] ;
 wire \top_ihp.oisc.regs[27][19] ;
 wire \top_ihp.oisc.regs[27][1] ;
 wire \top_ihp.oisc.regs[27][20] ;
 wire \top_ihp.oisc.regs[27][21] ;
 wire \top_ihp.oisc.regs[27][22] ;
 wire \top_ihp.oisc.regs[27][23] ;
 wire \top_ihp.oisc.regs[27][24] ;
 wire \top_ihp.oisc.regs[27][25] ;
 wire \top_ihp.oisc.regs[27][26] ;
 wire \top_ihp.oisc.regs[27][27] ;
 wire \top_ihp.oisc.regs[27][28] ;
 wire \top_ihp.oisc.regs[27][29] ;
 wire \top_ihp.oisc.regs[27][2] ;
 wire \top_ihp.oisc.regs[27][30] ;
 wire \top_ihp.oisc.regs[27][31] ;
 wire \top_ihp.oisc.regs[27][3] ;
 wire \top_ihp.oisc.regs[27][4] ;
 wire \top_ihp.oisc.regs[27][5] ;
 wire \top_ihp.oisc.regs[27][6] ;
 wire \top_ihp.oisc.regs[27][7] ;
 wire \top_ihp.oisc.regs[27][8] ;
 wire \top_ihp.oisc.regs[27][9] ;
 wire \top_ihp.oisc.regs[28][0] ;
 wire \top_ihp.oisc.regs[28][10] ;
 wire \top_ihp.oisc.regs[28][11] ;
 wire \top_ihp.oisc.regs[28][12] ;
 wire \top_ihp.oisc.regs[28][13] ;
 wire \top_ihp.oisc.regs[28][14] ;
 wire \top_ihp.oisc.regs[28][15] ;
 wire \top_ihp.oisc.regs[28][16] ;
 wire \top_ihp.oisc.regs[28][17] ;
 wire \top_ihp.oisc.regs[28][18] ;
 wire \top_ihp.oisc.regs[28][19] ;
 wire \top_ihp.oisc.regs[28][1] ;
 wire \top_ihp.oisc.regs[28][20] ;
 wire \top_ihp.oisc.regs[28][21] ;
 wire \top_ihp.oisc.regs[28][22] ;
 wire \top_ihp.oisc.regs[28][23] ;
 wire \top_ihp.oisc.regs[28][24] ;
 wire \top_ihp.oisc.regs[28][25] ;
 wire \top_ihp.oisc.regs[28][26] ;
 wire \top_ihp.oisc.regs[28][27] ;
 wire \top_ihp.oisc.regs[28][28] ;
 wire \top_ihp.oisc.regs[28][29] ;
 wire \top_ihp.oisc.regs[28][2] ;
 wire \top_ihp.oisc.regs[28][30] ;
 wire \top_ihp.oisc.regs[28][31] ;
 wire \top_ihp.oisc.regs[28][3] ;
 wire \top_ihp.oisc.regs[28][4] ;
 wire \top_ihp.oisc.regs[28][5] ;
 wire \top_ihp.oisc.regs[28][6] ;
 wire \top_ihp.oisc.regs[28][7] ;
 wire \top_ihp.oisc.regs[28][8] ;
 wire \top_ihp.oisc.regs[28][9] ;
 wire \top_ihp.oisc.regs[29][0] ;
 wire \top_ihp.oisc.regs[29][10] ;
 wire \top_ihp.oisc.regs[29][11] ;
 wire \top_ihp.oisc.regs[29][12] ;
 wire \top_ihp.oisc.regs[29][13] ;
 wire \top_ihp.oisc.regs[29][14] ;
 wire \top_ihp.oisc.regs[29][15] ;
 wire \top_ihp.oisc.regs[29][16] ;
 wire \top_ihp.oisc.regs[29][17] ;
 wire \top_ihp.oisc.regs[29][18] ;
 wire \top_ihp.oisc.regs[29][19] ;
 wire \top_ihp.oisc.regs[29][1] ;
 wire \top_ihp.oisc.regs[29][20] ;
 wire \top_ihp.oisc.regs[29][21] ;
 wire \top_ihp.oisc.regs[29][22] ;
 wire \top_ihp.oisc.regs[29][23] ;
 wire \top_ihp.oisc.regs[29][24] ;
 wire \top_ihp.oisc.regs[29][25] ;
 wire \top_ihp.oisc.regs[29][26] ;
 wire \top_ihp.oisc.regs[29][27] ;
 wire \top_ihp.oisc.regs[29][28] ;
 wire \top_ihp.oisc.regs[29][29] ;
 wire \top_ihp.oisc.regs[29][2] ;
 wire \top_ihp.oisc.regs[29][30] ;
 wire \top_ihp.oisc.regs[29][31] ;
 wire \top_ihp.oisc.regs[29][3] ;
 wire \top_ihp.oisc.regs[29][4] ;
 wire \top_ihp.oisc.regs[29][5] ;
 wire \top_ihp.oisc.regs[29][6] ;
 wire \top_ihp.oisc.regs[29][7] ;
 wire \top_ihp.oisc.regs[29][8] ;
 wire \top_ihp.oisc.regs[29][9] ;
 wire \top_ihp.oisc.regs[2][0] ;
 wire \top_ihp.oisc.regs[2][10] ;
 wire \top_ihp.oisc.regs[2][11] ;
 wire \top_ihp.oisc.regs[2][12] ;
 wire \top_ihp.oisc.regs[2][13] ;
 wire \top_ihp.oisc.regs[2][14] ;
 wire \top_ihp.oisc.regs[2][15] ;
 wire \top_ihp.oisc.regs[2][16] ;
 wire \top_ihp.oisc.regs[2][17] ;
 wire \top_ihp.oisc.regs[2][18] ;
 wire \top_ihp.oisc.regs[2][19] ;
 wire \top_ihp.oisc.regs[2][1] ;
 wire \top_ihp.oisc.regs[2][20] ;
 wire \top_ihp.oisc.regs[2][21] ;
 wire \top_ihp.oisc.regs[2][22] ;
 wire \top_ihp.oisc.regs[2][23] ;
 wire \top_ihp.oisc.regs[2][24] ;
 wire \top_ihp.oisc.regs[2][25] ;
 wire \top_ihp.oisc.regs[2][26] ;
 wire \top_ihp.oisc.regs[2][27] ;
 wire \top_ihp.oisc.regs[2][28] ;
 wire \top_ihp.oisc.regs[2][29] ;
 wire \top_ihp.oisc.regs[2][2] ;
 wire \top_ihp.oisc.regs[2][30] ;
 wire \top_ihp.oisc.regs[2][31] ;
 wire \top_ihp.oisc.regs[2][3] ;
 wire \top_ihp.oisc.regs[2][4] ;
 wire \top_ihp.oisc.regs[2][5] ;
 wire \top_ihp.oisc.regs[2][6] ;
 wire \top_ihp.oisc.regs[2][7] ;
 wire \top_ihp.oisc.regs[2][8] ;
 wire \top_ihp.oisc.regs[2][9] ;
 wire \top_ihp.oisc.regs[30][0] ;
 wire \top_ihp.oisc.regs[30][10] ;
 wire \top_ihp.oisc.regs[30][11] ;
 wire \top_ihp.oisc.regs[30][12] ;
 wire \top_ihp.oisc.regs[30][13] ;
 wire \top_ihp.oisc.regs[30][14] ;
 wire \top_ihp.oisc.regs[30][15] ;
 wire \top_ihp.oisc.regs[30][16] ;
 wire \top_ihp.oisc.regs[30][17] ;
 wire \top_ihp.oisc.regs[30][18] ;
 wire \top_ihp.oisc.regs[30][19] ;
 wire \top_ihp.oisc.regs[30][1] ;
 wire \top_ihp.oisc.regs[30][20] ;
 wire \top_ihp.oisc.regs[30][21] ;
 wire \top_ihp.oisc.regs[30][22] ;
 wire \top_ihp.oisc.regs[30][23] ;
 wire \top_ihp.oisc.regs[30][24] ;
 wire \top_ihp.oisc.regs[30][25] ;
 wire \top_ihp.oisc.regs[30][26] ;
 wire \top_ihp.oisc.regs[30][27] ;
 wire \top_ihp.oisc.regs[30][28] ;
 wire \top_ihp.oisc.regs[30][29] ;
 wire \top_ihp.oisc.regs[30][2] ;
 wire \top_ihp.oisc.regs[30][30] ;
 wire \top_ihp.oisc.regs[30][31] ;
 wire \top_ihp.oisc.regs[30][3] ;
 wire \top_ihp.oisc.regs[30][4] ;
 wire \top_ihp.oisc.regs[30][5] ;
 wire \top_ihp.oisc.regs[30][6] ;
 wire \top_ihp.oisc.regs[30][7] ;
 wire \top_ihp.oisc.regs[30][8] ;
 wire \top_ihp.oisc.regs[30][9] ;
 wire \top_ihp.oisc.regs[31][0] ;
 wire \top_ihp.oisc.regs[31][10] ;
 wire \top_ihp.oisc.regs[31][11] ;
 wire \top_ihp.oisc.regs[31][12] ;
 wire \top_ihp.oisc.regs[31][13] ;
 wire \top_ihp.oisc.regs[31][14] ;
 wire \top_ihp.oisc.regs[31][15] ;
 wire \top_ihp.oisc.regs[31][16] ;
 wire \top_ihp.oisc.regs[31][17] ;
 wire \top_ihp.oisc.regs[31][18] ;
 wire \top_ihp.oisc.regs[31][19] ;
 wire \top_ihp.oisc.regs[31][1] ;
 wire \top_ihp.oisc.regs[31][20] ;
 wire \top_ihp.oisc.regs[31][21] ;
 wire \top_ihp.oisc.regs[31][22] ;
 wire \top_ihp.oisc.regs[31][23] ;
 wire \top_ihp.oisc.regs[31][24] ;
 wire \top_ihp.oisc.regs[31][25] ;
 wire \top_ihp.oisc.regs[31][26] ;
 wire \top_ihp.oisc.regs[31][27] ;
 wire \top_ihp.oisc.regs[31][28] ;
 wire \top_ihp.oisc.regs[31][29] ;
 wire \top_ihp.oisc.regs[31][2] ;
 wire \top_ihp.oisc.regs[31][30] ;
 wire \top_ihp.oisc.regs[31][31] ;
 wire \top_ihp.oisc.regs[31][3] ;
 wire \top_ihp.oisc.regs[31][4] ;
 wire \top_ihp.oisc.regs[31][5] ;
 wire \top_ihp.oisc.regs[31][6] ;
 wire \top_ihp.oisc.regs[31][7] ;
 wire \top_ihp.oisc.regs[31][8] ;
 wire \top_ihp.oisc.regs[31][9] ;
 wire \top_ihp.oisc.regs[32][0] ;
 wire \top_ihp.oisc.regs[32][10] ;
 wire \top_ihp.oisc.regs[32][11] ;
 wire \top_ihp.oisc.regs[32][12] ;
 wire \top_ihp.oisc.regs[32][13] ;
 wire \top_ihp.oisc.regs[32][14] ;
 wire \top_ihp.oisc.regs[32][15] ;
 wire \top_ihp.oisc.regs[32][16] ;
 wire \top_ihp.oisc.regs[32][17] ;
 wire \top_ihp.oisc.regs[32][18] ;
 wire \top_ihp.oisc.regs[32][19] ;
 wire \top_ihp.oisc.regs[32][1] ;
 wire \top_ihp.oisc.regs[32][20] ;
 wire \top_ihp.oisc.regs[32][21] ;
 wire \top_ihp.oisc.regs[32][22] ;
 wire \top_ihp.oisc.regs[32][23] ;
 wire \top_ihp.oisc.regs[32][24] ;
 wire \top_ihp.oisc.regs[32][25] ;
 wire \top_ihp.oisc.regs[32][26] ;
 wire \top_ihp.oisc.regs[32][27] ;
 wire \top_ihp.oisc.regs[32][28] ;
 wire \top_ihp.oisc.regs[32][29] ;
 wire \top_ihp.oisc.regs[32][2] ;
 wire \top_ihp.oisc.regs[32][30] ;
 wire \top_ihp.oisc.regs[32][31] ;
 wire \top_ihp.oisc.regs[32][3] ;
 wire \top_ihp.oisc.regs[32][4] ;
 wire \top_ihp.oisc.regs[32][5] ;
 wire \top_ihp.oisc.regs[32][6] ;
 wire \top_ihp.oisc.regs[32][7] ;
 wire \top_ihp.oisc.regs[32][8] ;
 wire \top_ihp.oisc.regs[32][9] ;
 wire \top_ihp.oisc.regs[33][0] ;
 wire \top_ihp.oisc.regs[33][10] ;
 wire \top_ihp.oisc.regs[33][11] ;
 wire \top_ihp.oisc.regs[33][12] ;
 wire \top_ihp.oisc.regs[33][13] ;
 wire \top_ihp.oisc.regs[33][14] ;
 wire \top_ihp.oisc.regs[33][15] ;
 wire \top_ihp.oisc.regs[33][16] ;
 wire \top_ihp.oisc.regs[33][17] ;
 wire \top_ihp.oisc.regs[33][18] ;
 wire \top_ihp.oisc.regs[33][19] ;
 wire \top_ihp.oisc.regs[33][1] ;
 wire \top_ihp.oisc.regs[33][20] ;
 wire \top_ihp.oisc.regs[33][21] ;
 wire \top_ihp.oisc.regs[33][22] ;
 wire \top_ihp.oisc.regs[33][23] ;
 wire \top_ihp.oisc.regs[33][24] ;
 wire \top_ihp.oisc.regs[33][25] ;
 wire \top_ihp.oisc.regs[33][26] ;
 wire \top_ihp.oisc.regs[33][27] ;
 wire \top_ihp.oisc.regs[33][28] ;
 wire \top_ihp.oisc.regs[33][29] ;
 wire \top_ihp.oisc.regs[33][2] ;
 wire \top_ihp.oisc.regs[33][30] ;
 wire \top_ihp.oisc.regs[33][31] ;
 wire \top_ihp.oisc.regs[33][3] ;
 wire \top_ihp.oisc.regs[33][4] ;
 wire \top_ihp.oisc.regs[33][5] ;
 wire \top_ihp.oisc.regs[33][6] ;
 wire \top_ihp.oisc.regs[33][7] ;
 wire \top_ihp.oisc.regs[33][8] ;
 wire \top_ihp.oisc.regs[33][9] ;
 wire \top_ihp.oisc.regs[34][0] ;
 wire \top_ihp.oisc.regs[34][10] ;
 wire \top_ihp.oisc.regs[34][11] ;
 wire \top_ihp.oisc.regs[34][12] ;
 wire \top_ihp.oisc.regs[34][13] ;
 wire \top_ihp.oisc.regs[34][14] ;
 wire \top_ihp.oisc.regs[34][15] ;
 wire \top_ihp.oisc.regs[34][16] ;
 wire \top_ihp.oisc.regs[34][17] ;
 wire \top_ihp.oisc.regs[34][18] ;
 wire \top_ihp.oisc.regs[34][19] ;
 wire \top_ihp.oisc.regs[34][1] ;
 wire \top_ihp.oisc.regs[34][20] ;
 wire \top_ihp.oisc.regs[34][21] ;
 wire \top_ihp.oisc.regs[34][22] ;
 wire \top_ihp.oisc.regs[34][23] ;
 wire \top_ihp.oisc.regs[34][24] ;
 wire \top_ihp.oisc.regs[34][25] ;
 wire \top_ihp.oisc.regs[34][26] ;
 wire \top_ihp.oisc.regs[34][27] ;
 wire \top_ihp.oisc.regs[34][28] ;
 wire \top_ihp.oisc.regs[34][29] ;
 wire \top_ihp.oisc.regs[34][2] ;
 wire \top_ihp.oisc.regs[34][30] ;
 wire \top_ihp.oisc.regs[34][31] ;
 wire \top_ihp.oisc.regs[34][3] ;
 wire \top_ihp.oisc.regs[34][4] ;
 wire \top_ihp.oisc.regs[34][5] ;
 wire \top_ihp.oisc.regs[34][6] ;
 wire \top_ihp.oisc.regs[34][7] ;
 wire \top_ihp.oisc.regs[34][8] ;
 wire \top_ihp.oisc.regs[34][9] ;
 wire \top_ihp.oisc.regs[35][0] ;
 wire \top_ihp.oisc.regs[35][10] ;
 wire \top_ihp.oisc.regs[35][11] ;
 wire \top_ihp.oisc.regs[35][12] ;
 wire \top_ihp.oisc.regs[35][13] ;
 wire \top_ihp.oisc.regs[35][14] ;
 wire \top_ihp.oisc.regs[35][15] ;
 wire \top_ihp.oisc.regs[35][16] ;
 wire \top_ihp.oisc.regs[35][17] ;
 wire \top_ihp.oisc.regs[35][18] ;
 wire \top_ihp.oisc.regs[35][19] ;
 wire \top_ihp.oisc.regs[35][1] ;
 wire \top_ihp.oisc.regs[35][20] ;
 wire \top_ihp.oisc.regs[35][21] ;
 wire \top_ihp.oisc.regs[35][22] ;
 wire \top_ihp.oisc.regs[35][23] ;
 wire \top_ihp.oisc.regs[35][24] ;
 wire \top_ihp.oisc.regs[35][25] ;
 wire \top_ihp.oisc.regs[35][26] ;
 wire \top_ihp.oisc.regs[35][27] ;
 wire \top_ihp.oisc.regs[35][28] ;
 wire \top_ihp.oisc.regs[35][29] ;
 wire \top_ihp.oisc.regs[35][2] ;
 wire \top_ihp.oisc.regs[35][30] ;
 wire \top_ihp.oisc.regs[35][31] ;
 wire \top_ihp.oisc.regs[35][3] ;
 wire \top_ihp.oisc.regs[35][4] ;
 wire \top_ihp.oisc.regs[35][5] ;
 wire \top_ihp.oisc.regs[35][6] ;
 wire \top_ihp.oisc.regs[35][7] ;
 wire \top_ihp.oisc.regs[35][8] ;
 wire \top_ihp.oisc.regs[35][9] ;
 wire \top_ihp.oisc.regs[36][0] ;
 wire \top_ihp.oisc.regs[36][10] ;
 wire \top_ihp.oisc.regs[36][11] ;
 wire \top_ihp.oisc.regs[36][12] ;
 wire \top_ihp.oisc.regs[36][13] ;
 wire \top_ihp.oisc.regs[36][14] ;
 wire \top_ihp.oisc.regs[36][15] ;
 wire \top_ihp.oisc.regs[36][16] ;
 wire \top_ihp.oisc.regs[36][17] ;
 wire \top_ihp.oisc.regs[36][18] ;
 wire \top_ihp.oisc.regs[36][19] ;
 wire \top_ihp.oisc.regs[36][1] ;
 wire \top_ihp.oisc.regs[36][20] ;
 wire \top_ihp.oisc.regs[36][21] ;
 wire \top_ihp.oisc.regs[36][22] ;
 wire \top_ihp.oisc.regs[36][23] ;
 wire \top_ihp.oisc.regs[36][24] ;
 wire \top_ihp.oisc.regs[36][25] ;
 wire \top_ihp.oisc.regs[36][26] ;
 wire \top_ihp.oisc.regs[36][27] ;
 wire \top_ihp.oisc.regs[36][28] ;
 wire \top_ihp.oisc.regs[36][29] ;
 wire \top_ihp.oisc.regs[36][2] ;
 wire \top_ihp.oisc.regs[36][30] ;
 wire \top_ihp.oisc.regs[36][31] ;
 wire \top_ihp.oisc.regs[36][3] ;
 wire \top_ihp.oisc.regs[36][4] ;
 wire \top_ihp.oisc.regs[36][5] ;
 wire \top_ihp.oisc.regs[36][6] ;
 wire \top_ihp.oisc.regs[36][7] ;
 wire \top_ihp.oisc.regs[36][8] ;
 wire \top_ihp.oisc.regs[36][9] ;
 wire \top_ihp.oisc.regs[37][0] ;
 wire \top_ihp.oisc.regs[37][10] ;
 wire \top_ihp.oisc.regs[37][11] ;
 wire \top_ihp.oisc.regs[37][12] ;
 wire \top_ihp.oisc.regs[37][13] ;
 wire \top_ihp.oisc.regs[37][14] ;
 wire \top_ihp.oisc.regs[37][15] ;
 wire \top_ihp.oisc.regs[37][16] ;
 wire \top_ihp.oisc.regs[37][17] ;
 wire \top_ihp.oisc.regs[37][18] ;
 wire \top_ihp.oisc.regs[37][19] ;
 wire \top_ihp.oisc.regs[37][1] ;
 wire \top_ihp.oisc.regs[37][20] ;
 wire \top_ihp.oisc.regs[37][21] ;
 wire \top_ihp.oisc.regs[37][22] ;
 wire \top_ihp.oisc.regs[37][23] ;
 wire \top_ihp.oisc.regs[37][24] ;
 wire \top_ihp.oisc.regs[37][25] ;
 wire \top_ihp.oisc.regs[37][26] ;
 wire \top_ihp.oisc.regs[37][27] ;
 wire \top_ihp.oisc.regs[37][28] ;
 wire \top_ihp.oisc.regs[37][29] ;
 wire \top_ihp.oisc.regs[37][2] ;
 wire \top_ihp.oisc.regs[37][30] ;
 wire \top_ihp.oisc.regs[37][31] ;
 wire \top_ihp.oisc.regs[37][3] ;
 wire \top_ihp.oisc.regs[37][4] ;
 wire \top_ihp.oisc.regs[37][5] ;
 wire \top_ihp.oisc.regs[37][6] ;
 wire \top_ihp.oisc.regs[37][7] ;
 wire \top_ihp.oisc.regs[37][8] ;
 wire \top_ihp.oisc.regs[37][9] ;
 wire \top_ihp.oisc.regs[38][0] ;
 wire \top_ihp.oisc.regs[38][10] ;
 wire \top_ihp.oisc.regs[38][11] ;
 wire \top_ihp.oisc.regs[38][12] ;
 wire \top_ihp.oisc.regs[38][13] ;
 wire \top_ihp.oisc.regs[38][14] ;
 wire \top_ihp.oisc.regs[38][15] ;
 wire \top_ihp.oisc.regs[38][16] ;
 wire \top_ihp.oisc.regs[38][17] ;
 wire \top_ihp.oisc.regs[38][18] ;
 wire \top_ihp.oisc.regs[38][19] ;
 wire \top_ihp.oisc.regs[38][1] ;
 wire \top_ihp.oisc.regs[38][20] ;
 wire \top_ihp.oisc.regs[38][21] ;
 wire \top_ihp.oisc.regs[38][22] ;
 wire \top_ihp.oisc.regs[38][23] ;
 wire \top_ihp.oisc.regs[38][24] ;
 wire \top_ihp.oisc.regs[38][25] ;
 wire \top_ihp.oisc.regs[38][26] ;
 wire \top_ihp.oisc.regs[38][27] ;
 wire \top_ihp.oisc.regs[38][28] ;
 wire \top_ihp.oisc.regs[38][29] ;
 wire \top_ihp.oisc.regs[38][2] ;
 wire \top_ihp.oisc.regs[38][30] ;
 wire \top_ihp.oisc.regs[38][31] ;
 wire \top_ihp.oisc.regs[38][3] ;
 wire \top_ihp.oisc.regs[38][4] ;
 wire \top_ihp.oisc.regs[38][5] ;
 wire \top_ihp.oisc.regs[38][6] ;
 wire \top_ihp.oisc.regs[38][7] ;
 wire \top_ihp.oisc.regs[38][8] ;
 wire \top_ihp.oisc.regs[38][9] ;
 wire \top_ihp.oisc.regs[39][0] ;
 wire \top_ihp.oisc.regs[39][10] ;
 wire \top_ihp.oisc.regs[39][11] ;
 wire \top_ihp.oisc.regs[39][12] ;
 wire \top_ihp.oisc.regs[39][13] ;
 wire \top_ihp.oisc.regs[39][14] ;
 wire \top_ihp.oisc.regs[39][15] ;
 wire \top_ihp.oisc.regs[39][16] ;
 wire \top_ihp.oisc.regs[39][17] ;
 wire \top_ihp.oisc.regs[39][18] ;
 wire \top_ihp.oisc.regs[39][19] ;
 wire \top_ihp.oisc.regs[39][1] ;
 wire \top_ihp.oisc.regs[39][20] ;
 wire \top_ihp.oisc.regs[39][21] ;
 wire \top_ihp.oisc.regs[39][22] ;
 wire \top_ihp.oisc.regs[39][23] ;
 wire \top_ihp.oisc.regs[39][24] ;
 wire \top_ihp.oisc.regs[39][25] ;
 wire \top_ihp.oisc.regs[39][26] ;
 wire \top_ihp.oisc.regs[39][27] ;
 wire \top_ihp.oisc.regs[39][28] ;
 wire \top_ihp.oisc.regs[39][29] ;
 wire \top_ihp.oisc.regs[39][2] ;
 wire \top_ihp.oisc.regs[39][30] ;
 wire \top_ihp.oisc.regs[39][31] ;
 wire \top_ihp.oisc.regs[39][3] ;
 wire \top_ihp.oisc.regs[39][4] ;
 wire \top_ihp.oisc.regs[39][5] ;
 wire \top_ihp.oisc.regs[39][6] ;
 wire \top_ihp.oisc.regs[39][7] ;
 wire \top_ihp.oisc.regs[39][8] ;
 wire \top_ihp.oisc.regs[39][9] ;
 wire \top_ihp.oisc.regs[3][0] ;
 wire \top_ihp.oisc.regs[3][10] ;
 wire \top_ihp.oisc.regs[3][11] ;
 wire \top_ihp.oisc.regs[3][12] ;
 wire \top_ihp.oisc.regs[3][13] ;
 wire \top_ihp.oisc.regs[3][14] ;
 wire \top_ihp.oisc.regs[3][15] ;
 wire \top_ihp.oisc.regs[3][16] ;
 wire \top_ihp.oisc.regs[3][17] ;
 wire \top_ihp.oisc.regs[3][18] ;
 wire \top_ihp.oisc.regs[3][19] ;
 wire \top_ihp.oisc.regs[3][1] ;
 wire \top_ihp.oisc.regs[3][20] ;
 wire \top_ihp.oisc.regs[3][21] ;
 wire \top_ihp.oisc.regs[3][22] ;
 wire \top_ihp.oisc.regs[3][23] ;
 wire \top_ihp.oisc.regs[3][24] ;
 wire \top_ihp.oisc.regs[3][25] ;
 wire \top_ihp.oisc.regs[3][26] ;
 wire \top_ihp.oisc.regs[3][27] ;
 wire \top_ihp.oisc.regs[3][28] ;
 wire \top_ihp.oisc.regs[3][29] ;
 wire \top_ihp.oisc.regs[3][2] ;
 wire \top_ihp.oisc.regs[3][30] ;
 wire \top_ihp.oisc.regs[3][31] ;
 wire \top_ihp.oisc.regs[3][3] ;
 wire \top_ihp.oisc.regs[3][4] ;
 wire \top_ihp.oisc.regs[3][5] ;
 wire \top_ihp.oisc.regs[3][6] ;
 wire \top_ihp.oisc.regs[3][7] ;
 wire \top_ihp.oisc.regs[3][8] ;
 wire \top_ihp.oisc.regs[3][9] ;
 wire \top_ihp.oisc.regs[40][0] ;
 wire \top_ihp.oisc.regs[40][10] ;
 wire \top_ihp.oisc.regs[40][11] ;
 wire \top_ihp.oisc.regs[40][12] ;
 wire \top_ihp.oisc.regs[40][13] ;
 wire \top_ihp.oisc.regs[40][14] ;
 wire \top_ihp.oisc.regs[40][15] ;
 wire \top_ihp.oisc.regs[40][16] ;
 wire \top_ihp.oisc.regs[40][17] ;
 wire \top_ihp.oisc.regs[40][18] ;
 wire \top_ihp.oisc.regs[40][19] ;
 wire \top_ihp.oisc.regs[40][1] ;
 wire \top_ihp.oisc.regs[40][20] ;
 wire \top_ihp.oisc.regs[40][21] ;
 wire \top_ihp.oisc.regs[40][22] ;
 wire \top_ihp.oisc.regs[40][23] ;
 wire \top_ihp.oisc.regs[40][24] ;
 wire \top_ihp.oisc.regs[40][25] ;
 wire \top_ihp.oisc.regs[40][26] ;
 wire \top_ihp.oisc.regs[40][27] ;
 wire \top_ihp.oisc.regs[40][28] ;
 wire \top_ihp.oisc.regs[40][29] ;
 wire \top_ihp.oisc.regs[40][2] ;
 wire \top_ihp.oisc.regs[40][30] ;
 wire \top_ihp.oisc.regs[40][31] ;
 wire \top_ihp.oisc.regs[40][3] ;
 wire \top_ihp.oisc.regs[40][4] ;
 wire \top_ihp.oisc.regs[40][5] ;
 wire \top_ihp.oisc.regs[40][6] ;
 wire \top_ihp.oisc.regs[40][7] ;
 wire \top_ihp.oisc.regs[40][8] ;
 wire \top_ihp.oisc.regs[40][9] ;
 wire \top_ihp.oisc.regs[41][0] ;
 wire \top_ihp.oisc.regs[41][10] ;
 wire \top_ihp.oisc.regs[41][11] ;
 wire \top_ihp.oisc.regs[41][12] ;
 wire \top_ihp.oisc.regs[41][13] ;
 wire \top_ihp.oisc.regs[41][14] ;
 wire \top_ihp.oisc.regs[41][15] ;
 wire \top_ihp.oisc.regs[41][16] ;
 wire \top_ihp.oisc.regs[41][17] ;
 wire \top_ihp.oisc.regs[41][18] ;
 wire \top_ihp.oisc.regs[41][19] ;
 wire \top_ihp.oisc.regs[41][1] ;
 wire \top_ihp.oisc.regs[41][20] ;
 wire \top_ihp.oisc.regs[41][21] ;
 wire \top_ihp.oisc.regs[41][22] ;
 wire \top_ihp.oisc.regs[41][23] ;
 wire \top_ihp.oisc.regs[41][24] ;
 wire \top_ihp.oisc.regs[41][25] ;
 wire \top_ihp.oisc.regs[41][26] ;
 wire \top_ihp.oisc.regs[41][27] ;
 wire \top_ihp.oisc.regs[41][28] ;
 wire \top_ihp.oisc.regs[41][29] ;
 wire \top_ihp.oisc.regs[41][2] ;
 wire \top_ihp.oisc.regs[41][30] ;
 wire \top_ihp.oisc.regs[41][31] ;
 wire \top_ihp.oisc.regs[41][3] ;
 wire \top_ihp.oisc.regs[41][4] ;
 wire \top_ihp.oisc.regs[41][5] ;
 wire \top_ihp.oisc.regs[41][6] ;
 wire \top_ihp.oisc.regs[41][7] ;
 wire \top_ihp.oisc.regs[41][8] ;
 wire \top_ihp.oisc.regs[41][9] ;
 wire \top_ihp.oisc.regs[42][0] ;
 wire \top_ihp.oisc.regs[42][10] ;
 wire \top_ihp.oisc.regs[42][11] ;
 wire \top_ihp.oisc.regs[42][12] ;
 wire \top_ihp.oisc.regs[42][13] ;
 wire \top_ihp.oisc.regs[42][14] ;
 wire \top_ihp.oisc.regs[42][15] ;
 wire \top_ihp.oisc.regs[42][16] ;
 wire \top_ihp.oisc.regs[42][17] ;
 wire \top_ihp.oisc.regs[42][18] ;
 wire \top_ihp.oisc.regs[42][19] ;
 wire \top_ihp.oisc.regs[42][1] ;
 wire \top_ihp.oisc.regs[42][20] ;
 wire \top_ihp.oisc.regs[42][21] ;
 wire \top_ihp.oisc.regs[42][22] ;
 wire \top_ihp.oisc.regs[42][23] ;
 wire \top_ihp.oisc.regs[42][24] ;
 wire \top_ihp.oisc.regs[42][25] ;
 wire \top_ihp.oisc.regs[42][26] ;
 wire \top_ihp.oisc.regs[42][27] ;
 wire \top_ihp.oisc.regs[42][28] ;
 wire \top_ihp.oisc.regs[42][29] ;
 wire \top_ihp.oisc.regs[42][2] ;
 wire \top_ihp.oisc.regs[42][30] ;
 wire \top_ihp.oisc.regs[42][31] ;
 wire \top_ihp.oisc.regs[42][3] ;
 wire \top_ihp.oisc.regs[42][4] ;
 wire \top_ihp.oisc.regs[42][5] ;
 wire \top_ihp.oisc.regs[42][6] ;
 wire \top_ihp.oisc.regs[42][7] ;
 wire \top_ihp.oisc.regs[42][8] ;
 wire \top_ihp.oisc.regs[42][9] ;
 wire \top_ihp.oisc.regs[43][0] ;
 wire \top_ihp.oisc.regs[43][10] ;
 wire \top_ihp.oisc.regs[43][11] ;
 wire \top_ihp.oisc.regs[43][12] ;
 wire \top_ihp.oisc.regs[43][13] ;
 wire \top_ihp.oisc.regs[43][14] ;
 wire \top_ihp.oisc.regs[43][15] ;
 wire \top_ihp.oisc.regs[43][16] ;
 wire \top_ihp.oisc.regs[43][17] ;
 wire \top_ihp.oisc.regs[43][18] ;
 wire \top_ihp.oisc.regs[43][19] ;
 wire \top_ihp.oisc.regs[43][1] ;
 wire \top_ihp.oisc.regs[43][20] ;
 wire \top_ihp.oisc.regs[43][21] ;
 wire \top_ihp.oisc.regs[43][22] ;
 wire \top_ihp.oisc.regs[43][23] ;
 wire \top_ihp.oisc.regs[43][24] ;
 wire \top_ihp.oisc.regs[43][25] ;
 wire \top_ihp.oisc.regs[43][26] ;
 wire \top_ihp.oisc.regs[43][27] ;
 wire \top_ihp.oisc.regs[43][28] ;
 wire \top_ihp.oisc.regs[43][29] ;
 wire \top_ihp.oisc.regs[43][2] ;
 wire \top_ihp.oisc.regs[43][30] ;
 wire \top_ihp.oisc.regs[43][31] ;
 wire \top_ihp.oisc.regs[43][3] ;
 wire \top_ihp.oisc.regs[43][4] ;
 wire \top_ihp.oisc.regs[43][5] ;
 wire \top_ihp.oisc.regs[43][6] ;
 wire \top_ihp.oisc.regs[43][7] ;
 wire \top_ihp.oisc.regs[43][8] ;
 wire \top_ihp.oisc.regs[43][9] ;
 wire \top_ihp.oisc.regs[44][0] ;
 wire \top_ihp.oisc.regs[44][10] ;
 wire \top_ihp.oisc.regs[44][11] ;
 wire \top_ihp.oisc.regs[44][12] ;
 wire \top_ihp.oisc.regs[44][13] ;
 wire \top_ihp.oisc.regs[44][14] ;
 wire \top_ihp.oisc.regs[44][15] ;
 wire \top_ihp.oisc.regs[44][16] ;
 wire \top_ihp.oisc.regs[44][17] ;
 wire \top_ihp.oisc.regs[44][18] ;
 wire \top_ihp.oisc.regs[44][19] ;
 wire \top_ihp.oisc.regs[44][1] ;
 wire \top_ihp.oisc.regs[44][20] ;
 wire \top_ihp.oisc.regs[44][21] ;
 wire \top_ihp.oisc.regs[44][22] ;
 wire \top_ihp.oisc.regs[44][23] ;
 wire \top_ihp.oisc.regs[44][24] ;
 wire \top_ihp.oisc.regs[44][25] ;
 wire \top_ihp.oisc.regs[44][26] ;
 wire \top_ihp.oisc.regs[44][27] ;
 wire \top_ihp.oisc.regs[44][28] ;
 wire \top_ihp.oisc.regs[44][29] ;
 wire \top_ihp.oisc.regs[44][2] ;
 wire \top_ihp.oisc.regs[44][30] ;
 wire \top_ihp.oisc.regs[44][31] ;
 wire \top_ihp.oisc.regs[44][3] ;
 wire \top_ihp.oisc.regs[44][4] ;
 wire \top_ihp.oisc.regs[44][5] ;
 wire \top_ihp.oisc.regs[44][6] ;
 wire \top_ihp.oisc.regs[44][7] ;
 wire \top_ihp.oisc.regs[44][8] ;
 wire \top_ihp.oisc.regs[44][9] ;
 wire \top_ihp.oisc.regs[45][0] ;
 wire \top_ihp.oisc.regs[45][10] ;
 wire \top_ihp.oisc.regs[45][11] ;
 wire \top_ihp.oisc.regs[45][12] ;
 wire \top_ihp.oisc.regs[45][13] ;
 wire \top_ihp.oisc.regs[45][14] ;
 wire \top_ihp.oisc.regs[45][15] ;
 wire \top_ihp.oisc.regs[45][16] ;
 wire \top_ihp.oisc.regs[45][17] ;
 wire \top_ihp.oisc.regs[45][18] ;
 wire \top_ihp.oisc.regs[45][19] ;
 wire \top_ihp.oisc.regs[45][1] ;
 wire \top_ihp.oisc.regs[45][20] ;
 wire \top_ihp.oisc.regs[45][21] ;
 wire \top_ihp.oisc.regs[45][22] ;
 wire \top_ihp.oisc.regs[45][23] ;
 wire \top_ihp.oisc.regs[45][24] ;
 wire \top_ihp.oisc.regs[45][25] ;
 wire \top_ihp.oisc.regs[45][26] ;
 wire \top_ihp.oisc.regs[45][27] ;
 wire \top_ihp.oisc.regs[45][28] ;
 wire \top_ihp.oisc.regs[45][29] ;
 wire \top_ihp.oisc.regs[45][2] ;
 wire \top_ihp.oisc.regs[45][30] ;
 wire \top_ihp.oisc.regs[45][31] ;
 wire \top_ihp.oisc.regs[45][3] ;
 wire \top_ihp.oisc.regs[45][4] ;
 wire \top_ihp.oisc.regs[45][5] ;
 wire \top_ihp.oisc.regs[45][6] ;
 wire \top_ihp.oisc.regs[45][7] ;
 wire \top_ihp.oisc.regs[45][8] ;
 wire \top_ihp.oisc.regs[45][9] ;
 wire \top_ihp.oisc.regs[46][0] ;
 wire \top_ihp.oisc.regs[46][10] ;
 wire \top_ihp.oisc.regs[46][11] ;
 wire \top_ihp.oisc.regs[46][12] ;
 wire \top_ihp.oisc.regs[46][13] ;
 wire \top_ihp.oisc.regs[46][14] ;
 wire \top_ihp.oisc.regs[46][15] ;
 wire \top_ihp.oisc.regs[46][16] ;
 wire \top_ihp.oisc.regs[46][17] ;
 wire \top_ihp.oisc.regs[46][18] ;
 wire \top_ihp.oisc.regs[46][19] ;
 wire \top_ihp.oisc.regs[46][1] ;
 wire \top_ihp.oisc.regs[46][20] ;
 wire \top_ihp.oisc.regs[46][21] ;
 wire \top_ihp.oisc.regs[46][22] ;
 wire \top_ihp.oisc.regs[46][23] ;
 wire \top_ihp.oisc.regs[46][24] ;
 wire \top_ihp.oisc.regs[46][25] ;
 wire \top_ihp.oisc.regs[46][26] ;
 wire \top_ihp.oisc.regs[46][27] ;
 wire \top_ihp.oisc.regs[46][28] ;
 wire \top_ihp.oisc.regs[46][29] ;
 wire \top_ihp.oisc.regs[46][2] ;
 wire \top_ihp.oisc.regs[46][30] ;
 wire \top_ihp.oisc.regs[46][31] ;
 wire \top_ihp.oisc.regs[46][3] ;
 wire \top_ihp.oisc.regs[46][4] ;
 wire \top_ihp.oisc.regs[46][5] ;
 wire \top_ihp.oisc.regs[46][6] ;
 wire \top_ihp.oisc.regs[46][7] ;
 wire \top_ihp.oisc.regs[46][8] ;
 wire \top_ihp.oisc.regs[46][9] ;
 wire \top_ihp.oisc.regs[47][0] ;
 wire \top_ihp.oisc.regs[47][10] ;
 wire \top_ihp.oisc.regs[47][11] ;
 wire \top_ihp.oisc.regs[47][12] ;
 wire \top_ihp.oisc.regs[47][13] ;
 wire \top_ihp.oisc.regs[47][14] ;
 wire \top_ihp.oisc.regs[47][15] ;
 wire \top_ihp.oisc.regs[47][16] ;
 wire \top_ihp.oisc.regs[47][17] ;
 wire \top_ihp.oisc.regs[47][18] ;
 wire \top_ihp.oisc.regs[47][19] ;
 wire \top_ihp.oisc.regs[47][1] ;
 wire \top_ihp.oisc.regs[47][20] ;
 wire \top_ihp.oisc.regs[47][21] ;
 wire \top_ihp.oisc.regs[47][22] ;
 wire \top_ihp.oisc.regs[47][23] ;
 wire \top_ihp.oisc.regs[47][24] ;
 wire \top_ihp.oisc.regs[47][25] ;
 wire \top_ihp.oisc.regs[47][26] ;
 wire \top_ihp.oisc.regs[47][27] ;
 wire \top_ihp.oisc.regs[47][28] ;
 wire \top_ihp.oisc.regs[47][29] ;
 wire \top_ihp.oisc.regs[47][2] ;
 wire \top_ihp.oisc.regs[47][30] ;
 wire \top_ihp.oisc.regs[47][31] ;
 wire \top_ihp.oisc.regs[47][3] ;
 wire \top_ihp.oisc.regs[47][4] ;
 wire \top_ihp.oisc.regs[47][5] ;
 wire \top_ihp.oisc.regs[47][6] ;
 wire \top_ihp.oisc.regs[47][7] ;
 wire \top_ihp.oisc.regs[47][8] ;
 wire \top_ihp.oisc.regs[47][9] ;
 wire \top_ihp.oisc.regs[48][0] ;
 wire \top_ihp.oisc.regs[48][10] ;
 wire \top_ihp.oisc.regs[48][11] ;
 wire \top_ihp.oisc.regs[48][12] ;
 wire \top_ihp.oisc.regs[48][13] ;
 wire \top_ihp.oisc.regs[48][14] ;
 wire \top_ihp.oisc.regs[48][15] ;
 wire \top_ihp.oisc.regs[48][16] ;
 wire \top_ihp.oisc.regs[48][17] ;
 wire \top_ihp.oisc.regs[48][18] ;
 wire \top_ihp.oisc.regs[48][19] ;
 wire \top_ihp.oisc.regs[48][1] ;
 wire \top_ihp.oisc.regs[48][20] ;
 wire \top_ihp.oisc.regs[48][21] ;
 wire \top_ihp.oisc.regs[48][22] ;
 wire \top_ihp.oisc.regs[48][23] ;
 wire \top_ihp.oisc.regs[48][24] ;
 wire \top_ihp.oisc.regs[48][25] ;
 wire \top_ihp.oisc.regs[48][26] ;
 wire \top_ihp.oisc.regs[48][27] ;
 wire \top_ihp.oisc.regs[48][28] ;
 wire \top_ihp.oisc.regs[48][29] ;
 wire \top_ihp.oisc.regs[48][2] ;
 wire \top_ihp.oisc.regs[48][30] ;
 wire \top_ihp.oisc.regs[48][31] ;
 wire \top_ihp.oisc.regs[48][3] ;
 wire \top_ihp.oisc.regs[48][4] ;
 wire \top_ihp.oisc.regs[48][5] ;
 wire \top_ihp.oisc.regs[48][6] ;
 wire \top_ihp.oisc.regs[48][7] ;
 wire \top_ihp.oisc.regs[48][8] ;
 wire \top_ihp.oisc.regs[48][9] ;
 wire \top_ihp.oisc.regs[49][0] ;
 wire \top_ihp.oisc.regs[49][10] ;
 wire \top_ihp.oisc.regs[49][11] ;
 wire \top_ihp.oisc.regs[49][12] ;
 wire \top_ihp.oisc.regs[49][13] ;
 wire \top_ihp.oisc.regs[49][14] ;
 wire \top_ihp.oisc.regs[49][15] ;
 wire \top_ihp.oisc.regs[49][16] ;
 wire \top_ihp.oisc.regs[49][17] ;
 wire \top_ihp.oisc.regs[49][18] ;
 wire \top_ihp.oisc.regs[49][19] ;
 wire \top_ihp.oisc.regs[49][1] ;
 wire \top_ihp.oisc.regs[49][20] ;
 wire \top_ihp.oisc.regs[49][21] ;
 wire \top_ihp.oisc.regs[49][22] ;
 wire \top_ihp.oisc.regs[49][23] ;
 wire \top_ihp.oisc.regs[49][24] ;
 wire \top_ihp.oisc.regs[49][25] ;
 wire \top_ihp.oisc.regs[49][26] ;
 wire \top_ihp.oisc.regs[49][27] ;
 wire \top_ihp.oisc.regs[49][28] ;
 wire \top_ihp.oisc.regs[49][29] ;
 wire \top_ihp.oisc.regs[49][2] ;
 wire \top_ihp.oisc.regs[49][30] ;
 wire \top_ihp.oisc.regs[49][31] ;
 wire \top_ihp.oisc.regs[49][3] ;
 wire \top_ihp.oisc.regs[49][4] ;
 wire \top_ihp.oisc.regs[49][5] ;
 wire \top_ihp.oisc.regs[49][6] ;
 wire \top_ihp.oisc.regs[49][7] ;
 wire \top_ihp.oisc.regs[49][8] ;
 wire \top_ihp.oisc.regs[49][9] ;
 wire \top_ihp.oisc.regs[4][0] ;
 wire \top_ihp.oisc.regs[4][10] ;
 wire \top_ihp.oisc.regs[4][11] ;
 wire \top_ihp.oisc.regs[4][12] ;
 wire \top_ihp.oisc.regs[4][13] ;
 wire \top_ihp.oisc.regs[4][14] ;
 wire \top_ihp.oisc.regs[4][15] ;
 wire \top_ihp.oisc.regs[4][16] ;
 wire \top_ihp.oisc.regs[4][17] ;
 wire \top_ihp.oisc.regs[4][18] ;
 wire \top_ihp.oisc.regs[4][19] ;
 wire \top_ihp.oisc.regs[4][1] ;
 wire \top_ihp.oisc.regs[4][20] ;
 wire \top_ihp.oisc.regs[4][21] ;
 wire \top_ihp.oisc.regs[4][22] ;
 wire \top_ihp.oisc.regs[4][23] ;
 wire \top_ihp.oisc.regs[4][24] ;
 wire \top_ihp.oisc.regs[4][25] ;
 wire \top_ihp.oisc.regs[4][26] ;
 wire \top_ihp.oisc.regs[4][27] ;
 wire \top_ihp.oisc.regs[4][28] ;
 wire \top_ihp.oisc.regs[4][29] ;
 wire \top_ihp.oisc.regs[4][2] ;
 wire \top_ihp.oisc.regs[4][30] ;
 wire \top_ihp.oisc.regs[4][31] ;
 wire \top_ihp.oisc.regs[4][3] ;
 wire \top_ihp.oisc.regs[4][4] ;
 wire \top_ihp.oisc.regs[4][5] ;
 wire \top_ihp.oisc.regs[4][6] ;
 wire \top_ihp.oisc.regs[4][7] ;
 wire \top_ihp.oisc.regs[4][8] ;
 wire \top_ihp.oisc.regs[4][9] ;
 wire \top_ihp.oisc.regs[50][0] ;
 wire \top_ihp.oisc.regs[50][10] ;
 wire \top_ihp.oisc.regs[50][11] ;
 wire \top_ihp.oisc.regs[50][12] ;
 wire \top_ihp.oisc.regs[50][13] ;
 wire \top_ihp.oisc.regs[50][14] ;
 wire \top_ihp.oisc.regs[50][15] ;
 wire \top_ihp.oisc.regs[50][16] ;
 wire \top_ihp.oisc.regs[50][17] ;
 wire \top_ihp.oisc.regs[50][18] ;
 wire \top_ihp.oisc.regs[50][19] ;
 wire \top_ihp.oisc.regs[50][1] ;
 wire \top_ihp.oisc.regs[50][20] ;
 wire \top_ihp.oisc.regs[50][21] ;
 wire \top_ihp.oisc.regs[50][22] ;
 wire \top_ihp.oisc.regs[50][23] ;
 wire \top_ihp.oisc.regs[50][24] ;
 wire \top_ihp.oisc.regs[50][25] ;
 wire \top_ihp.oisc.regs[50][26] ;
 wire \top_ihp.oisc.regs[50][27] ;
 wire \top_ihp.oisc.regs[50][28] ;
 wire \top_ihp.oisc.regs[50][29] ;
 wire \top_ihp.oisc.regs[50][2] ;
 wire \top_ihp.oisc.regs[50][30] ;
 wire \top_ihp.oisc.regs[50][31] ;
 wire \top_ihp.oisc.regs[50][3] ;
 wire \top_ihp.oisc.regs[50][4] ;
 wire \top_ihp.oisc.regs[50][5] ;
 wire \top_ihp.oisc.regs[50][6] ;
 wire \top_ihp.oisc.regs[50][7] ;
 wire \top_ihp.oisc.regs[50][8] ;
 wire \top_ihp.oisc.regs[50][9] ;
 wire \top_ihp.oisc.regs[51][0] ;
 wire \top_ihp.oisc.regs[51][10] ;
 wire \top_ihp.oisc.regs[51][11] ;
 wire \top_ihp.oisc.regs[51][12] ;
 wire \top_ihp.oisc.regs[51][13] ;
 wire \top_ihp.oisc.regs[51][14] ;
 wire \top_ihp.oisc.regs[51][15] ;
 wire \top_ihp.oisc.regs[51][16] ;
 wire \top_ihp.oisc.regs[51][17] ;
 wire \top_ihp.oisc.regs[51][18] ;
 wire \top_ihp.oisc.regs[51][19] ;
 wire \top_ihp.oisc.regs[51][1] ;
 wire \top_ihp.oisc.regs[51][20] ;
 wire \top_ihp.oisc.regs[51][21] ;
 wire \top_ihp.oisc.regs[51][22] ;
 wire \top_ihp.oisc.regs[51][23] ;
 wire \top_ihp.oisc.regs[51][24] ;
 wire \top_ihp.oisc.regs[51][25] ;
 wire \top_ihp.oisc.regs[51][26] ;
 wire \top_ihp.oisc.regs[51][27] ;
 wire \top_ihp.oisc.regs[51][28] ;
 wire \top_ihp.oisc.regs[51][29] ;
 wire \top_ihp.oisc.regs[51][2] ;
 wire \top_ihp.oisc.regs[51][30] ;
 wire \top_ihp.oisc.regs[51][31] ;
 wire \top_ihp.oisc.regs[51][3] ;
 wire \top_ihp.oisc.regs[51][4] ;
 wire \top_ihp.oisc.regs[51][5] ;
 wire \top_ihp.oisc.regs[51][6] ;
 wire \top_ihp.oisc.regs[51][7] ;
 wire \top_ihp.oisc.regs[51][8] ;
 wire \top_ihp.oisc.regs[51][9] ;
 wire \top_ihp.oisc.regs[52][0] ;
 wire \top_ihp.oisc.regs[52][10] ;
 wire \top_ihp.oisc.regs[52][11] ;
 wire \top_ihp.oisc.regs[52][12] ;
 wire \top_ihp.oisc.regs[52][13] ;
 wire \top_ihp.oisc.regs[52][14] ;
 wire \top_ihp.oisc.regs[52][15] ;
 wire \top_ihp.oisc.regs[52][16] ;
 wire \top_ihp.oisc.regs[52][17] ;
 wire \top_ihp.oisc.regs[52][18] ;
 wire \top_ihp.oisc.regs[52][19] ;
 wire \top_ihp.oisc.regs[52][1] ;
 wire \top_ihp.oisc.regs[52][20] ;
 wire \top_ihp.oisc.regs[52][21] ;
 wire \top_ihp.oisc.regs[52][22] ;
 wire \top_ihp.oisc.regs[52][23] ;
 wire \top_ihp.oisc.regs[52][24] ;
 wire \top_ihp.oisc.regs[52][25] ;
 wire \top_ihp.oisc.regs[52][26] ;
 wire \top_ihp.oisc.regs[52][27] ;
 wire \top_ihp.oisc.regs[52][28] ;
 wire \top_ihp.oisc.regs[52][29] ;
 wire \top_ihp.oisc.regs[52][2] ;
 wire \top_ihp.oisc.regs[52][30] ;
 wire \top_ihp.oisc.regs[52][31] ;
 wire \top_ihp.oisc.regs[52][3] ;
 wire \top_ihp.oisc.regs[52][4] ;
 wire \top_ihp.oisc.regs[52][5] ;
 wire \top_ihp.oisc.regs[52][6] ;
 wire \top_ihp.oisc.regs[52][7] ;
 wire \top_ihp.oisc.regs[52][8] ;
 wire \top_ihp.oisc.regs[52][9] ;
 wire \top_ihp.oisc.regs[53][0] ;
 wire \top_ihp.oisc.regs[53][10] ;
 wire \top_ihp.oisc.regs[53][11] ;
 wire \top_ihp.oisc.regs[53][12] ;
 wire \top_ihp.oisc.regs[53][13] ;
 wire \top_ihp.oisc.regs[53][14] ;
 wire \top_ihp.oisc.regs[53][15] ;
 wire \top_ihp.oisc.regs[53][16] ;
 wire \top_ihp.oisc.regs[53][17] ;
 wire \top_ihp.oisc.regs[53][18] ;
 wire \top_ihp.oisc.regs[53][19] ;
 wire \top_ihp.oisc.regs[53][1] ;
 wire \top_ihp.oisc.regs[53][20] ;
 wire \top_ihp.oisc.regs[53][21] ;
 wire \top_ihp.oisc.regs[53][22] ;
 wire \top_ihp.oisc.regs[53][23] ;
 wire \top_ihp.oisc.regs[53][24] ;
 wire \top_ihp.oisc.regs[53][25] ;
 wire \top_ihp.oisc.regs[53][26] ;
 wire \top_ihp.oisc.regs[53][27] ;
 wire \top_ihp.oisc.regs[53][28] ;
 wire \top_ihp.oisc.regs[53][29] ;
 wire \top_ihp.oisc.regs[53][2] ;
 wire \top_ihp.oisc.regs[53][30] ;
 wire \top_ihp.oisc.regs[53][31] ;
 wire \top_ihp.oisc.regs[53][3] ;
 wire \top_ihp.oisc.regs[53][4] ;
 wire \top_ihp.oisc.regs[53][5] ;
 wire \top_ihp.oisc.regs[53][6] ;
 wire \top_ihp.oisc.regs[53][7] ;
 wire \top_ihp.oisc.regs[53][8] ;
 wire \top_ihp.oisc.regs[53][9] ;
 wire \top_ihp.oisc.regs[54][0] ;
 wire \top_ihp.oisc.regs[54][10] ;
 wire \top_ihp.oisc.regs[54][11] ;
 wire \top_ihp.oisc.regs[54][12] ;
 wire \top_ihp.oisc.regs[54][13] ;
 wire \top_ihp.oisc.regs[54][14] ;
 wire \top_ihp.oisc.regs[54][15] ;
 wire \top_ihp.oisc.regs[54][16] ;
 wire \top_ihp.oisc.regs[54][17] ;
 wire \top_ihp.oisc.regs[54][18] ;
 wire \top_ihp.oisc.regs[54][19] ;
 wire \top_ihp.oisc.regs[54][1] ;
 wire \top_ihp.oisc.regs[54][20] ;
 wire \top_ihp.oisc.regs[54][21] ;
 wire \top_ihp.oisc.regs[54][22] ;
 wire \top_ihp.oisc.regs[54][23] ;
 wire \top_ihp.oisc.regs[54][24] ;
 wire \top_ihp.oisc.regs[54][25] ;
 wire \top_ihp.oisc.regs[54][26] ;
 wire \top_ihp.oisc.regs[54][27] ;
 wire \top_ihp.oisc.regs[54][28] ;
 wire \top_ihp.oisc.regs[54][29] ;
 wire \top_ihp.oisc.regs[54][2] ;
 wire \top_ihp.oisc.regs[54][30] ;
 wire \top_ihp.oisc.regs[54][31] ;
 wire \top_ihp.oisc.regs[54][3] ;
 wire \top_ihp.oisc.regs[54][4] ;
 wire \top_ihp.oisc.regs[54][5] ;
 wire \top_ihp.oisc.regs[54][6] ;
 wire \top_ihp.oisc.regs[54][7] ;
 wire \top_ihp.oisc.regs[54][8] ;
 wire \top_ihp.oisc.regs[54][9] ;
 wire \top_ihp.oisc.regs[55][0] ;
 wire \top_ihp.oisc.regs[55][10] ;
 wire \top_ihp.oisc.regs[55][11] ;
 wire \top_ihp.oisc.regs[55][12] ;
 wire \top_ihp.oisc.regs[55][13] ;
 wire \top_ihp.oisc.regs[55][14] ;
 wire \top_ihp.oisc.regs[55][15] ;
 wire \top_ihp.oisc.regs[55][16] ;
 wire \top_ihp.oisc.regs[55][17] ;
 wire \top_ihp.oisc.regs[55][18] ;
 wire \top_ihp.oisc.regs[55][19] ;
 wire \top_ihp.oisc.regs[55][1] ;
 wire \top_ihp.oisc.regs[55][20] ;
 wire \top_ihp.oisc.regs[55][21] ;
 wire \top_ihp.oisc.regs[55][22] ;
 wire \top_ihp.oisc.regs[55][23] ;
 wire \top_ihp.oisc.regs[55][24] ;
 wire \top_ihp.oisc.regs[55][25] ;
 wire \top_ihp.oisc.regs[55][26] ;
 wire \top_ihp.oisc.regs[55][27] ;
 wire \top_ihp.oisc.regs[55][28] ;
 wire \top_ihp.oisc.regs[55][29] ;
 wire \top_ihp.oisc.regs[55][2] ;
 wire \top_ihp.oisc.regs[55][30] ;
 wire \top_ihp.oisc.regs[55][31] ;
 wire \top_ihp.oisc.regs[55][3] ;
 wire \top_ihp.oisc.regs[55][4] ;
 wire \top_ihp.oisc.regs[55][5] ;
 wire \top_ihp.oisc.regs[55][6] ;
 wire \top_ihp.oisc.regs[55][7] ;
 wire \top_ihp.oisc.regs[55][8] ;
 wire \top_ihp.oisc.regs[55][9] ;
 wire \top_ihp.oisc.regs[56][0] ;
 wire \top_ihp.oisc.regs[56][10] ;
 wire \top_ihp.oisc.regs[56][11] ;
 wire \top_ihp.oisc.regs[56][12] ;
 wire \top_ihp.oisc.regs[56][13] ;
 wire \top_ihp.oisc.regs[56][14] ;
 wire \top_ihp.oisc.regs[56][15] ;
 wire \top_ihp.oisc.regs[56][16] ;
 wire \top_ihp.oisc.regs[56][17] ;
 wire \top_ihp.oisc.regs[56][18] ;
 wire \top_ihp.oisc.regs[56][19] ;
 wire \top_ihp.oisc.regs[56][1] ;
 wire \top_ihp.oisc.regs[56][20] ;
 wire \top_ihp.oisc.regs[56][21] ;
 wire \top_ihp.oisc.regs[56][22] ;
 wire \top_ihp.oisc.regs[56][23] ;
 wire \top_ihp.oisc.regs[56][24] ;
 wire \top_ihp.oisc.regs[56][25] ;
 wire \top_ihp.oisc.regs[56][26] ;
 wire \top_ihp.oisc.regs[56][27] ;
 wire \top_ihp.oisc.regs[56][28] ;
 wire \top_ihp.oisc.regs[56][29] ;
 wire \top_ihp.oisc.regs[56][2] ;
 wire \top_ihp.oisc.regs[56][30] ;
 wire \top_ihp.oisc.regs[56][31] ;
 wire \top_ihp.oisc.regs[56][3] ;
 wire \top_ihp.oisc.regs[56][4] ;
 wire \top_ihp.oisc.regs[56][5] ;
 wire \top_ihp.oisc.regs[56][6] ;
 wire \top_ihp.oisc.regs[56][7] ;
 wire \top_ihp.oisc.regs[56][8] ;
 wire \top_ihp.oisc.regs[56][9] ;
 wire \top_ihp.oisc.regs[57][0] ;
 wire \top_ihp.oisc.regs[57][10] ;
 wire \top_ihp.oisc.regs[57][11] ;
 wire \top_ihp.oisc.regs[57][12] ;
 wire \top_ihp.oisc.regs[57][13] ;
 wire \top_ihp.oisc.regs[57][14] ;
 wire \top_ihp.oisc.regs[57][15] ;
 wire \top_ihp.oisc.regs[57][16] ;
 wire \top_ihp.oisc.regs[57][17] ;
 wire \top_ihp.oisc.regs[57][18] ;
 wire \top_ihp.oisc.regs[57][19] ;
 wire \top_ihp.oisc.regs[57][1] ;
 wire \top_ihp.oisc.regs[57][20] ;
 wire \top_ihp.oisc.regs[57][21] ;
 wire \top_ihp.oisc.regs[57][22] ;
 wire \top_ihp.oisc.regs[57][23] ;
 wire \top_ihp.oisc.regs[57][24] ;
 wire \top_ihp.oisc.regs[57][25] ;
 wire \top_ihp.oisc.regs[57][26] ;
 wire \top_ihp.oisc.regs[57][27] ;
 wire \top_ihp.oisc.regs[57][28] ;
 wire \top_ihp.oisc.regs[57][29] ;
 wire \top_ihp.oisc.regs[57][2] ;
 wire \top_ihp.oisc.regs[57][30] ;
 wire \top_ihp.oisc.regs[57][31] ;
 wire \top_ihp.oisc.regs[57][3] ;
 wire \top_ihp.oisc.regs[57][4] ;
 wire \top_ihp.oisc.regs[57][5] ;
 wire \top_ihp.oisc.regs[57][6] ;
 wire \top_ihp.oisc.regs[57][7] ;
 wire \top_ihp.oisc.regs[57][8] ;
 wire \top_ihp.oisc.regs[57][9] ;
 wire \top_ihp.oisc.regs[58][0] ;
 wire \top_ihp.oisc.regs[58][10] ;
 wire \top_ihp.oisc.regs[58][11] ;
 wire \top_ihp.oisc.regs[58][12] ;
 wire \top_ihp.oisc.regs[58][13] ;
 wire \top_ihp.oisc.regs[58][14] ;
 wire \top_ihp.oisc.regs[58][15] ;
 wire \top_ihp.oisc.regs[58][16] ;
 wire \top_ihp.oisc.regs[58][17] ;
 wire \top_ihp.oisc.regs[58][18] ;
 wire \top_ihp.oisc.regs[58][19] ;
 wire \top_ihp.oisc.regs[58][1] ;
 wire \top_ihp.oisc.regs[58][20] ;
 wire \top_ihp.oisc.regs[58][21] ;
 wire \top_ihp.oisc.regs[58][22] ;
 wire \top_ihp.oisc.regs[58][23] ;
 wire \top_ihp.oisc.regs[58][24] ;
 wire \top_ihp.oisc.regs[58][25] ;
 wire \top_ihp.oisc.regs[58][26] ;
 wire \top_ihp.oisc.regs[58][27] ;
 wire \top_ihp.oisc.regs[58][28] ;
 wire \top_ihp.oisc.regs[58][29] ;
 wire \top_ihp.oisc.regs[58][2] ;
 wire \top_ihp.oisc.regs[58][30] ;
 wire \top_ihp.oisc.regs[58][31] ;
 wire \top_ihp.oisc.regs[58][3] ;
 wire \top_ihp.oisc.regs[58][4] ;
 wire \top_ihp.oisc.regs[58][5] ;
 wire \top_ihp.oisc.regs[58][6] ;
 wire \top_ihp.oisc.regs[58][7] ;
 wire \top_ihp.oisc.regs[58][8] ;
 wire \top_ihp.oisc.regs[58][9] ;
 wire \top_ihp.oisc.regs[59][0] ;
 wire \top_ihp.oisc.regs[59][10] ;
 wire \top_ihp.oisc.regs[59][11] ;
 wire \top_ihp.oisc.regs[59][12] ;
 wire \top_ihp.oisc.regs[59][13] ;
 wire \top_ihp.oisc.regs[59][14] ;
 wire \top_ihp.oisc.regs[59][15] ;
 wire \top_ihp.oisc.regs[59][16] ;
 wire \top_ihp.oisc.regs[59][17] ;
 wire \top_ihp.oisc.regs[59][18] ;
 wire \top_ihp.oisc.regs[59][19] ;
 wire \top_ihp.oisc.regs[59][1] ;
 wire \top_ihp.oisc.regs[59][20] ;
 wire \top_ihp.oisc.regs[59][21] ;
 wire \top_ihp.oisc.regs[59][22] ;
 wire \top_ihp.oisc.regs[59][23] ;
 wire \top_ihp.oisc.regs[59][24] ;
 wire \top_ihp.oisc.regs[59][25] ;
 wire \top_ihp.oisc.regs[59][26] ;
 wire \top_ihp.oisc.regs[59][27] ;
 wire \top_ihp.oisc.regs[59][28] ;
 wire \top_ihp.oisc.regs[59][29] ;
 wire \top_ihp.oisc.regs[59][2] ;
 wire \top_ihp.oisc.regs[59][30] ;
 wire \top_ihp.oisc.regs[59][31] ;
 wire \top_ihp.oisc.regs[59][3] ;
 wire \top_ihp.oisc.regs[59][4] ;
 wire \top_ihp.oisc.regs[59][5] ;
 wire \top_ihp.oisc.regs[59][6] ;
 wire \top_ihp.oisc.regs[59][7] ;
 wire \top_ihp.oisc.regs[59][8] ;
 wire \top_ihp.oisc.regs[59][9] ;
 wire \top_ihp.oisc.regs[5][0] ;
 wire \top_ihp.oisc.regs[5][10] ;
 wire \top_ihp.oisc.regs[5][11] ;
 wire \top_ihp.oisc.regs[5][12] ;
 wire \top_ihp.oisc.regs[5][13] ;
 wire \top_ihp.oisc.regs[5][14] ;
 wire \top_ihp.oisc.regs[5][15] ;
 wire \top_ihp.oisc.regs[5][16] ;
 wire \top_ihp.oisc.regs[5][17] ;
 wire \top_ihp.oisc.regs[5][18] ;
 wire \top_ihp.oisc.regs[5][19] ;
 wire \top_ihp.oisc.regs[5][1] ;
 wire \top_ihp.oisc.regs[5][20] ;
 wire \top_ihp.oisc.regs[5][21] ;
 wire \top_ihp.oisc.regs[5][22] ;
 wire \top_ihp.oisc.regs[5][23] ;
 wire \top_ihp.oisc.regs[5][24] ;
 wire \top_ihp.oisc.regs[5][25] ;
 wire \top_ihp.oisc.regs[5][26] ;
 wire \top_ihp.oisc.regs[5][27] ;
 wire \top_ihp.oisc.regs[5][28] ;
 wire \top_ihp.oisc.regs[5][29] ;
 wire \top_ihp.oisc.regs[5][2] ;
 wire \top_ihp.oisc.regs[5][30] ;
 wire \top_ihp.oisc.regs[5][31] ;
 wire \top_ihp.oisc.regs[5][3] ;
 wire \top_ihp.oisc.regs[5][4] ;
 wire \top_ihp.oisc.regs[5][5] ;
 wire \top_ihp.oisc.regs[5][6] ;
 wire \top_ihp.oisc.regs[5][7] ;
 wire \top_ihp.oisc.regs[5][8] ;
 wire \top_ihp.oisc.regs[5][9] ;
 wire \top_ihp.oisc.regs[60][0] ;
 wire \top_ihp.oisc.regs[60][10] ;
 wire \top_ihp.oisc.regs[60][11] ;
 wire \top_ihp.oisc.regs[60][12] ;
 wire \top_ihp.oisc.regs[60][13] ;
 wire \top_ihp.oisc.regs[60][14] ;
 wire \top_ihp.oisc.regs[60][15] ;
 wire \top_ihp.oisc.regs[60][16] ;
 wire \top_ihp.oisc.regs[60][17] ;
 wire \top_ihp.oisc.regs[60][18] ;
 wire \top_ihp.oisc.regs[60][19] ;
 wire \top_ihp.oisc.regs[60][1] ;
 wire \top_ihp.oisc.regs[60][20] ;
 wire \top_ihp.oisc.regs[60][21] ;
 wire \top_ihp.oisc.regs[60][22] ;
 wire \top_ihp.oisc.regs[60][23] ;
 wire \top_ihp.oisc.regs[60][24] ;
 wire \top_ihp.oisc.regs[60][25] ;
 wire \top_ihp.oisc.regs[60][26] ;
 wire \top_ihp.oisc.regs[60][27] ;
 wire \top_ihp.oisc.regs[60][28] ;
 wire \top_ihp.oisc.regs[60][29] ;
 wire \top_ihp.oisc.regs[60][2] ;
 wire \top_ihp.oisc.regs[60][30] ;
 wire \top_ihp.oisc.regs[60][31] ;
 wire \top_ihp.oisc.regs[60][3] ;
 wire \top_ihp.oisc.regs[60][4] ;
 wire \top_ihp.oisc.regs[60][5] ;
 wire \top_ihp.oisc.regs[60][6] ;
 wire \top_ihp.oisc.regs[60][7] ;
 wire \top_ihp.oisc.regs[60][8] ;
 wire \top_ihp.oisc.regs[60][9] ;
 wire \top_ihp.oisc.regs[61][0] ;
 wire \top_ihp.oisc.regs[61][10] ;
 wire \top_ihp.oisc.regs[61][11] ;
 wire \top_ihp.oisc.regs[61][12] ;
 wire \top_ihp.oisc.regs[61][13] ;
 wire \top_ihp.oisc.regs[61][14] ;
 wire \top_ihp.oisc.regs[61][15] ;
 wire \top_ihp.oisc.regs[61][16] ;
 wire \top_ihp.oisc.regs[61][17] ;
 wire \top_ihp.oisc.regs[61][18] ;
 wire \top_ihp.oisc.regs[61][19] ;
 wire \top_ihp.oisc.regs[61][1] ;
 wire \top_ihp.oisc.regs[61][20] ;
 wire \top_ihp.oisc.regs[61][21] ;
 wire \top_ihp.oisc.regs[61][22] ;
 wire \top_ihp.oisc.regs[61][23] ;
 wire \top_ihp.oisc.regs[61][24] ;
 wire \top_ihp.oisc.regs[61][25] ;
 wire \top_ihp.oisc.regs[61][26] ;
 wire \top_ihp.oisc.regs[61][27] ;
 wire \top_ihp.oisc.regs[61][28] ;
 wire \top_ihp.oisc.regs[61][29] ;
 wire \top_ihp.oisc.regs[61][2] ;
 wire \top_ihp.oisc.regs[61][30] ;
 wire \top_ihp.oisc.regs[61][31] ;
 wire \top_ihp.oisc.regs[61][3] ;
 wire \top_ihp.oisc.regs[61][4] ;
 wire \top_ihp.oisc.regs[61][5] ;
 wire \top_ihp.oisc.regs[61][6] ;
 wire \top_ihp.oisc.regs[61][7] ;
 wire \top_ihp.oisc.regs[61][8] ;
 wire \top_ihp.oisc.regs[61][9] ;
 wire \top_ihp.oisc.regs[62][0] ;
 wire \top_ihp.oisc.regs[62][10] ;
 wire \top_ihp.oisc.regs[62][11] ;
 wire \top_ihp.oisc.regs[62][12] ;
 wire \top_ihp.oisc.regs[62][13] ;
 wire \top_ihp.oisc.regs[62][14] ;
 wire \top_ihp.oisc.regs[62][15] ;
 wire \top_ihp.oisc.regs[62][16] ;
 wire \top_ihp.oisc.regs[62][17] ;
 wire \top_ihp.oisc.regs[62][18] ;
 wire \top_ihp.oisc.regs[62][19] ;
 wire \top_ihp.oisc.regs[62][1] ;
 wire \top_ihp.oisc.regs[62][20] ;
 wire \top_ihp.oisc.regs[62][21] ;
 wire \top_ihp.oisc.regs[62][22] ;
 wire \top_ihp.oisc.regs[62][23] ;
 wire \top_ihp.oisc.regs[62][24] ;
 wire \top_ihp.oisc.regs[62][25] ;
 wire \top_ihp.oisc.regs[62][26] ;
 wire \top_ihp.oisc.regs[62][27] ;
 wire \top_ihp.oisc.regs[62][28] ;
 wire \top_ihp.oisc.regs[62][29] ;
 wire \top_ihp.oisc.regs[62][2] ;
 wire \top_ihp.oisc.regs[62][30] ;
 wire \top_ihp.oisc.regs[62][31] ;
 wire \top_ihp.oisc.regs[62][3] ;
 wire \top_ihp.oisc.regs[62][4] ;
 wire \top_ihp.oisc.regs[62][5] ;
 wire \top_ihp.oisc.regs[62][6] ;
 wire \top_ihp.oisc.regs[62][7] ;
 wire \top_ihp.oisc.regs[62][8] ;
 wire \top_ihp.oisc.regs[62][9] ;
 wire \top_ihp.oisc.regs[63][0] ;
 wire \top_ihp.oisc.regs[63][10] ;
 wire \top_ihp.oisc.regs[63][11] ;
 wire \top_ihp.oisc.regs[63][12] ;
 wire \top_ihp.oisc.regs[63][13] ;
 wire \top_ihp.oisc.regs[63][14] ;
 wire \top_ihp.oisc.regs[63][15] ;
 wire \top_ihp.oisc.regs[63][16] ;
 wire \top_ihp.oisc.regs[63][17] ;
 wire \top_ihp.oisc.regs[63][18] ;
 wire \top_ihp.oisc.regs[63][19] ;
 wire \top_ihp.oisc.regs[63][1] ;
 wire \top_ihp.oisc.regs[63][20] ;
 wire \top_ihp.oisc.regs[63][21] ;
 wire \top_ihp.oisc.regs[63][22] ;
 wire \top_ihp.oisc.regs[63][23] ;
 wire \top_ihp.oisc.regs[63][24] ;
 wire \top_ihp.oisc.regs[63][25] ;
 wire \top_ihp.oisc.regs[63][26] ;
 wire \top_ihp.oisc.regs[63][27] ;
 wire \top_ihp.oisc.regs[63][28] ;
 wire \top_ihp.oisc.regs[63][29] ;
 wire \top_ihp.oisc.regs[63][2] ;
 wire \top_ihp.oisc.regs[63][30] ;
 wire \top_ihp.oisc.regs[63][31] ;
 wire \top_ihp.oisc.regs[63][3] ;
 wire \top_ihp.oisc.regs[63][4] ;
 wire \top_ihp.oisc.regs[63][5] ;
 wire \top_ihp.oisc.regs[63][6] ;
 wire \top_ihp.oisc.regs[63][7] ;
 wire \top_ihp.oisc.regs[63][8] ;
 wire \top_ihp.oisc.regs[63][9] ;
 wire \top_ihp.oisc.regs[6][0] ;
 wire \top_ihp.oisc.regs[6][10] ;
 wire \top_ihp.oisc.regs[6][11] ;
 wire \top_ihp.oisc.regs[6][12] ;
 wire \top_ihp.oisc.regs[6][13] ;
 wire \top_ihp.oisc.regs[6][14] ;
 wire \top_ihp.oisc.regs[6][15] ;
 wire \top_ihp.oisc.regs[6][16] ;
 wire \top_ihp.oisc.regs[6][17] ;
 wire \top_ihp.oisc.regs[6][18] ;
 wire \top_ihp.oisc.regs[6][19] ;
 wire \top_ihp.oisc.regs[6][1] ;
 wire \top_ihp.oisc.regs[6][20] ;
 wire \top_ihp.oisc.regs[6][21] ;
 wire \top_ihp.oisc.regs[6][22] ;
 wire \top_ihp.oisc.regs[6][23] ;
 wire \top_ihp.oisc.regs[6][24] ;
 wire \top_ihp.oisc.regs[6][25] ;
 wire \top_ihp.oisc.regs[6][26] ;
 wire \top_ihp.oisc.regs[6][27] ;
 wire \top_ihp.oisc.regs[6][28] ;
 wire \top_ihp.oisc.regs[6][29] ;
 wire \top_ihp.oisc.regs[6][2] ;
 wire \top_ihp.oisc.regs[6][30] ;
 wire \top_ihp.oisc.regs[6][31] ;
 wire \top_ihp.oisc.regs[6][3] ;
 wire \top_ihp.oisc.regs[6][4] ;
 wire \top_ihp.oisc.regs[6][5] ;
 wire \top_ihp.oisc.regs[6][6] ;
 wire \top_ihp.oisc.regs[6][7] ;
 wire \top_ihp.oisc.regs[6][8] ;
 wire \top_ihp.oisc.regs[6][9] ;
 wire \top_ihp.oisc.regs[7][0] ;
 wire \top_ihp.oisc.regs[7][10] ;
 wire \top_ihp.oisc.regs[7][11] ;
 wire \top_ihp.oisc.regs[7][12] ;
 wire \top_ihp.oisc.regs[7][13] ;
 wire \top_ihp.oisc.regs[7][14] ;
 wire \top_ihp.oisc.regs[7][15] ;
 wire \top_ihp.oisc.regs[7][16] ;
 wire \top_ihp.oisc.regs[7][17] ;
 wire \top_ihp.oisc.regs[7][18] ;
 wire \top_ihp.oisc.regs[7][19] ;
 wire \top_ihp.oisc.regs[7][1] ;
 wire \top_ihp.oisc.regs[7][20] ;
 wire \top_ihp.oisc.regs[7][21] ;
 wire \top_ihp.oisc.regs[7][22] ;
 wire \top_ihp.oisc.regs[7][23] ;
 wire \top_ihp.oisc.regs[7][24] ;
 wire \top_ihp.oisc.regs[7][25] ;
 wire \top_ihp.oisc.regs[7][26] ;
 wire \top_ihp.oisc.regs[7][27] ;
 wire \top_ihp.oisc.regs[7][28] ;
 wire \top_ihp.oisc.regs[7][29] ;
 wire \top_ihp.oisc.regs[7][2] ;
 wire \top_ihp.oisc.regs[7][30] ;
 wire \top_ihp.oisc.regs[7][31] ;
 wire \top_ihp.oisc.regs[7][3] ;
 wire \top_ihp.oisc.regs[7][4] ;
 wire \top_ihp.oisc.regs[7][5] ;
 wire \top_ihp.oisc.regs[7][6] ;
 wire \top_ihp.oisc.regs[7][7] ;
 wire \top_ihp.oisc.regs[7][8] ;
 wire \top_ihp.oisc.regs[7][9] ;
 wire \top_ihp.oisc.regs[8][0] ;
 wire \top_ihp.oisc.regs[8][10] ;
 wire \top_ihp.oisc.regs[8][11] ;
 wire \top_ihp.oisc.regs[8][12] ;
 wire \top_ihp.oisc.regs[8][13] ;
 wire \top_ihp.oisc.regs[8][14] ;
 wire \top_ihp.oisc.regs[8][15] ;
 wire \top_ihp.oisc.regs[8][16] ;
 wire \top_ihp.oisc.regs[8][17] ;
 wire \top_ihp.oisc.regs[8][18] ;
 wire \top_ihp.oisc.regs[8][19] ;
 wire \top_ihp.oisc.regs[8][1] ;
 wire \top_ihp.oisc.regs[8][20] ;
 wire \top_ihp.oisc.regs[8][21] ;
 wire \top_ihp.oisc.regs[8][22] ;
 wire \top_ihp.oisc.regs[8][23] ;
 wire \top_ihp.oisc.regs[8][24] ;
 wire \top_ihp.oisc.regs[8][25] ;
 wire \top_ihp.oisc.regs[8][26] ;
 wire \top_ihp.oisc.regs[8][27] ;
 wire \top_ihp.oisc.regs[8][28] ;
 wire \top_ihp.oisc.regs[8][29] ;
 wire \top_ihp.oisc.regs[8][2] ;
 wire \top_ihp.oisc.regs[8][30] ;
 wire \top_ihp.oisc.regs[8][31] ;
 wire \top_ihp.oisc.regs[8][3] ;
 wire \top_ihp.oisc.regs[8][4] ;
 wire \top_ihp.oisc.regs[8][5] ;
 wire \top_ihp.oisc.regs[8][6] ;
 wire \top_ihp.oisc.regs[8][7] ;
 wire \top_ihp.oisc.regs[8][8] ;
 wire \top_ihp.oisc.regs[8][9] ;
 wire \top_ihp.oisc.regs[9][0] ;
 wire \top_ihp.oisc.regs[9][10] ;
 wire \top_ihp.oisc.regs[9][11] ;
 wire \top_ihp.oisc.regs[9][12] ;
 wire \top_ihp.oisc.regs[9][13] ;
 wire \top_ihp.oisc.regs[9][14] ;
 wire \top_ihp.oisc.regs[9][15] ;
 wire \top_ihp.oisc.regs[9][16] ;
 wire \top_ihp.oisc.regs[9][17] ;
 wire \top_ihp.oisc.regs[9][18] ;
 wire \top_ihp.oisc.regs[9][19] ;
 wire \top_ihp.oisc.regs[9][1] ;
 wire \top_ihp.oisc.regs[9][20] ;
 wire \top_ihp.oisc.regs[9][21] ;
 wire \top_ihp.oisc.regs[9][22] ;
 wire \top_ihp.oisc.regs[9][23] ;
 wire \top_ihp.oisc.regs[9][24] ;
 wire \top_ihp.oisc.regs[9][25] ;
 wire \top_ihp.oisc.regs[9][26] ;
 wire \top_ihp.oisc.regs[9][27] ;
 wire \top_ihp.oisc.regs[9][28] ;
 wire \top_ihp.oisc.regs[9][29] ;
 wire \top_ihp.oisc.regs[9][2] ;
 wire \top_ihp.oisc.regs[9][30] ;
 wire \top_ihp.oisc.regs[9][31] ;
 wire \top_ihp.oisc.regs[9][3] ;
 wire \top_ihp.oisc.regs[9][4] ;
 wire \top_ihp.oisc.regs[9][5] ;
 wire \top_ihp.oisc.regs[9][6] ;
 wire \top_ihp.oisc.regs[9][7] ;
 wire \top_ihp.oisc.regs[9][8] ;
 wire \top_ihp.oisc.regs[9][9] ;
 wire \top_ihp.oisc.state[0] ;
 wire \top_ihp.oisc.state[1] ;
 wire \top_ihp.oisc.state[2] ;
 wire \top_ihp.oisc.state[3] ;
 wire \top_ihp.oisc.state[4] ;
 wire \top_ihp.oisc.state[5] ;
 wire \top_ihp.oisc.state[6] ;
 wire \top_ihp.oisc.wb_adr_o[0] ;
 wire \top_ihp.oisc.wb_adr_o[1] ;
 wire \top_ihp.oisc.wb_dat_o[0] ;
 wire \top_ihp.oisc.wb_dat_o[10] ;
 wire \top_ihp.oisc.wb_dat_o[11] ;
 wire \top_ihp.oisc.wb_dat_o[12] ;
 wire \top_ihp.oisc.wb_dat_o[13] ;
 wire \top_ihp.oisc.wb_dat_o[14] ;
 wire \top_ihp.oisc.wb_dat_o[15] ;
 wire \top_ihp.oisc.wb_dat_o[16] ;
 wire \top_ihp.oisc.wb_dat_o[17] ;
 wire \top_ihp.oisc.wb_dat_o[18] ;
 wire \top_ihp.oisc.wb_dat_o[19] ;
 wire \top_ihp.oisc.wb_dat_o[1] ;
 wire \top_ihp.oisc.wb_dat_o[20] ;
 wire \top_ihp.oisc.wb_dat_o[21] ;
 wire \top_ihp.oisc.wb_dat_o[22] ;
 wire \top_ihp.oisc.wb_dat_o[23] ;
 wire \top_ihp.oisc.wb_dat_o[24] ;
 wire \top_ihp.oisc.wb_dat_o[25] ;
 wire \top_ihp.oisc.wb_dat_o[26] ;
 wire \top_ihp.oisc.wb_dat_o[27] ;
 wire \top_ihp.oisc.wb_dat_o[28] ;
 wire \top_ihp.oisc.wb_dat_o[29] ;
 wire \top_ihp.oisc.wb_dat_o[2] ;
 wire \top_ihp.oisc.wb_dat_o[30] ;
 wire \top_ihp.oisc.wb_dat_o[31] ;
 wire \top_ihp.oisc.wb_dat_o[3] ;
 wire \top_ihp.oisc.wb_dat_o[4] ;
 wire \top_ihp.oisc.wb_dat_o[5] ;
 wire \top_ihp.oisc.wb_dat_o[6] ;
 wire \top_ihp.oisc.wb_dat_o[7] ;
 wire \top_ihp.oisc.wb_dat_o[8] ;
 wire \top_ihp.oisc.wb_dat_o[9] ;
 wire \top_ihp.ram_clk_o ;
 wire \top_ihp.ram_cs_o ;
 wire \top_ihp.ram_data_o ;
 wire \top_ihp.rom_clk_o ;
 wire \top_ihp.rom_cs_o ;
 wire \top_ihp.rom_data_o ;
 wire \top_ihp.spi_clk_o ;
 wire \top_ihp.spi_cs_o_1 ;
 wire \top_ihp.spi_cs_o_2 ;
 wire \top_ihp.spi_cs_o_3 ;
 wire \top_ihp.spi_data_o ;
 wire \top_ihp.tx ;
 wire \top_ihp.wb_ack_gpio ;
 wire \top_ihp.wb_ack_spi ;
 wire \top_ihp.wb_ack_uart ;
 wire \top_ihp.wb_dati_gpio[0] ;
 wire \top_ihp.wb_dati_ram[0] ;
 wire \top_ihp.wb_dati_ram[10] ;
 wire \top_ihp.wb_dati_ram[11] ;
 wire \top_ihp.wb_dati_ram[12] ;
 wire \top_ihp.wb_dati_ram[13] ;
 wire \top_ihp.wb_dati_ram[14] ;
 wire \top_ihp.wb_dati_ram[15] ;
 wire \top_ihp.wb_dati_ram[16] ;
 wire \top_ihp.wb_dati_ram[17] ;
 wire \top_ihp.wb_dati_ram[18] ;
 wire \top_ihp.wb_dati_ram[19] ;
 wire \top_ihp.wb_dati_ram[1] ;
 wire \top_ihp.wb_dati_ram[20] ;
 wire \top_ihp.wb_dati_ram[21] ;
 wire \top_ihp.wb_dati_ram[22] ;
 wire \top_ihp.wb_dati_ram[23] ;
 wire \top_ihp.wb_dati_ram[24] ;
 wire \top_ihp.wb_dati_ram[25] ;
 wire \top_ihp.wb_dati_ram[26] ;
 wire \top_ihp.wb_dati_ram[27] ;
 wire \top_ihp.wb_dati_ram[28] ;
 wire \top_ihp.wb_dati_ram[29] ;
 wire \top_ihp.wb_dati_ram[2] ;
 wire \top_ihp.wb_dati_ram[30] ;
 wire \top_ihp.wb_dati_ram[31] ;
 wire \top_ihp.wb_dati_ram[3] ;
 wire \top_ihp.wb_dati_ram[4] ;
 wire \top_ihp.wb_dati_ram[5] ;
 wire \top_ihp.wb_dati_ram[6] ;
 wire \top_ihp.wb_dati_ram[7] ;
 wire \top_ihp.wb_dati_ram[8] ;
 wire \top_ihp.wb_dati_ram[9] ;
 wire \top_ihp.wb_dati_rom[0] ;
 wire \top_ihp.wb_dati_rom[10] ;
 wire \top_ihp.wb_dati_rom[11] ;
 wire \top_ihp.wb_dati_rom[12] ;
 wire \top_ihp.wb_dati_rom[13] ;
 wire \top_ihp.wb_dati_rom[14] ;
 wire \top_ihp.wb_dati_rom[15] ;
 wire \top_ihp.wb_dati_rom[16] ;
 wire \top_ihp.wb_dati_rom[17] ;
 wire \top_ihp.wb_dati_rom[18] ;
 wire \top_ihp.wb_dati_rom[19] ;
 wire \top_ihp.wb_dati_rom[1] ;
 wire \top_ihp.wb_dati_rom[20] ;
 wire \top_ihp.wb_dati_rom[21] ;
 wire \top_ihp.wb_dati_rom[22] ;
 wire \top_ihp.wb_dati_rom[23] ;
 wire \top_ihp.wb_dati_rom[24] ;
 wire \top_ihp.wb_dati_rom[25] ;
 wire \top_ihp.wb_dati_rom[26] ;
 wire \top_ihp.wb_dati_rom[27] ;
 wire \top_ihp.wb_dati_rom[28] ;
 wire \top_ihp.wb_dati_rom[29] ;
 wire \top_ihp.wb_dati_rom[2] ;
 wire \top_ihp.wb_dati_rom[30] ;
 wire \top_ihp.wb_dati_rom[31] ;
 wire \top_ihp.wb_dati_rom[3] ;
 wire \top_ihp.wb_dati_rom[4] ;
 wire \top_ihp.wb_dati_rom[5] ;
 wire \top_ihp.wb_dati_rom[6] ;
 wire \top_ihp.wb_dati_rom[7] ;
 wire \top_ihp.wb_dati_rom[8] ;
 wire \top_ihp.wb_dati_rom[9] ;
 wire \top_ihp.wb_dati_spi[0] ;
 wire \top_ihp.wb_dati_spi[10] ;
 wire \top_ihp.wb_dati_spi[11] ;
 wire \top_ihp.wb_dati_spi[12] ;
 wire \top_ihp.wb_dati_spi[13] ;
 wire \top_ihp.wb_dati_spi[14] ;
 wire \top_ihp.wb_dati_spi[15] ;
 wire \top_ihp.wb_dati_spi[16] ;
 wire \top_ihp.wb_dati_spi[17] ;
 wire \top_ihp.wb_dati_spi[18] ;
 wire \top_ihp.wb_dati_spi[19] ;
 wire \top_ihp.wb_dati_spi[1] ;
 wire \top_ihp.wb_dati_spi[20] ;
 wire \top_ihp.wb_dati_spi[21] ;
 wire \top_ihp.wb_dati_spi[22] ;
 wire \top_ihp.wb_dati_spi[23] ;
 wire \top_ihp.wb_dati_spi[24] ;
 wire \top_ihp.wb_dati_spi[25] ;
 wire \top_ihp.wb_dati_spi[26] ;
 wire \top_ihp.wb_dati_spi[27] ;
 wire \top_ihp.wb_dati_spi[28] ;
 wire \top_ihp.wb_dati_spi[29] ;
 wire \top_ihp.wb_dati_spi[2] ;
 wire \top_ihp.wb_dati_spi[30] ;
 wire \top_ihp.wb_dati_spi[31] ;
 wire \top_ihp.wb_dati_spi[3] ;
 wire \top_ihp.wb_dati_spi[4] ;
 wire \top_ihp.wb_dati_spi[5] ;
 wire \top_ihp.wb_dati_spi[6] ;
 wire \top_ihp.wb_dati_spi[7] ;
 wire \top_ihp.wb_dati_spi[8] ;
 wire \top_ihp.wb_dati_spi[9] ;
 wire \top_ihp.wb_dati_uart[0] ;
 wire \top_ihp.wb_dati_uart[1] ;
 wire \top_ihp.wb_dati_uart[2] ;
 wire \top_ihp.wb_dati_uart[3] ;
 wire \top_ihp.wb_dati_uart[4] ;
 wire \top_ihp.wb_dati_uart[5] ;
 wire \top_ihp.wb_dati_uart[6] ;
 wire \top_ihp.wb_dati_uart[7] ;
 wire \top_ihp.wb_emem.bit_counter[0] ;
 wire \top_ihp.wb_emem.bit_counter[1] ;
 wire \top_ihp.wb_emem.bit_counter[2] ;
 wire \top_ihp.wb_emem.bit_counter[3] ;
 wire \top_ihp.wb_emem.bit_counter[4] ;
 wire \top_ihp.wb_emem.bit_counter[5] ;
 wire \top_ihp.wb_emem.bit_counter[6] ;
 wire \top_ihp.wb_emem.bit_counter[7] ;
 wire \top_ihp.wb_emem.cmd[32] ;
 wire \top_ihp.wb_emem.cmd[33] ;
 wire \top_ihp.wb_emem.cmd[34] ;
 wire \top_ihp.wb_emem.cmd[35] ;
 wire \top_ihp.wb_emem.cmd[36] ;
 wire \top_ihp.wb_emem.cmd[37] ;
 wire \top_ihp.wb_emem.cmd[38] ;
 wire \top_ihp.wb_emem.cmd[39] ;
 wire \top_ihp.wb_emem.cmd[40] ;
 wire \top_ihp.wb_emem.cmd[41] ;
 wire \top_ihp.wb_emem.cmd[42] ;
 wire \top_ihp.wb_emem.cmd[43] ;
 wire \top_ihp.wb_emem.cmd[44] ;
 wire \top_ihp.wb_emem.cmd[45] ;
 wire \top_ihp.wb_emem.cmd[46] ;
 wire \top_ihp.wb_emem.cmd[47] ;
 wire \top_ihp.wb_emem.cmd[48] ;
 wire \top_ihp.wb_emem.cmd[49] ;
 wire \top_ihp.wb_emem.cmd[50] ;
 wire \top_ihp.wb_emem.cmd[51] ;
 wire \top_ihp.wb_emem.cmd[52] ;
 wire \top_ihp.wb_emem.cmd[53] ;
 wire \top_ihp.wb_emem.cmd[54] ;
 wire \top_ihp.wb_emem.cmd[55] ;
 wire \top_ihp.wb_emem.cmd[56] ;
 wire \top_ihp.wb_emem.cmd[57] ;
 wire \top_ihp.wb_emem.cmd[58] ;
 wire \top_ihp.wb_emem.cmd[59] ;
 wire \top_ihp.wb_emem.cmd[60] ;
 wire \top_ihp.wb_emem.cmd[61] ;
 wire \top_ihp.wb_emem.cmd[62] ;
 wire \top_ihp.wb_emem.cmd[63] ;
 wire \top_ihp.wb_emem.last_bit ;
 wire \top_ihp.wb_emem.last_wait ;
 wire \top_ihp.wb_emem.nbits[3] ;
 wire \top_ihp.wb_emem.nbits[4] ;
 wire \top_ihp.wb_emem.nbits[5] ;
 wire \top_ihp.wb_emem.nbits[6] ;
 wire \top_ihp.wb_emem.state[0] ;
 wire \top_ihp.wb_emem.state[1] ;
 wire \top_ihp.wb_emem.state[2] ;
 wire \top_ihp.wb_emem.state[3] ;
 wire \top_ihp.wb_emem.wait_counter[0] ;
 wire \top_ihp.wb_emem.wait_counter[1] ;
 wire \top_ihp.wb_emem.wait_counter[2] ;
 wire \top_ihp.wb_emem.wait_counter[3] ;
 wire \top_ihp.wb_emem.wait_counter[4] ;
 wire \top_ihp.wb_emem.wait_counter[5] ;
 wire \top_ihp.wb_emem.wait_counter[6] ;
 wire \top_ihp.wb_emem.wait_counter[7] ;
 wire \top_ihp.wb_imem.bits_left[0] ;
 wire \top_ihp.wb_imem.bits_left[1] ;
 wire \top_ihp.wb_imem.bits_left[2] ;
 wire \top_ihp.wb_imem.bits_left[3] ;
 wire \top_ihp.wb_imem.bits_left[4] ;
 wire \top_ihp.wb_imem.bits_left[5] ;
 wire \top_ihp.wb_imem.state[0] ;
 wire \top_ihp.wb_imem.state[1] ;
 wire \top_ihp.wb_imem.state[2] ;
 wire \top_ihp.wb_spi.bits_left[0] ;
 wire \top_ihp.wb_spi.bits_left[1] ;
 wire \top_ihp.wb_spi.bits_left[2] ;
 wire \top_ihp.wb_spi.bits_left[3] ;
 wire \top_ihp.wb_spi.bits_left[4] ;
 wire \top_ihp.wb_spi.bits_left[5] ;
 wire \top_ihp.wb_spi.spi_clk_cnt[0] ;
 wire \top_ihp.wb_spi.state ;
 wire \top_ihp.wb_uart.rx_ready ;
 wire \top_ihp.wb_uart.state[0] ;
 wire \top_ihp.wb_uart.state[1] ;
 wire \top_ihp.wb_uart.tx_ready ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[0] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[1] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[2] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[3] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[0] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[10] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[11] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[12] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[13] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[14] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[15] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[16] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[17] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[18] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[19] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[1] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[20] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[21] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[22] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[23] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[24] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[25] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[26] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[27] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[28] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[29] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[2] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[30] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[31] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[3] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[4] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[5] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[6] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[7] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[8] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[9] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[0] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[1] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[2] ;
 wire \top_ihp.wb_uart.uart_rx.state[0] ;
 wire \top_ihp.wb_uart.uart_rx.state[1] ;
 wire \top_ihp.wb_uart.uart_rx.state[2] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[0] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[1] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[2] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[3] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[0] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[10] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[11] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[12] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[13] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[14] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[15] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[16] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[17] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[18] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[19] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[1] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[20] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[21] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[22] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[23] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[24] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[25] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[26] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[27] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[28] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[29] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[2] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[30] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[31] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[3] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[4] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[5] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[6] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[7] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[8] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[9] ;
 wire \top_ihp.wb_uart.uart_tx.next_state[0] ;
 wire \top_ihp.wb_uart.uart_tx.next_state[1] ;
 wire \top_ihp.wb_uart.uart_tx.state[0] ;
 wire \top_ihp.wb_uart.uart_tx.state[1] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[0] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[1] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[2] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[3] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[4] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[5] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[6] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _13211_ (.A(\top_ihp.oisc.state[1] ),
    .X(_07417_));
 sg13g2_buf_1 _13212_ (.A(_07417_),
    .X(_07418_));
 sg13g2_buf_1 _13213_ (.A(\top_ihp.oisc.decoder.decoded[10] ),
    .X(_07419_));
 sg13g2_buf_1 _13214_ (.A(\top_ihp.oisc.decoder.decoded[11] ),
    .X(_07420_));
 sg13g2_nor2_1 _13215_ (.A(_07419_),
    .B(_07420_),
    .Y(_07421_));
 sg13g2_buf_1 _13216_ (.A(\top_ihp.oisc.state[5] ),
    .X(_07422_));
 sg13g2_buf_1 _13217_ (.A(_07422_),
    .X(_07423_));
 sg13g2_buf_2 _13218_ (.A(\top_ihp.oisc.micro_op[1] ),
    .X(_07424_));
 sg13g2_buf_2 _13219_ (.A(\top_ihp.oisc.micro_op[0] ),
    .X(_07425_));
 sg13g2_buf_2 _13220_ (.A(\top_ihp.oisc.micro_op[4] ),
    .X(_07426_));
 sg13g2_and4_1 _13221_ (.A(_07424_),
    .B(_07425_),
    .C(_07426_),
    .D(\top_ihp.oisc.micro_state[2] ),
    .X(_07427_));
 sg13g2_buf_1 _13222_ (.A(_07427_),
    .X(_07428_));
 sg13g2_buf_2 _13223_ (.A(\top_ihp.oisc.micro_op[3] ),
    .X(_07429_));
 sg13g2_buf_2 _13224_ (.A(\top_ihp.oisc.micro_op[2] ),
    .X(_07430_));
 sg13g2_buf_1 _13225_ (.A(\top_ihp.oisc.micro_op[5] ),
    .X(_07431_));
 sg13g2_and3_1 _13226_ (.X(_07432_),
    .A(_07429_),
    .B(_07430_),
    .C(_07431_));
 sg13g2_buf_1 _13227_ (.A(_07432_),
    .X(_07433_));
 sg13g2_and2_1 _13228_ (.A(_07428_),
    .B(_07433_),
    .X(_07434_));
 sg13g2_buf_1 _13229_ (.A(_07434_),
    .X(_07435_));
 sg13g2_buf_8 _13230_ (.A(_07435_),
    .X(_07436_));
 sg13g2_and2_1 _13231_ (.A(net1016),
    .B(net879),
    .X(_07437_));
 sg13g2_nand2b_1 _13232_ (.Y(_07438_),
    .B(_07437_),
    .A_N(_07421_));
 sg13g2_nor2_1 _13233_ (.A(net1017),
    .B(_07438_),
    .Y(_07439_));
 sg13g2_buf_1 _13234_ (.A(_07439_),
    .X(_07440_));
 sg13g2_buf_1 _13235_ (.A(net807),
    .X(_07441_));
 sg13g2_buf_2 _13236_ (.A(\top_ihp.oisc.op_a[23] ),
    .X(_07442_));
 sg13g2_buf_1 _13237_ (.A(\top_ihp.oisc.op_b[23] ),
    .X(_07443_));
 sg13g2_buf_2 _13238_ (.A(\top_ihp.oisc.op_a[22] ),
    .X(_07444_));
 sg13g2_buf_1 _13239_ (.A(\top_ihp.oisc.op_b[22] ),
    .X(_07445_));
 sg13g2_nor2b_1 _13240_ (.A(_07444_),
    .B_N(net1044),
    .Y(_07446_));
 sg13g2_nor2_1 _13241_ (.A(_07443_),
    .B(_07446_),
    .Y(_07447_));
 sg13g2_nand2_1 _13242_ (.Y(_07448_),
    .A(_07443_),
    .B(_07446_));
 sg13g2_o21ai_1 _13243_ (.B1(_07448_),
    .Y(_07449_),
    .A1(_07442_),
    .A2(_07447_));
 sg13g2_buf_2 _13244_ (.A(\top_ihp.oisc.op_a[20] ),
    .X(_07450_));
 sg13g2_inv_1 _13245_ (.Y(_07451_),
    .A(_07450_));
 sg13g2_buf_2 _13246_ (.A(\top_ihp.oisc.op_b[20] ),
    .X(_07452_));
 sg13g2_buf_1 _13247_ (.A(\top_ihp.oisc.op_b[19] ),
    .X(_07453_));
 sg13g2_inv_1 _13248_ (.Y(_07454_),
    .A(_07453_));
 sg13g2_buf_2 _13249_ (.A(\top_ihp.oisc.op_a[18] ),
    .X(_07455_));
 sg13g2_buf_1 _13250_ (.A(\top_ihp.oisc.op_b[18] ),
    .X(_07456_));
 sg13g2_nand2b_1 _13251_ (.Y(_07457_),
    .B(_07456_),
    .A_N(net1043));
 sg13g2_nand2_1 _13252_ (.Y(_07458_),
    .A(_07454_),
    .B(_07457_));
 sg13g2_buf_1 _13253_ (.A(\top_ihp.oisc.op_a[19] ),
    .X(_07459_));
 sg13g2_o21ai_1 _13254_ (.B1(net1042),
    .Y(_07460_),
    .A1(_07454_),
    .A2(_07457_));
 sg13g2_buf_2 _13255_ (.A(\top_ihp.oisc.op_a[21] ),
    .X(_07461_));
 sg13g2_buf_1 _13256_ (.A(\top_ihp.oisc.op_b[21] ),
    .X(_07462_));
 sg13g2_nor2b_1 _13257_ (.A(_07461_),
    .B_N(_07462_),
    .Y(_07463_));
 sg13g2_buf_2 _13258_ (.A(_07463_),
    .X(_07464_));
 sg13g2_a221oi_1 _13259_ (.B2(_07460_),
    .C1(_07464_),
    .B1(_07458_),
    .A1(_07451_),
    .Y(_07465_),
    .A2(_07452_));
 sg13g2_nand2b_1 _13260_ (.Y(_07466_),
    .B(_07450_),
    .A_N(_07452_));
 sg13g2_nand2b_1 _13261_ (.Y(_07467_),
    .B(_07461_),
    .A_N(_07462_));
 sg13g2_o21ai_1 _13262_ (.B1(_07467_),
    .Y(_07468_),
    .A1(_07464_),
    .A2(_07466_));
 sg13g2_or2_1 _13263_ (.X(_07469_),
    .B(_07468_),
    .A(_07465_));
 sg13g2_buf_1 _13264_ (.A(_07469_),
    .X(_07470_));
 sg13g2_nand2b_1 _13265_ (.Y(_07471_),
    .B(_07470_),
    .A_N(_07449_));
 sg13g2_buf_1 _13266_ (.A(\top_ihp.oisc.op_b[2] ),
    .X(_07472_));
 sg13g2_nor2b_1 _13267_ (.A(_07472_),
    .B_N(\top_ihp.oisc.op_a[2] ),
    .Y(_07473_));
 sg13g2_buf_2 _13268_ (.A(\top_ihp.oisc.op_b[0] ),
    .X(_07474_));
 sg13g2_buf_8 _13269_ (.A(\top_ihp.oisc.op_a[0] ),
    .X(_07475_));
 sg13g2_nand2b_1 _13270_ (.Y(_07476_),
    .B(_07475_),
    .A_N(_07474_));
 sg13g2_buf_1 _13271_ (.A(\top_ihp.oisc.op_b[1] ),
    .X(_07477_));
 sg13g2_buf_1 _13272_ (.A(\top_ihp.oisc.op_a[1] ),
    .X(_07478_));
 sg13g2_nand2b_1 _13273_ (.Y(_07479_),
    .B(net1041),
    .A_N(_07477_));
 sg13g2_nor2b_1 _13274_ (.A(net1041),
    .B_N(_07477_),
    .Y(_07480_));
 sg13g2_a21oi_2 _13275_ (.B1(_07480_),
    .Y(_07481_),
    .A2(_07479_),
    .A1(_07476_));
 sg13g2_buf_1 _13276_ (.A(\top_ihp.oisc.op_a[2] ),
    .X(_07482_));
 sg13g2_nand2b_1 _13277_ (.Y(_07483_),
    .B(_07472_),
    .A_N(net1040));
 sg13g2_o21ai_1 _13278_ (.B1(_07483_),
    .Y(_07484_),
    .A1(_07473_),
    .A2(_07481_));
 sg13g2_buf_2 _13279_ (.A(\top_ihp.oisc.op_b[3] ),
    .X(_07485_));
 sg13g2_buf_1 _13280_ (.A(\top_ihp.oisc.op_b[4] ),
    .X(_07486_));
 sg13g2_buf_1 _13281_ (.A(\top_ihp.oisc.op_a[4] ),
    .X(_07487_));
 sg13g2_nand2b_1 _13282_ (.Y(_07488_),
    .B(net1039),
    .A_N(_07486_));
 sg13g2_buf_1 _13283_ (.A(\top_ihp.oisc.op_b[5] ),
    .X(_07489_));
 sg13g2_buf_2 _13284_ (.A(\top_ihp.oisc.op_a[5] ),
    .X(_07490_));
 sg13g2_nand2b_1 _13285_ (.Y(_07491_),
    .B(net1038),
    .A_N(_07489_));
 sg13g2_and3_1 _13286_ (.X(_07492_),
    .A(_07485_),
    .B(_07488_),
    .C(_07491_));
 sg13g2_nor2b_1 _13287_ (.A(net1040),
    .B_N(_07472_),
    .Y(_07493_));
 sg13g2_nor2_1 _13288_ (.A(_07485_),
    .B(_07493_),
    .Y(_07494_));
 sg13g2_o21ai_1 _13289_ (.B1(_07494_),
    .Y(_07495_),
    .A1(_07473_),
    .A2(_07481_));
 sg13g2_buf_2 _13290_ (.A(\top_ihp.oisc.op_a[3] ),
    .X(_07496_));
 sg13g2_nand2b_1 _13291_ (.Y(_07497_),
    .B(_07486_),
    .A_N(net1039));
 sg13g2_nand2b_1 _13292_ (.Y(_07498_),
    .B(_07489_),
    .A_N(net1038));
 sg13g2_nand4_1 _13293_ (.B(_07491_),
    .C(_07497_),
    .A(_07488_),
    .Y(_07499_),
    .D(_07498_));
 sg13g2_nor2_1 _13294_ (.A(net1037),
    .B(_07499_),
    .Y(_07500_));
 sg13g2_nor2b_1 _13295_ (.A(net1039),
    .B_N(_07486_),
    .Y(_07501_));
 sg13g2_inv_1 _13296_ (.Y(_07502_),
    .A(_07489_));
 sg13g2_a21oi_1 _13297_ (.A1(_07502_),
    .A2(_07497_),
    .Y(_07503_),
    .B1(net1038));
 sg13g2_a21o_1 _13298_ (.A2(_07501_),
    .A1(_07489_),
    .B1(_07503_),
    .X(_07504_));
 sg13g2_a221oi_1 _13299_ (.B2(_07500_),
    .C1(_07504_),
    .B1(_07495_),
    .A1(_07484_),
    .Y(_07505_),
    .A2(_07492_));
 sg13g2_buf_2 _13300_ (.A(_07505_),
    .X(_07506_));
 sg13g2_buf_2 _13301_ (.A(\top_ihp.oisc.op_a[16] ),
    .X(_07507_));
 sg13g2_buf_2 _13302_ (.A(\top_ihp.oisc.op_b[16] ),
    .X(_07508_));
 sg13g2_xnor2_1 _13303_ (.Y(_07509_),
    .A(_07507_),
    .B(_07508_));
 sg13g2_buf_1 _13304_ (.A(\top_ihp.oisc.op_a[15] ),
    .X(_07510_));
 sg13g2_buf_1 _13305_ (.A(\top_ihp.oisc.op_b[15] ),
    .X(_07511_));
 sg13g2_nand2b_1 _13306_ (.Y(_07512_),
    .B(_07511_),
    .A_N(net1036));
 sg13g2_nand2b_1 _13307_ (.Y(_07513_),
    .B(net1036),
    .A_N(_07511_));
 sg13g2_and3_1 _13308_ (.X(_07514_),
    .A(_07509_),
    .B(_07512_),
    .C(_07513_));
 sg13g2_buf_2 _13309_ (.A(_07514_),
    .X(_07515_));
 sg13g2_buf_2 _13310_ (.A(\top_ihp.oisc.op_b[17] ),
    .X(_07516_));
 sg13g2_buf_1 _13311_ (.A(\top_ihp.oisc.op_a[17] ),
    .X(_07517_));
 sg13g2_nor2b_1 _13312_ (.A(_07516_),
    .B_N(net1035),
    .Y(_07518_));
 sg13g2_nor2b_1 _13313_ (.A(net1035),
    .B_N(_07516_),
    .Y(_07519_));
 sg13g2_buf_2 _13314_ (.A(_07519_),
    .X(_07520_));
 sg13g2_buf_2 _13315_ (.A(\top_ihp.oisc.op_a[14] ),
    .X(_07521_));
 sg13g2_buf_1 _13316_ (.A(\top_ihp.oisc.op_b[14] ),
    .X(_07522_));
 sg13g2_xor2_1 _13317_ (.B(_07522_),
    .A(_07521_),
    .X(_07523_));
 sg13g2_nor3_1 _13318_ (.A(_07518_),
    .B(_07520_),
    .C(_07523_),
    .Y(_07524_));
 sg13g2_buf_1 _13319_ (.A(\top_ihp.oisc.op_a[13] ),
    .X(_07525_));
 sg13g2_buf_2 _13320_ (.A(\top_ihp.oisc.op_b[13] ),
    .X(_07526_));
 sg13g2_xor2_1 _13321_ (.B(_07526_),
    .A(net1034),
    .X(_07527_));
 sg13g2_buf_2 _13322_ (.A(\top_ihp.oisc.op_a[12] ),
    .X(_07528_));
 sg13g2_buf_2 _13323_ (.A(\top_ihp.oisc.op_b[12] ),
    .X(_07529_));
 sg13g2_xor2_1 _13324_ (.B(_07529_),
    .A(_07528_),
    .X(_07530_));
 sg13g2_buf_2 _13325_ (.A(\top_ihp.oisc.op_a[11] ),
    .X(_07531_));
 sg13g2_buf_2 _13326_ (.A(\top_ihp.oisc.op_b[11] ),
    .X(_07532_));
 sg13g2_xor2_1 _13327_ (.B(_07532_),
    .A(_07531_),
    .X(_07533_));
 sg13g2_buf_2 _13328_ (.A(\top_ihp.oisc.op_a[10] ),
    .X(_07534_));
 sg13g2_buf_2 _13329_ (.A(\top_ihp.oisc.op_b[10] ),
    .X(_07535_));
 sg13g2_xor2_1 _13330_ (.B(_07535_),
    .A(_07534_),
    .X(_07536_));
 sg13g2_nor4_1 _13331_ (.A(_07527_),
    .B(_07530_),
    .C(_07533_),
    .D(_07536_),
    .Y(_07537_));
 sg13g2_nand3_1 _13332_ (.B(_07524_),
    .C(_07537_),
    .A(_07515_),
    .Y(_07538_));
 sg13g2_buf_8 _13333_ (.A(\top_ihp.oisc.op_a[7] ),
    .X(_07539_));
 sg13g2_buf_2 _13334_ (.A(\top_ihp.oisc.op_b[7] ),
    .X(_07540_));
 sg13g2_nor2b_1 _13335_ (.A(net1033),
    .B_N(_07540_),
    .Y(_07541_));
 sg13g2_nor2b_1 _13336_ (.A(_07540_),
    .B_N(\top_ihp.oisc.op_a[7] ),
    .Y(_07542_));
 sg13g2_buf_1 _13337_ (.A(\top_ihp.oisc.op_a[8] ),
    .X(_07543_));
 sg13g2_buf_2 _13338_ (.A(\top_ihp.oisc.op_b[8] ),
    .X(_07544_));
 sg13g2_xor2_1 _13339_ (.B(_07544_),
    .A(_07543_),
    .X(_07545_));
 sg13g2_or3_1 _13340_ (.A(_07541_),
    .B(_07542_),
    .C(_07545_),
    .X(_07546_));
 sg13g2_buf_2 _13341_ (.A(\top_ihp.oisc.op_a[9] ),
    .X(_07547_));
 sg13g2_buf_1 _13342_ (.A(\top_ihp.oisc.op_b[9] ),
    .X(_07548_));
 sg13g2_xor2_1 _13343_ (.B(_07548_),
    .A(net1032),
    .X(_07549_));
 sg13g2_buf_1 _13344_ (.A(\top_ihp.oisc.op_a[6] ),
    .X(_07550_));
 sg13g2_buf_2 _13345_ (.A(\top_ihp.oisc.op_b[6] ),
    .X(_07551_));
 sg13g2_inv_1 _13346_ (.Y(_07552_),
    .A(_07551_));
 sg13g2_nor2_1 _13347_ (.A(net1031),
    .B(_07552_),
    .Y(_07553_));
 sg13g2_nor2b_1 _13348_ (.A(_07551_),
    .B_N(\top_ihp.oisc.op_a[6] ),
    .Y(_07554_));
 sg13g2_or4_1 _13349_ (.A(_07546_),
    .B(_07549_),
    .C(_07553_),
    .D(_07554_),
    .X(_07555_));
 sg13g2_nor2_1 _13350_ (.A(_07538_),
    .B(_07555_),
    .Y(_07556_));
 sg13g2_nor2b_1 _13351_ (.A(_07506_),
    .B_N(_07556_),
    .Y(_07557_));
 sg13g2_inv_1 _13352_ (.Y(_07558_),
    .A(_07516_));
 sg13g2_inv_1 _13353_ (.Y(_07559_),
    .A(_07511_));
 sg13g2_nand2b_1 _13354_ (.Y(_07560_),
    .B(_07522_),
    .A_N(_07521_));
 sg13g2_nor2_1 _13355_ (.A(_07559_),
    .B(_07560_),
    .Y(_07561_));
 sg13g2_a21oi_1 _13356_ (.A1(_07559_),
    .A2(_07560_),
    .Y(_07562_),
    .B1(_07510_));
 sg13g2_o21ai_1 _13357_ (.B1(_07508_),
    .Y(_07563_),
    .A1(_07561_),
    .A2(_07562_));
 sg13g2_nor3_1 _13358_ (.A(_07508_),
    .B(_07561_),
    .C(_07562_),
    .Y(_07564_));
 sg13g2_a221oi_1 _13359_ (.B2(_07563_),
    .C1(_07564_),
    .B1(_07507_),
    .A1(net1035),
    .Y(_07565_),
    .A2(_07558_));
 sg13g2_or2_1 _13360_ (.X(_07566_),
    .B(_07565_),
    .A(_07520_));
 sg13g2_nor2b_1 _13361_ (.A(_07534_),
    .B_N(_07535_),
    .Y(_07567_));
 sg13g2_buf_1 _13362_ (.A(_07567_),
    .X(_07568_));
 sg13g2_nor2_1 _13363_ (.A(_07532_),
    .B(_07568_),
    .Y(_07569_));
 sg13g2_inv_1 _13364_ (.Y(_07570_),
    .A(_07531_));
 sg13g2_a21oi_1 _13365_ (.A1(_07532_),
    .A2(_07568_),
    .Y(_07571_),
    .B1(_07570_));
 sg13g2_inv_1 _13366_ (.Y(_07572_),
    .A(_07528_));
 sg13g2_nor2b_1 _13367_ (.A(net1034),
    .B_N(_07526_),
    .Y(_07573_));
 sg13g2_a21oi_1 _13368_ (.A1(_07572_),
    .A2(_07529_),
    .Y(_07574_),
    .B1(_07573_));
 sg13g2_o21ai_1 _13369_ (.B1(_07574_),
    .Y(_07575_),
    .A1(_07569_),
    .A2(_07571_));
 sg13g2_inv_1 _13370_ (.Y(_07576_),
    .A(_07526_));
 sg13g2_nor3_1 _13371_ (.A(_07572_),
    .B(_07529_),
    .C(_07573_),
    .Y(_07577_));
 sg13g2_a21oi_1 _13372_ (.A1(net1034),
    .A2(_07576_),
    .Y(_07578_),
    .B1(_07577_));
 sg13g2_and4_1 _13373_ (.A(_07515_),
    .B(_07524_),
    .C(_07575_),
    .D(_07578_),
    .X(_07579_));
 sg13g2_buf_2 _13374_ (.A(_07543_),
    .X(_07580_));
 sg13g2_inv_1 _13375_ (.Y(_07581_),
    .A(_07544_));
 sg13g2_nand2_1 _13376_ (.Y(_07582_),
    .A(net1015),
    .B(_07581_));
 sg13g2_inv_1 _13377_ (.Y(_07583_),
    .A(_07540_));
 sg13g2_nand2b_1 _13378_ (.Y(_07584_),
    .B(_07544_),
    .A_N(net1015));
 sg13g2_nand2b_1 _13379_ (.Y(_07585_),
    .B(_07551_),
    .A_N(_07550_));
 sg13g2_nand3_1 _13380_ (.B(_07584_),
    .C(_07585_),
    .A(_07583_),
    .Y(_07586_));
 sg13g2_nand3b_1 _13381_ (.B(_07551_),
    .C(_07540_),
    .Y(_07587_),
    .A_N(_07550_));
 sg13g2_nand3_1 _13382_ (.B(_07584_),
    .C(_07587_),
    .A(net1033),
    .Y(_07588_));
 sg13g2_nand4_1 _13383_ (.B(_07582_),
    .C(_07586_),
    .A(_07548_),
    .Y(_07589_),
    .D(_07588_));
 sg13g2_nand2_1 _13384_ (.Y(_07590_),
    .A(net1033),
    .B(_07587_));
 sg13g2_a221oi_1 _13385_ (.B2(_07585_),
    .C1(net1032),
    .B1(_07583_),
    .A1(net1015),
    .Y(_07591_),
    .A2(_07581_));
 sg13g2_inv_1 _13386_ (.Y(_07592_),
    .A(_07548_));
 sg13g2_a21oi_1 _13387_ (.A1(_07592_),
    .A2(_07584_),
    .Y(_07593_),
    .B1(net1032));
 sg13g2_a21oi_1 _13388_ (.A1(_07590_),
    .A2(_07591_),
    .Y(_07594_),
    .B1(_07593_));
 sg13g2_a21oi_1 _13389_ (.A1(_07589_),
    .A2(_07594_),
    .Y(_07595_),
    .B1(_07538_));
 sg13g2_or2_1 _13390_ (.X(_07596_),
    .B(_07595_),
    .A(_07579_));
 sg13g2_or4_1 _13391_ (.A(_07471_),
    .B(_07557_),
    .C(_07566_),
    .D(_07596_),
    .X(_07597_));
 sg13g2_buf_1 _13392_ (.A(_07597_),
    .X(_07598_));
 sg13g2_xnor2_1 _13393_ (.Y(_07599_),
    .A(_07444_),
    .B(net1044));
 sg13g2_xnor2_1 _13394_ (.Y(_07600_),
    .A(_07442_),
    .B(_07443_));
 sg13g2_a21oi_1 _13395_ (.A1(_07599_),
    .A2(_07600_),
    .Y(_07601_),
    .B1(_07449_));
 sg13g2_nor2_1 _13396_ (.A(_07465_),
    .B(_07468_),
    .Y(_07602_));
 sg13g2_nor2b_1 _13397_ (.A(_07462_),
    .B_N(_07461_),
    .Y(_07603_));
 sg13g2_xor2_1 _13398_ (.B(_07453_),
    .A(net1042),
    .X(_07604_));
 sg13g2_xnor2_1 _13399_ (.Y(_07605_),
    .A(_07450_),
    .B(_07452_));
 sg13g2_nand2b_1 _13400_ (.Y(_07606_),
    .B(_07605_),
    .A_N(_07604_));
 sg13g2_buf_1 _13401_ (.A(_07606_),
    .X(_07607_));
 sg13g2_xor2_1 _13402_ (.B(_07456_),
    .A(net1043),
    .X(_07608_));
 sg13g2_nor4_1 _13403_ (.A(_07464_),
    .B(_07603_),
    .C(_07607_),
    .D(_07608_),
    .Y(_07609_));
 sg13g2_nor3_1 _13404_ (.A(_07449_),
    .B(_07602_),
    .C(_07609_),
    .Y(_07610_));
 sg13g2_nor2_2 _13405_ (.A(_07601_),
    .B(_07610_),
    .Y(_07611_));
 sg13g2_buf_2 _13406_ (.A(\top_ihp.oisc.op_b[24] ),
    .X(_07612_));
 sg13g2_inv_1 _13407_ (.Y(_07613_),
    .A(_07612_));
 sg13g2_buf_1 _13408_ (.A(\top_ihp.oisc.op_a[26] ),
    .X(_07614_));
 sg13g2_buf_2 _13409_ (.A(\top_ihp.oisc.op_b[26] ),
    .X(_07615_));
 sg13g2_nor2b_1 _13410_ (.A(net1030),
    .B_N(_07615_),
    .Y(_07616_));
 sg13g2_inv_2 _13411_ (.Y(_07617_),
    .A(net1030));
 sg13g2_nor2_1 _13412_ (.A(_07615_),
    .B(_07617_),
    .Y(_07618_));
 sg13g2_or2_1 _13413_ (.X(_07619_),
    .B(_07618_),
    .A(_07616_));
 sg13g2_buf_1 _13414_ (.A(_07619_),
    .X(_07620_));
 sg13g2_buf_1 _13415_ (.A(\top_ihp.oisc.op_a[25] ),
    .X(_07621_));
 sg13g2_buf_1 _13416_ (.A(\top_ihp.oisc.op_b[25] ),
    .X(_07622_));
 sg13g2_nand2b_1 _13417_ (.Y(_07623_),
    .B(_07622_),
    .A_N(_07621_));
 sg13g2_buf_2 _13418_ (.A(_07623_),
    .X(_07624_));
 sg13g2_nand3_1 _13419_ (.B(net904),
    .C(_07624_),
    .A(_07613_),
    .Y(_07625_));
 sg13g2_buf_2 _13420_ (.A(\top_ihp.oisc.op_a[24] ),
    .X(_07626_));
 sg13g2_nand3_1 _13421_ (.B(net904),
    .C(_07624_),
    .A(net1029),
    .Y(_07627_));
 sg13g2_a22oi_1 _13422_ (.Y(_07628_),
    .B1(_07625_),
    .B2(_07627_),
    .A2(_07611_),
    .A1(_07598_));
 sg13g2_nor4_1 _13423_ (.A(_07471_),
    .B(_07557_),
    .C(_07566_),
    .D(_07596_),
    .Y(_07629_));
 sg13g2_buf_2 _13424_ (.A(_07629_),
    .X(_07630_));
 sg13g2_or2_1 _13425_ (.X(_07631_),
    .B(_07610_),
    .A(_07601_));
 sg13g2_buf_1 _13426_ (.A(_07631_),
    .X(_07632_));
 sg13g2_nor2b_1 _13427_ (.A(_07622_),
    .B_N(_07621_),
    .Y(_07633_));
 sg13g2_buf_1 _13428_ (.A(_07633_),
    .X(_07634_));
 sg13g2_nand2b_1 _13429_ (.Y(_07635_),
    .B(_07612_),
    .A_N(net985));
 sg13g2_nor4_2 _13430_ (.A(net904),
    .B(_07630_),
    .C(_07632_),
    .Y(_07636_),
    .D(_07635_));
 sg13g2_or2_1 _13431_ (.X(_07637_),
    .B(net985),
    .A(net1029));
 sg13g2_nor4_1 _13432_ (.A(net904),
    .B(_07630_),
    .C(_07632_),
    .D(_07637_),
    .Y(_07638_));
 sg13g2_nand2_1 _13433_ (.Y(_07639_),
    .A(_07620_),
    .B(_07634_));
 sg13g2_nand4_1 _13434_ (.B(_07613_),
    .C(net904),
    .A(net1029),
    .Y(_07640_),
    .D(_07624_));
 sg13g2_nor2_1 _13435_ (.A(net904),
    .B(_07624_),
    .Y(_07641_));
 sg13g2_nand2b_1 _13436_ (.Y(_07642_),
    .B(_07612_),
    .A_N(net1029));
 sg13g2_nor3_1 _13437_ (.A(net904),
    .B(_07642_),
    .C(net985),
    .Y(_07643_));
 sg13g2_nor2_1 _13438_ (.A(_07641_),
    .B(_07643_),
    .Y(_07644_));
 sg13g2_nand3_1 _13439_ (.B(_07640_),
    .C(_07644_),
    .A(_07639_),
    .Y(_07645_));
 sg13g2_nor4_2 _13440_ (.A(_07628_),
    .B(_07636_),
    .C(_07638_),
    .Y(_07646_),
    .D(_07645_));
 sg13g2_inv_1 _13441_ (.Y(_07647_),
    .A(_07417_));
 sg13g2_buf_1 _13442_ (.A(_07647_),
    .X(_07648_));
 sg13g2_nor2_1 _13443_ (.A(_07648_),
    .B(_07617_),
    .Y(_07649_));
 sg13g2_a21oi_1 _13444_ (.A1(net777),
    .A2(_07646_),
    .Y(_07650_),
    .B1(_07649_));
 sg13g2_buf_1 _13445_ (.A(\top_ihp.wb_spi.state ),
    .X(_07651_));
 sg13g2_inv_2 _13446_ (.Y(_07652_),
    .A(_07651_));
 sg13g2_inv_1 _13447_ (.Y(_07653_),
    .A(_07419_));
 sg13g2_nand2_1 _13448_ (.Y(_07654_),
    .A(_07422_),
    .B(_07435_));
 sg13g2_nor2_1 _13449_ (.A(_07653_),
    .B(_07654_),
    .Y(_07655_));
 sg13g2_buf_2 _13450_ (.A(_07655_),
    .X(_07656_));
 sg13g2_buf_1 _13451_ (.A(_07656_),
    .X(_07657_));
 sg13g2_buf_1 _13452_ (.A(net824),
    .X(_07658_));
 sg13g2_nand2_1 _13453_ (.Y(_07659_),
    .A(_07652_),
    .B(net806));
 sg13g2_buf_1 _13454_ (.A(\top_ihp.wb_spi.bits_left[0] ),
    .X(_07660_));
 sg13g2_inv_1 _13455_ (.Y(_07661_),
    .A(\top_ihp.wb_spi.bits_left[1] ));
 sg13g2_buf_1 _13456_ (.A(\top_ihp.wb_spi.bits_left[2] ),
    .X(_07662_));
 sg13g2_nand2b_1 _13457_ (.Y(_07663_),
    .B(\top_ihp.spi_clk_o ),
    .A_N(\top_ihp.wb_spi.spi_clk_cnt[0] ));
 sg13g2_buf_1 _13458_ (.A(_07663_),
    .X(_07664_));
 sg13g2_nor2_1 _13459_ (.A(_07662_),
    .B(_07664_),
    .Y(_07665_));
 sg13g2_buf_1 _13460_ (.A(\top_ihp.wb_spi.bits_left[4] ),
    .X(_07666_));
 sg13g2_nor2_1 _13461_ (.A(_07666_),
    .B(\top_ihp.wb_spi.bits_left[5] ),
    .Y(_07667_));
 sg13g2_nand4_1 _13462_ (.B(_07661_),
    .C(_07665_),
    .A(_07660_),
    .Y(_07668_),
    .D(_07667_));
 sg13g2_o21ai_1 _13463_ (.B1(_07651_),
    .Y(_07669_),
    .A1(\top_ihp.wb_spi.bits_left[3] ),
    .A2(_07668_));
 sg13g2_o21ai_1 _13464_ (.B1(_07669_),
    .Y(_13210_),
    .A1(_07650_),
    .A2(_07659_));
 sg13g2_inv_1 _13465_ (.Y(_07670_),
    .A(_07669_));
 sg13g2_a21o_1 _13466_ (.A2(_07646_),
    .A1(net777),
    .B1(_07649_),
    .X(_07671_));
 sg13g2_nand2_1 _13467_ (.Y(_07672_),
    .A(_07419_),
    .B(_07437_));
 sg13g2_buf_2 _13468_ (.A(_07672_),
    .X(_07673_));
 sg13g2_buf_1 _13469_ (.A(_07651_),
    .X(_07674_));
 sg13g2_buf_1 _13470_ (.A(net1014),
    .X(_07675_));
 sg13g2_a21oi_1 _13471_ (.A1(_07671_),
    .A2(_07673_),
    .Y(_07676_),
    .B1(_07675_));
 sg13g2_nor2_1 _13472_ (.A(_07670_),
    .B(_07676_),
    .Y(_13209_));
 sg13g2_inv_1 _13473_ (.Y(_07677_),
    .A(_00072_));
 sg13g2_buf_1 _13474_ (.A(_07418_),
    .X(_07678_));
 sg13g2_buf_1 _13475_ (.A(\top_ihp.oisc.op_a[28] ),
    .X(_07679_));
 sg13g2_buf_1 _13476_ (.A(\top_ihp.oisc.op_b[28] ),
    .X(_07680_));
 sg13g2_buf_2 _13477_ (.A(\top_ihp.oisc.op_a[27] ),
    .X(_07681_));
 sg13g2_buf_1 _13478_ (.A(\top_ihp.oisc.op_b[27] ),
    .X(_07682_));
 sg13g2_nand2b_1 _13479_ (.Y(_07683_),
    .B(_07682_),
    .A_N(_07681_));
 sg13g2_buf_1 _13480_ (.A(_07683_),
    .X(_07684_));
 sg13g2_o21ai_1 _13481_ (.B1(_07624_),
    .Y(_07685_),
    .A1(_07642_),
    .A2(net985));
 sg13g2_nand2_1 _13482_ (.Y(_07686_),
    .A(_07617_),
    .B(_07685_));
 sg13g2_o21ai_1 _13483_ (.B1(_07615_),
    .Y(_07687_),
    .A1(_07617_),
    .A2(_07685_));
 sg13g2_and2_1 _13484_ (.A(_07686_),
    .B(_07687_),
    .X(_07688_));
 sg13g2_nor2b_1 _13485_ (.A(_07682_),
    .B_N(_07681_),
    .Y(_07689_));
 sg13g2_buf_1 _13486_ (.A(_07689_),
    .X(_07690_));
 sg13g2_a21o_1 _13487_ (.A2(_07688_),
    .A1(_07684_),
    .B1(_07690_),
    .X(_07691_));
 sg13g2_buf_1 _13488_ (.A(_07691_),
    .X(_07692_));
 sg13g2_xnor2_1 _13489_ (.Y(_07693_),
    .A(net1029),
    .B(_07612_));
 sg13g2_nor2b_1 _13490_ (.A(_07621_),
    .B_N(_07622_),
    .Y(_07694_));
 sg13g2_nor2b_1 _13491_ (.A(_07681_),
    .B_N(_07682_),
    .Y(_07695_));
 sg13g2_or2_1 _13492_ (.X(_07696_),
    .B(_07690_),
    .A(_07695_));
 sg13g2_buf_1 _13493_ (.A(_07696_),
    .X(_07697_));
 sg13g2_nor4_2 _13494_ (.A(net904),
    .B(_07694_),
    .C(net985),
    .Y(_07698_),
    .D(_07697_));
 sg13g2_nand2_2 _13495_ (.Y(_07699_),
    .A(_07693_),
    .B(_07698_));
 sg13g2_nand3_1 _13496_ (.B(_07692_),
    .C(_07699_),
    .A(net1027),
    .Y(_07700_));
 sg13g2_o21ai_1 _13497_ (.B1(_07700_),
    .Y(_07701_),
    .A1(net1027),
    .A2(_07692_));
 sg13g2_nand2_1 _13498_ (.Y(_07702_),
    .A(net1027),
    .B(_07692_));
 sg13g2_a21oi_1 _13499_ (.A1(_07598_),
    .A2(_07611_),
    .Y(_07703_),
    .B1(_07702_));
 sg13g2_nor4_2 _13500_ (.A(net1027),
    .B(_07630_),
    .C(_07632_),
    .Y(_07704_),
    .D(_07699_));
 sg13g2_or3_1 _13501_ (.A(_07701_),
    .B(_07703_),
    .C(_07704_),
    .X(_07705_));
 sg13g2_inv_1 _13502_ (.Y(_07706_),
    .A(net1028));
 sg13g2_nand2b_1 _13503_ (.Y(_07707_),
    .B(net984),
    .A_N(_07438_));
 sg13g2_buf_2 _13504_ (.A(_07707_),
    .X(_07708_));
 sg13g2_nor2_1 _13505_ (.A(_07706_),
    .B(_07708_),
    .Y(_07709_));
 sg13g2_nand2_1 _13506_ (.Y(_07710_),
    .A(_07706_),
    .B(net807));
 sg13g2_nor4_1 _13507_ (.A(_07701_),
    .B(_07703_),
    .C(_07704_),
    .D(_07710_),
    .Y(_07711_));
 sg13g2_a221oi_1 _13508_ (.B2(_07709_),
    .C1(_07711_),
    .B1(_07705_),
    .A1(_07678_),
    .Y(_07712_),
    .A2(net1028));
 sg13g2_nor2_1 _13509_ (.A(_07677_),
    .B(_07712_),
    .Y(_00003_));
 sg13g2_buf_2 _13510_ (.A(\top_ihp.wb_imem.state[0] ),
    .X(_07713_));
 sg13g2_inv_1 _13511_ (.Y(_07714_),
    .A(_07713_));
 sg13g2_buf_1 _13512_ (.A(\top_ihp.oisc.op_a[30] ),
    .X(_07715_));
 sg13g2_and2_1 _13513_ (.A(net1017),
    .B(net1026),
    .X(_07716_));
 sg13g2_nand3b_1 _13514_ (.B(_07598_),
    .C(_07611_),
    .Y(_07717_),
    .A_N(_07699_));
 sg13g2_a21oi_1 _13515_ (.A1(_07684_),
    .A2(_07688_),
    .Y(_07718_),
    .B1(_07690_));
 sg13g2_buf_1 _13516_ (.A(\top_ihp.oisc.op_b[30] ),
    .X(_07719_));
 sg13g2_xor2_1 _13517_ (.B(net1026),
    .A(_07719_),
    .X(_07720_));
 sg13g2_buf_2 _13518_ (.A(\top_ihp.oisc.op_a[29] ),
    .X(_07721_));
 sg13g2_buf_2 _13519_ (.A(\top_ihp.oisc.op_b[29] ),
    .X(_07722_));
 sg13g2_nor2b_1 _13520_ (.A(net1028),
    .B_N(net1027),
    .Y(_07723_));
 sg13g2_nor2_1 _13521_ (.A(_07722_),
    .B(_07723_),
    .Y(_07724_));
 sg13g2_nand2_1 _13522_ (.Y(_07725_),
    .A(_07722_),
    .B(_07723_));
 sg13g2_o21ai_1 _13523_ (.B1(_07725_),
    .Y(_07726_),
    .A1(_07721_),
    .A2(_07724_));
 sg13g2_xnor2_1 _13524_ (.Y(_07727_),
    .A(_07720_),
    .B(_07726_));
 sg13g2_nor2_1 _13525_ (.A(_07718_),
    .B(_07727_),
    .Y(_07728_));
 sg13g2_nand2b_1 _13526_ (.Y(_07729_),
    .B(net1028),
    .A_N(net1027));
 sg13g2_buf_1 _13527_ (.A(_07729_),
    .X(_07730_));
 sg13g2_nand2_1 _13528_ (.Y(_07731_),
    .A(_07722_),
    .B(_07730_));
 sg13g2_nor2_1 _13529_ (.A(_07722_),
    .B(_07730_),
    .Y(_07732_));
 sg13g2_a21oi_1 _13530_ (.A1(_07721_),
    .A2(_07731_),
    .Y(_07733_),
    .B1(_07732_));
 sg13g2_xor2_1 _13531_ (.B(_07733_),
    .A(_07720_),
    .X(_07734_));
 sg13g2_inv_1 _13532_ (.Y(_07735_),
    .A(_07734_));
 sg13g2_nor4_1 _13533_ (.A(_07630_),
    .B(_07632_),
    .C(_07699_),
    .D(_07735_),
    .Y(_07736_));
 sg13g2_a221oi_1 _13534_ (.B2(_07718_),
    .C1(_07736_),
    .B1(_07734_),
    .A1(_07717_),
    .Y(_07737_),
    .A2(_07728_));
 sg13g2_buf_2 _13535_ (.A(_07737_),
    .X(_07738_));
 sg13g2_nor2_1 _13536_ (.A(_07708_),
    .B(_07656_),
    .Y(_07739_));
 sg13g2_a22oi_1 _13537_ (.Y(_07740_),
    .B1(_07738_),
    .B2(_07739_),
    .A2(_07716_),
    .A1(_07673_));
 sg13g2_buf_2 _13538_ (.A(_07740_),
    .X(_07741_));
 sg13g2_buf_8 _13539_ (.A(\top_ihp.wb_imem.bits_left[2] ),
    .X(_07742_));
 sg13g2_buf_2 _13540_ (.A(\top_ihp.wb_imem.bits_left[4] ),
    .X(_07743_));
 sg13g2_nor4_2 _13541_ (.A(_07742_),
    .B(\top_ihp.wb_imem.bits_left[3] ),
    .C(\top_ihp.wb_imem.bits_left[5] ),
    .Y(_07744_),
    .D(_07743_));
 sg13g2_buf_1 _13542_ (.A(\top_ihp.wb_imem.bits_left[1] ),
    .X(_07745_));
 sg13g2_buf_2 _13543_ (.A(\top_ihp.wb_imem.bits_left[0] ),
    .X(_07746_));
 sg13g2_nor2b_1 _13544_ (.A(_07745_),
    .B_N(_07746_),
    .Y(_07747_));
 sg13g2_and2_1 _13545_ (.A(_07744_),
    .B(_07747_),
    .X(_07748_));
 sg13g2_buf_1 _13546_ (.A(_07748_),
    .X(_07749_));
 sg13g2_buf_2 _13547_ (.A(\top_ihp.wb_imem.state[2] ),
    .X(_07750_));
 sg13g2_nand2b_1 _13548_ (.Y(_07751_),
    .B(_07750_),
    .A_N(_07749_));
 sg13g2_o21ai_1 _13549_ (.B1(_07751_),
    .Y(_00001_),
    .A1(_07714_),
    .A2(_07741_));
 sg13g2_buf_1 _13550_ (.A(_00077_),
    .X(_07752_));
 sg13g2_nor2_1 _13551_ (.A(_07746_),
    .B(_07745_),
    .Y(_07753_));
 sg13g2_buf_2 _13552_ (.A(_07753_),
    .X(_07754_));
 sg13g2_and2_1 _13553_ (.A(_07744_),
    .B(_07754_),
    .X(_07755_));
 sg13g2_buf_8 _13554_ (.A(_07755_),
    .X(_07756_));
 sg13g2_buf_8 _13555_ (.A(net878),
    .X(_07757_));
 sg13g2_buf_8 _13556_ (.A(_07757_),
    .X(_07758_));
 sg13g2_nand2_1 _13557_ (.Y(_07759_),
    .A(_07750_),
    .B(_07749_));
 sg13g2_o21ai_1 _13558_ (.B1(_07759_),
    .Y(_00000_),
    .A1(_07752_),
    .A2(net846));
 sg13g2_buf_1 _13559_ (.A(\top_ihp.wb_uart.uart_rx.state[0] ),
    .X(_07760_));
 sg13g2_inv_2 _13560_ (.Y(_07761_),
    .A(_07760_));
 sg13g2_buf_1 _13561_ (.A(\top_ihp.wb_uart.uart_rx.state[1] ),
    .X(_07762_));
 sg13g2_inv_1 _13562_ (.Y(_07763_),
    .A(net1025));
 sg13g2_buf_1 _13563_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ),
    .X(_07764_));
 sg13g2_buf_1 _13564_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ),
    .X(_07765_));
 sg13g2_buf_1 _13565_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[13] ),
    .X(_07766_));
 sg13g2_nor4_1 _13566_ (.A(_07764_),
    .B(_07765_),
    .C(_07766_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ),
    .Y(_07767_));
 sg13g2_buf_1 _13567_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ),
    .X(_07768_));
 sg13g2_buf_1 _13568_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[18] ),
    .X(_07769_));
 sg13g2_buf_1 _13569_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ),
    .X(_07770_));
 sg13g2_nor4_1 _13570_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .B(_07768_),
    .C(_07769_),
    .D(_07770_),
    .Y(_07771_));
 sg13g2_buf_1 _13571_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[23] ),
    .X(_07772_));
 sg13g2_buf_1 _13572_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ),
    .X(_07773_));
 sg13g2_nor4_1 _13573_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ),
    .B(_07772_),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .D(_07773_),
    .Y(_07774_));
 sg13g2_buf_1 _13574_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ),
    .X(_07775_));
 sg13g2_nor3_1 _13575_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .B(_07775_),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ),
    .Y(_07776_));
 sg13g2_nand4_1 _13576_ (.B(_07771_),
    .C(_07774_),
    .A(_07767_),
    .Y(_07777_),
    .D(_07776_));
 sg13g2_buf_1 _13577_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[29] ),
    .X(_07778_));
 sg13g2_nor4_1 _13578_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .D(_07778_),
    .Y(_07779_));
 sg13g2_buf_1 _13579_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[11] ),
    .X(_07780_));
 sg13g2_buf_1 _13580_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ),
    .X(_07781_));
 sg13g2_buf_1 _13581_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .X(_07782_));
 sg13g2_nor4_1 _13582_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .B(_07780_),
    .C(_07781_),
    .D(_07782_),
    .Y(_07783_));
 sg13g2_nand2_1 _13583_ (.Y(_07784_),
    .A(_07779_),
    .B(_07783_));
 sg13g2_buf_8 _13584_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[0] ),
    .X(_07785_));
 sg13g2_inv_1 _13585_ (.Y(_07786_),
    .A(_07785_));
 sg13g2_buf_1 _13586_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ),
    .X(_07787_));
 sg13g2_inv_1 _13587_ (.Y(_07788_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ));
 sg13g2_buf_1 _13588_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[4] ),
    .X(_07789_));
 sg13g2_inv_1 _13589_ (.Y(_07790_),
    .A(_07789_));
 sg13g2_buf_1 _13590_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ),
    .X(_07791_));
 sg13g2_nor4_1 _13591_ (.A(_07788_),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ),
    .C(_07790_),
    .D(_07791_),
    .Y(_07792_));
 sg13g2_nand3_1 _13592_ (.B(_07787_),
    .C(_07792_),
    .A(_07786_),
    .Y(_07793_));
 sg13g2_buf_8 _13593_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[2] ),
    .X(_07794_));
 sg13g2_buf_8 _13594_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[3] ),
    .X(_07795_));
 sg13g2_buf_8 _13595_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[1] ),
    .X(_07796_));
 sg13g2_nand3b_1 _13596_ (.B(_07795_),
    .C(_07796_),
    .Y(_07797_),
    .A_N(_07794_));
 sg13g2_nor4_1 _13597_ (.A(_07777_),
    .B(_07784_),
    .C(_07793_),
    .D(_07797_),
    .Y(_07798_));
 sg13g2_buf_1 _13598_ (.A(_07798_),
    .X(_07799_));
 sg13g2_nand2_1 _13599_ (.Y(_07800_),
    .A(net1044),
    .B(_07464_));
 sg13g2_inv_1 _13600_ (.Y(_07801_),
    .A(_07444_));
 sg13g2_o21ai_1 _13601_ (.B1(_07801_),
    .Y(_07802_),
    .A1(net1044),
    .A2(_07464_));
 sg13g2_nand2_1 _13602_ (.Y(_07803_),
    .A(_07600_),
    .B(_07693_));
 sg13g2_a21oi_1 _13603_ (.A1(_07800_),
    .A2(_07802_),
    .Y(_07804_),
    .B1(_07803_));
 sg13g2_nor2b_1 _13604_ (.A(_07442_),
    .B_N(_07443_),
    .Y(_07805_));
 sg13g2_nand2_1 _13605_ (.Y(_07806_),
    .A(_07612_),
    .B(_07805_));
 sg13g2_nor2_1 _13606_ (.A(_07612_),
    .B(_07805_),
    .Y(_07807_));
 sg13g2_a21oi_1 _13607_ (.A1(net1029),
    .A2(_07806_),
    .Y(_07808_),
    .B1(_07807_));
 sg13g2_or2_1 _13608_ (.X(_07809_),
    .B(_07808_),
    .A(_07804_));
 sg13g2_buf_1 _13609_ (.A(_07809_),
    .X(_07810_));
 sg13g2_inv_1 _13610_ (.Y(_07811_),
    .A(_07621_));
 sg13g2_a21oi_1 _13611_ (.A1(_07622_),
    .A2(_07810_),
    .Y(_07812_),
    .B1(_07811_));
 sg13g2_nor2_1 _13612_ (.A(_07622_),
    .B(_07810_),
    .Y(_07813_));
 sg13g2_a21oi_1 _13613_ (.A1(_07706_),
    .A2(_07695_),
    .Y(_07814_),
    .B1(net1027));
 sg13g2_a21oi_1 _13614_ (.A1(net1028),
    .A2(_07684_),
    .Y(_07815_),
    .B1(_07814_));
 sg13g2_nor2_1 _13615_ (.A(_07616_),
    .B(_07815_),
    .Y(_07816_));
 sg13g2_o21ai_1 _13616_ (.B1(_07816_),
    .Y(_07817_),
    .A1(_07812_),
    .A2(_07813_));
 sg13g2_a21oi_1 _13617_ (.A1(_07618_),
    .A2(_07684_),
    .Y(_07818_),
    .B1(_07690_));
 sg13g2_o21ai_1 _13618_ (.B1(_07730_),
    .Y(_07819_),
    .A1(_07723_),
    .A2(_07818_));
 sg13g2_nor3_1 _13619_ (.A(_07722_),
    .B(_07708_),
    .C(_07819_),
    .Y(_07820_));
 sg13g2_a21o_1 _13620_ (.A2(_07820_),
    .A1(_07817_),
    .B1(net1017),
    .X(_07821_));
 sg13g2_buf_2 _13621_ (.A(\top_ihp.oisc.decoder.instruction[12] ),
    .X(_07822_));
 sg13g2_buf_1 _13622_ (.A(\top_ihp.oisc.decoder.instruction[13] ),
    .X(_07823_));
 sg13g2_buf_1 _13623_ (.A(_00070_),
    .X(_07824_));
 sg13g2_nand2_1 _13624_ (.Y(_07825_),
    .A(_07823_),
    .B(_07824_));
 sg13g2_o21ai_1 _13625_ (.B1(_07647_),
    .Y(_07826_),
    .A1(_07421_),
    .A2(_07654_));
 sg13g2_o21ai_1 _13626_ (.B1(_07826_),
    .Y(_07827_),
    .A1(_07822_),
    .A2(_07825_));
 sg13g2_buf_2 _13627_ (.A(_07827_),
    .X(_07828_));
 sg13g2_inv_1 _13628_ (.Y(_07829_),
    .A(_07824_));
 sg13g2_nor2_2 _13629_ (.A(_07823_),
    .B(_07829_),
    .Y(_07830_));
 sg13g2_or2_1 _13630_ (.X(_07831_),
    .B(_07830_),
    .A(_07828_));
 sg13g2_buf_1 _13631_ (.A(_07831_),
    .X(_07832_));
 sg13g2_and2_1 _13632_ (.A(_07721_),
    .B(_07832_),
    .X(_07833_));
 sg13g2_nor2b_1 _13633_ (.A(_07721_),
    .B_N(_07722_),
    .Y(_07834_));
 sg13g2_and3_1 _13634_ (.X(_07835_),
    .A(_07440_),
    .B(_07832_),
    .C(_07834_));
 sg13g2_nand2_1 _13635_ (.Y(_07836_),
    .A(_07706_),
    .B(net1027));
 sg13g2_nand2_1 _13636_ (.Y(_07837_),
    .A(_07730_),
    .B(_07818_));
 sg13g2_nand2_1 _13637_ (.Y(_07838_),
    .A(_07836_),
    .B(_07837_));
 sg13g2_and2_1 _13638_ (.A(_07838_),
    .B(_07817_),
    .X(_07839_));
 sg13g2_a22oi_1 _13639_ (.Y(_07840_),
    .B1(_07835_),
    .B2(_07839_),
    .A2(_07833_),
    .A1(_07821_));
 sg13g2_nand3b_1 _13640_ (.B(_07467_),
    .C(_07599_),
    .Y(_07841_),
    .A_N(_07464_));
 sg13g2_buf_1 _13641_ (.A(_07841_),
    .X(_07842_));
 sg13g2_nand2b_1 _13642_ (.Y(_07843_),
    .B(_07698_),
    .A_N(_07803_));
 sg13g2_nand2_1 _13643_ (.Y(_07844_),
    .A(_07836_),
    .B(_07730_));
 sg13g2_nor3_1 _13644_ (.A(_07842_),
    .B(_07843_),
    .C(_07844_),
    .Y(_07845_));
 sg13g2_nor2_1 _13645_ (.A(net1037),
    .B(_07473_),
    .Y(_07846_));
 sg13g2_inv_1 _13646_ (.Y(_07847_),
    .A(_07472_));
 sg13g2_nor2b_1 _13647_ (.A(_07474_),
    .B_N(_07475_),
    .Y(_07848_));
 sg13g2_a221oi_1 _13648_ (.B2(_07848_),
    .C1(\top_ihp.oisc.op_a[3] ),
    .B1(net1041),
    .A1(net1040),
    .Y(_07849_),
    .A2(_07847_));
 sg13g2_inv_1 _13649_ (.Y(_07850_),
    .A(_07477_));
 sg13g2_o21ai_1 _13650_ (.B1(_07850_),
    .Y(_07851_),
    .A1(_07478_),
    .A2(_07848_));
 sg13g2_a221oi_1 _13651_ (.B2(_07851_),
    .C1(_07485_),
    .B1(_07849_),
    .A1(_07493_),
    .Y(_07852_),
    .A2(_07846_));
 sg13g2_nand2_1 _13652_ (.Y(_07853_),
    .A(net1040),
    .B(_07847_));
 sg13g2_a21o_1 _13653_ (.A2(_07479_),
    .A1(_07476_),
    .B1(_07480_),
    .X(_07854_));
 sg13g2_nand2_1 _13654_ (.Y(_07855_),
    .A(net1037),
    .B(_07483_));
 sg13g2_a21oi_1 _13655_ (.A1(_07853_),
    .A2(_07854_),
    .Y(_07856_),
    .B1(_07855_));
 sg13g2_o21ai_1 _13656_ (.B1(net1031),
    .Y(_07857_),
    .A1(_07552_),
    .A2(_07498_));
 sg13g2_nand2_1 _13657_ (.Y(_07858_),
    .A(_07552_),
    .B(_07498_));
 sg13g2_a21oi_1 _13658_ (.A1(_07857_),
    .A2(_07858_),
    .Y(_07859_),
    .B1(_07501_));
 sg13g2_o21ai_1 _13659_ (.B1(_07859_),
    .Y(_07860_),
    .A1(_07852_),
    .A2(_07856_));
 sg13g2_nor2b_1 _13660_ (.A(_07486_),
    .B_N(net1039),
    .Y(_07861_));
 sg13g2_a21oi_1 _13661_ (.A1(_07502_),
    .A2(_07861_),
    .Y(_07862_),
    .B1(net1038));
 sg13g2_nor2_1 _13662_ (.A(_07502_),
    .B(_07861_),
    .Y(_07863_));
 sg13g2_nor4_1 _13663_ (.A(_07541_),
    .B(_07542_),
    .C(_07545_),
    .D(_07554_),
    .Y(_07864_));
 sg13g2_o21ai_1 _13664_ (.B1(_07864_),
    .Y(_07865_),
    .A1(_07862_),
    .A2(_07863_));
 sg13g2_nand2b_1 _13665_ (.Y(_07866_),
    .B(_07553_),
    .A_N(_07546_));
 sg13g2_or4_1 _13666_ (.A(_07530_),
    .B(_07533_),
    .C(_07536_),
    .D(_07549_),
    .X(_07867_));
 sg13g2_a21oi_1 _13667_ (.A1(_07865_),
    .A2(_07866_),
    .Y(_07868_),
    .B1(_07867_));
 sg13g2_or2_1 _13668_ (.X(_07869_),
    .B(_07568_),
    .A(_07548_));
 sg13g2_nand2b_1 _13669_ (.Y(_07870_),
    .B(net1032),
    .A_N(_07568_));
 sg13g2_nand2b_1 _13670_ (.Y(_07871_),
    .B(_07540_),
    .A_N(net1033));
 sg13g2_a21oi_1 _13671_ (.A1(_07581_),
    .A2(_07871_),
    .Y(_07872_),
    .B1(net1015));
 sg13g2_a221oi_1 _13672_ (.B2(_07870_),
    .C1(_07872_),
    .B1(_07869_),
    .A1(_07544_),
    .Y(_07873_),
    .A2(_07541_));
 sg13g2_nand2_1 _13673_ (.Y(_07874_),
    .A(net1032),
    .B(_07592_));
 sg13g2_nand2b_1 _13674_ (.Y(_07875_),
    .B(_07534_),
    .A_N(_07535_));
 sg13g2_o21ai_1 _13675_ (.B1(_07875_),
    .Y(_07876_),
    .A1(_07568_),
    .A2(_07874_));
 sg13g2_nor2_1 _13676_ (.A(_07873_),
    .B(_07876_),
    .Y(_07877_));
 sg13g2_nor2_1 _13677_ (.A(_07530_),
    .B(_07533_),
    .Y(_07878_));
 sg13g2_nor2b_1 _13678_ (.A(_07531_),
    .B_N(_07532_),
    .Y(_07879_));
 sg13g2_nor2_1 _13679_ (.A(_07529_),
    .B(_07879_),
    .Y(_07880_));
 sg13g2_a21oi_1 _13680_ (.A1(_07529_),
    .A2(_07879_),
    .Y(_07881_),
    .B1(_07572_));
 sg13g2_nor2_1 _13681_ (.A(_07880_),
    .B(_07881_),
    .Y(_07882_));
 sg13g2_a221oi_1 _13682_ (.B2(_07878_),
    .C1(_07882_),
    .B1(_07877_),
    .A1(_07860_),
    .Y(_07883_),
    .A2(_07868_));
 sg13g2_buf_2 _13683_ (.A(_07883_),
    .X(_07884_));
 sg13g2_nor2_1 _13684_ (.A(_07523_),
    .B(_07527_),
    .Y(_07885_));
 sg13g2_nor2_1 _13685_ (.A(_07518_),
    .B(_07520_),
    .Y(_07886_));
 sg13g2_nand2b_1 _13686_ (.Y(_07887_),
    .B(_07886_),
    .A_N(_07608_));
 sg13g2_nor2_1 _13687_ (.A(_07607_),
    .B(_07887_),
    .Y(_07888_));
 sg13g2_nand3_1 _13688_ (.B(_07885_),
    .C(_07888_),
    .A(_07515_),
    .Y(_07889_));
 sg13g2_inv_2 _13689_ (.Y(_07890_),
    .A(_07456_));
 sg13g2_nand2b_1 _13690_ (.Y(_07891_),
    .B(_07516_),
    .A_N(net1035));
 sg13g2_nor2_1 _13691_ (.A(_07890_),
    .B(_07891_),
    .Y(_07892_));
 sg13g2_a21oi_1 _13692_ (.A1(_07890_),
    .A2(_07891_),
    .Y(_07893_),
    .B1(net1043));
 sg13g2_nor3_1 _13693_ (.A(_07453_),
    .B(_07892_),
    .C(_07893_),
    .Y(_07894_));
 sg13g2_o21ai_1 _13694_ (.B1(_07453_),
    .Y(_07895_),
    .A1(_07892_),
    .A2(_07893_));
 sg13g2_o21ai_1 _13695_ (.B1(_07895_),
    .Y(_07896_),
    .A1(net1042),
    .A2(_07894_));
 sg13g2_inv_1 _13696_ (.Y(_07897_),
    .A(_07515_));
 sg13g2_inv_1 _13697_ (.Y(_07898_),
    .A(_07522_));
 sg13g2_nand2b_1 _13698_ (.Y(_07899_),
    .B(_07526_),
    .A_N(net1034));
 sg13g2_o21ai_1 _13699_ (.B1(_07521_),
    .Y(_07900_),
    .A1(_07898_),
    .A2(_07899_));
 sg13g2_o21ai_1 _13700_ (.B1(_07900_),
    .Y(_07901_),
    .A1(_07522_),
    .A2(_07573_));
 sg13g2_nand2b_1 _13701_ (.Y(_07902_),
    .B(_07512_),
    .A_N(_07508_));
 sg13g2_buf_1 _13702_ (.A(_07902_),
    .X(_07903_));
 sg13g2_nor2b_1 _13703_ (.A(net1036),
    .B_N(_07511_),
    .Y(_07904_));
 sg13g2_inv_1 _13704_ (.Y(_07905_),
    .A(_07507_));
 sg13g2_a21o_1 _13705_ (.A2(_07904_),
    .A1(_07508_),
    .B1(_07905_),
    .X(_07906_));
 sg13g2_buf_1 _13706_ (.A(_07906_),
    .X(_07907_));
 sg13g2_nand2_1 _13707_ (.Y(_07908_),
    .A(_07903_),
    .B(_07907_));
 sg13g2_o21ai_1 _13708_ (.B1(_07908_),
    .Y(_07909_),
    .A1(_07897_),
    .A2(_07901_));
 sg13g2_nor2b_1 _13709_ (.A(_07450_),
    .B_N(_07452_),
    .Y(_07910_));
 sg13g2_a221oi_1 _13710_ (.B2(_07888_),
    .C1(_07910_),
    .B1(_07909_),
    .A1(_07466_),
    .Y(_07911_),
    .A2(_07896_));
 sg13g2_o21ai_1 _13711_ (.B1(_07911_),
    .Y(_07912_),
    .A1(_07884_),
    .A2(_07889_));
 sg13g2_buf_2 _13712_ (.A(_07912_),
    .X(_07913_));
 sg13g2_nand2b_1 _13713_ (.Y(_07914_),
    .B(_07721_),
    .A_N(_07722_));
 sg13g2_nand2b_1 _13714_ (.Y(_07915_),
    .B(_07914_),
    .A_N(_07834_));
 sg13g2_buf_1 _13715_ (.A(_07915_),
    .X(_07916_));
 sg13g2_a221oi_1 _13716_ (.B2(_07913_),
    .C1(_07916_),
    .B1(_07845_),
    .A1(_07838_),
    .Y(_07917_),
    .A2(_07817_));
 sg13g2_and3_1 _13717_ (.X(_07918_),
    .A(_07913_),
    .B(_07845_),
    .C(_07916_));
 sg13g2_and2_1 _13718_ (.A(net807),
    .B(_07832_),
    .X(_07919_));
 sg13g2_o21ai_1 _13719_ (.B1(_07919_),
    .Y(_07920_),
    .A1(_07917_),
    .A2(_07918_));
 sg13g2_a21o_1 _13720_ (.A2(_07920_),
    .A1(_07840_),
    .B1(_07656_),
    .X(_07921_));
 sg13g2_buf_1 _13721_ (.A(_07921_),
    .X(_07922_));
 sg13g2_nand2_1 _13722_ (.Y(_07923_),
    .A(_07763_),
    .B(_07922_));
 sg13g2_o21ai_1 _13723_ (.B1(_07923_),
    .Y(_07924_),
    .A1(_07763_),
    .A2(net877));
 sg13g2_buf_2 _13724_ (.A(_00080_),
    .X(_07925_));
 sg13g2_buf_2 _13725_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[2] ),
    .X(_07926_));
 sg13g2_nand2_1 _13726_ (.Y(_07927_),
    .A(_07926_),
    .B(net877));
 sg13g2_buf_2 _13727_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[0] ),
    .X(_07928_));
 sg13g2_buf_1 _13728_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[1] ),
    .X(_07929_));
 sg13g2_nand2_1 _13729_ (.Y(_07930_),
    .A(_07928_),
    .B(_07929_));
 sg13g2_or3_1 _13730_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .B(_07927_),
    .C(_07930_),
    .X(_07931_));
 sg13g2_buf_1 _13731_ (.A(_07931_),
    .X(_07932_));
 sg13g2_a21o_1 _13732_ (.A2(_07932_),
    .A1(net1025),
    .B1(_07761_),
    .X(_07933_));
 sg13g2_buf_1 _13733_ (.A(\top_ihp.wb_uart.uart_rx.state[2] ),
    .X(_07934_));
 sg13g2_nor2_1 _13734_ (.A(_07761_),
    .B(_07934_),
    .Y(_07935_));
 sg13g2_buf_2 _13735_ (.A(ui_in[0]),
    .X(_07936_));
 sg13g2_inv_1 _13736_ (.Y(_07937_),
    .A(_07936_));
 sg13g2_nor2_1 _13737_ (.A(net1025),
    .B(_07937_),
    .Y(_07938_));
 sg13g2_a22oi_1 _13738_ (.Y(_07939_),
    .B1(_07935_),
    .B2(_07938_),
    .A2(_07933_),
    .A1(_07925_));
 sg13g2_a21oi_1 _13739_ (.A1(_07761_),
    .A2(_07924_),
    .Y(\top_ihp.wb_uart.uart_rx.next_state[0] ),
    .B1(_07939_));
 sg13g2_o21ai_1 _13740_ (.B1(_07925_),
    .Y(_07940_),
    .A1(_07761_),
    .A2(_07932_));
 sg13g2_nand3_1 _13741_ (.B(_07937_),
    .C(_07935_),
    .A(_07763_),
    .Y(_07941_));
 sg13g2_o21ai_1 _13742_ (.B1(_07941_),
    .Y(\top_ihp.wb_uart.uart_rx.next_state[1] ),
    .A1(_07763_),
    .A2(_07940_));
 sg13g2_nand3_1 _13743_ (.B(_07760_),
    .C(_07925_),
    .A(_07762_),
    .Y(_07942_));
 sg13g2_buf_1 _13744_ (.A(_07942_),
    .X(_07943_));
 sg13g2_nor2_1 _13745_ (.A(net1025),
    .B(_07760_),
    .Y(_07944_));
 sg13g2_nand2_1 _13746_ (.Y(_07945_),
    .A(_07934_),
    .B(_07944_));
 sg13g2_or2_1 _13747_ (.X(_07946_),
    .B(_07945_),
    .A(net877));
 sg13g2_o21ai_1 _13748_ (.B1(_07946_),
    .Y(\top_ihp.wb_uart.uart_rx.next_state[2] ),
    .A1(_07932_),
    .A2(_07943_));
 sg13g2_nor3_1 _13749_ (.A(net1025),
    .B(_07760_),
    .C(_07934_),
    .Y(_07947_));
 sg13g2_nor2b_1 _13750_ (.A(net877),
    .B_N(_07944_),
    .Y(_07948_));
 sg13g2_o21ai_1 _13751_ (.B1(_07922_),
    .Y(_07949_),
    .A1(_07947_),
    .A2(_07948_));
 sg13g2_nand2_1 _13752_ (.Y(_07950_),
    .A(_07760_),
    .B(net877));
 sg13g2_a21oi_1 _13753_ (.A1(_07925_),
    .A2(_07950_),
    .Y(_07951_),
    .B1(_07763_));
 sg13g2_nor3_1 _13754_ (.A(net1025),
    .B(_07761_),
    .C(_07936_),
    .Y(_07952_));
 sg13g2_nor3_1 _13755_ (.A(_07934_),
    .B(_07951_),
    .C(_07952_),
    .Y(_07953_));
 sg13g2_nor3_1 _13756_ (.A(_07763_),
    .B(_07760_),
    .C(net877),
    .Y(_07954_));
 sg13g2_nand2_1 _13757_ (.Y(_07955_),
    .A(_07953_),
    .B(_07954_));
 sg13g2_and3_1 _13758_ (.X(_07956_),
    .A(net1025),
    .B(_07925_),
    .C(_07932_));
 sg13g2_nor3_1 _13759_ (.A(net1025),
    .B(_07934_),
    .C(_07937_),
    .Y(_07957_));
 sg13g2_nor3_1 _13760_ (.A(_07761_),
    .B(_07956_),
    .C(_07957_),
    .Y(_07958_));
 sg13g2_a21oi_1 _13761_ (.A1(_07761_),
    .A2(_07925_),
    .Y(_07959_),
    .B1(_07958_));
 sg13g2_o21ai_1 _13762_ (.B1(_07959_),
    .Y(_07960_),
    .A1(_07953_),
    .A2(_07948_));
 sg13g2_and3_1 _13763_ (.X(_07961_),
    .A(_07949_),
    .B(_07955_),
    .C(_07960_));
 sg13g2_buf_1 _13764_ (.A(_07961_),
    .X(_07962_));
 sg13g2_buf_1 _13765_ (.A(_07962_),
    .X(_07963_));
 sg13g2_nor2_1 _13766_ (.A(_07785_),
    .B(net254),
    .Y(_00004_));
 sg13g2_xnor2_1 _13767_ (.Y(_07964_),
    .A(_07785_),
    .B(_07796_));
 sg13g2_nor2_1 _13768_ (.A(net254),
    .B(_07964_),
    .Y(_00015_));
 sg13g2_nand2_1 _13769_ (.Y(_07965_),
    .A(_07785_),
    .B(_07796_));
 sg13g2_xor2_1 _13770_ (.B(_07965_),
    .A(_07794_),
    .X(_07966_));
 sg13g2_nor2_1 _13771_ (.A(net254),
    .B(_07966_),
    .Y(_00026_));
 sg13g2_nand3_1 _13772_ (.B(_07796_),
    .C(_07794_),
    .A(_07785_),
    .Y(_07967_));
 sg13g2_xor2_1 _13773_ (.B(_07967_),
    .A(_07795_),
    .X(_07968_));
 sg13g2_nor2_1 _13774_ (.A(_07963_),
    .B(_07968_),
    .Y(_00029_));
 sg13g2_and4_1 _13775_ (.A(_07785_),
    .B(_07796_),
    .C(_07795_),
    .D(_07794_),
    .X(_07969_));
 sg13g2_buf_2 _13776_ (.A(_07969_),
    .X(_07970_));
 sg13g2_xnor2_1 _13777_ (.Y(_07971_),
    .A(_07789_),
    .B(_07970_));
 sg13g2_nor2_1 _13778_ (.A(net254),
    .B(_07971_),
    .Y(_00030_));
 sg13g2_nand2_1 _13779_ (.Y(_07972_),
    .A(_07789_),
    .B(_07970_));
 sg13g2_xnor2_1 _13780_ (.Y(_07973_),
    .A(_00079_),
    .B(_07972_));
 sg13g2_nor2_1 _13781_ (.A(net254),
    .B(_07973_),
    .Y(_00031_));
 sg13g2_nand3_1 _13782_ (.B(_07791_),
    .C(_07970_),
    .A(_07789_),
    .Y(_07974_));
 sg13g2_xnor2_1 _13783_ (.Y(_07975_),
    .A(_07788_),
    .B(_07974_));
 sg13g2_nor2_1 _13784_ (.A(net254),
    .B(_07975_),
    .Y(_00032_));
 sg13g2_inv_1 _13785_ (.Y(_07976_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ));
 sg13g2_nand4_1 _13786_ (.B(_07789_),
    .C(_07791_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ),
    .Y(_07977_),
    .D(_07970_));
 sg13g2_xnor2_1 _13787_ (.Y(_07978_),
    .A(_07976_),
    .B(_07977_));
 sg13g2_nor2_1 _13788_ (.A(net254),
    .B(_07978_),
    .Y(_00033_));
 sg13g2_nor2_2 _13789_ (.A(_07976_),
    .B(_07977_),
    .Y(_07979_));
 sg13g2_xnor2_1 _13790_ (.Y(_07980_),
    .A(_07787_),
    .B(_07979_));
 sg13g2_nor2_1 _13791_ (.A(net254),
    .B(_07980_),
    .Y(_00034_));
 sg13g2_nand2_1 _13792_ (.Y(_07981_),
    .A(_07787_),
    .B(_07979_));
 sg13g2_xor2_1 _13793_ (.B(_07981_),
    .A(_07781_),
    .X(_07982_));
 sg13g2_nor2_1 _13794_ (.A(_07963_),
    .B(_07982_),
    .Y(_00035_));
 sg13g2_buf_1 _13795_ (.A(_07962_),
    .X(_07983_));
 sg13g2_nand3_1 _13796_ (.B(_07781_),
    .C(_07979_),
    .A(_07787_),
    .Y(_07984_));
 sg13g2_xor2_1 _13797_ (.B(_07984_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .X(_07985_));
 sg13g2_nor2_1 _13798_ (.A(net253),
    .B(_07985_),
    .Y(_00005_));
 sg13g2_and4_1 _13799_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .B(_07787_),
    .C(_07781_),
    .D(_07979_),
    .X(_07986_));
 sg13g2_buf_1 _13800_ (.A(_07986_),
    .X(_07987_));
 sg13g2_xnor2_1 _13801_ (.Y(_07988_),
    .A(_07780_),
    .B(_07987_));
 sg13g2_nor2_1 _13802_ (.A(net253),
    .B(_07988_),
    .Y(_00006_));
 sg13g2_nand2_1 _13803_ (.Y(_07989_),
    .A(_07780_),
    .B(_07987_));
 sg13g2_xor2_1 _13804_ (.B(_07989_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .X(_07990_));
 sg13g2_nor2_1 _13805_ (.A(net253),
    .B(_07990_),
    .Y(_00007_));
 sg13g2_and3_1 _13806_ (.X(_07991_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .B(_07780_),
    .C(_07987_));
 sg13g2_buf_1 _13807_ (.A(_07991_),
    .X(_07992_));
 sg13g2_xnor2_1 _13808_ (.Y(_07993_),
    .A(_07766_),
    .B(_07992_));
 sg13g2_nor2_1 _13809_ (.A(_07983_),
    .B(_07993_),
    .Y(_00008_));
 sg13g2_nand2_1 _13810_ (.Y(_07994_),
    .A(_07766_),
    .B(_07992_));
 sg13g2_xor2_1 _13811_ (.B(_07994_),
    .A(_07765_),
    .X(_07995_));
 sg13g2_nor2_1 _13812_ (.A(_07983_),
    .B(_07995_),
    .Y(_00009_));
 sg13g2_nand3_1 _13813_ (.B(_07766_),
    .C(_07992_),
    .A(_07765_),
    .Y(_07996_));
 sg13g2_xor2_1 _13814_ (.B(_07996_),
    .A(_07764_),
    .X(_07997_));
 sg13g2_nor2_1 _13815_ (.A(net253),
    .B(_07997_),
    .Y(_00010_));
 sg13g2_inv_1 _13816_ (.Y(_07998_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ));
 sg13g2_nand4_1 _13817_ (.B(_07765_),
    .C(_07766_),
    .A(_07764_),
    .Y(_07999_),
    .D(_07992_));
 sg13g2_xnor2_1 _13818_ (.Y(_08000_),
    .A(_07998_),
    .B(_07999_));
 sg13g2_nor2_1 _13819_ (.A(net253),
    .B(_08000_),
    .Y(_00011_));
 sg13g2_nor2_1 _13820_ (.A(_07998_),
    .B(_07999_),
    .Y(_08001_));
 sg13g2_xnor2_1 _13821_ (.Y(_08002_),
    .A(_07770_),
    .B(_08001_));
 sg13g2_nor2_1 _13822_ (.A(net253),
    .B(_08002_),
    .Y(_00012_));
 sg13g2_and2_1 _13823_ (.A(_07770_),
    .B(_08001_),
    .X(_08003_));
 sg13g2_buf_1 _13824_ (.A(_08003_),
    .X(_08004_));
 sg13g2_xnor2_1 _13825_ (.Y(_08005_),
    .A(_07769_),
    .B(_08004_));
 sg13g2_nor2_1 _13826_ (.A(net253),
    .B(_08005_),
    .Y(_00013_));
 sg13g2_nand2_1 _13827_ (.Y(_08006_),
    .A(_07769_),
    .B(_08004_));
 sg13g2_xor2_1 _13828_ (.B(_08006_),
    .A(_07768_),
    .X(_08007_));
 sg13g2_nor2_1 _13829_ (.A(net253),
    .B(_08007_),
    .Y(_00014_));
 sg13g2_buf_1 _13830_ (.A(_07962_),
    .X(_08008_));
 sg13g2_nand3_1 _13831_ (.B(_07769_),
    .C(_08004_),
    .A(_07768_),
    .Y(_08009_));
 sg13g2_xor2_1 _13832_ (.B(_08009_),
    .A(_07773_),
    .X(_08010_));
 sg13g2_nor2_1 _13833_ (.A(net252),
    .B(_08010_),
    .Y(_00016_));
 sg13g2_nand4_1 _13834_ (.B(_07768_),
    .C(_07769_),
    .A(_07773_),
    .Y(_08011_),
    .D(_08004_));
 sg13g2_xor2_1 _13835_ (.B(_08011_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .X(_08012_));
 sg13g2_nor2_1 _13836_ (.A(net252),
    .B(_08012_),
    .Y(_00017_));
 sg13g2_nand3_1 _13837_ (.B(_07768_),
    .C(_07769_),
    .A(_07773_),
    .Y(_08013_));
 sg13g2_nand2_1 _13838_ (.Y(_08014_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .B(_07770_));
 sg13g2_nor2_1 _13839_ (.A(_08013_),
    .B(_08014_),
    .Y(_08015_));
 sg13g2_nand2_1 _13840_ (.Y(_08016_),
    .A(_08001_),
    .B(_08015_));
 sg13g2_xor2_1 _13841_ (.B(_08016_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .X(_08017_));
 sg13g2_nor2_1 _13842_ (.A(net252),
    .B(_08017_),
    .Y(_00018_));
 sg13g2_and4_1 _13843_ (.A(_07764_),
    .B(_07765_),
    .C(_07766_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ),
    .X(_08018_));
 sg13g2_and4_1 _13844_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .B(_07992_),
    .C(_08015_),
    .D(_08018_),
    .X(_08019_));
 sg13g2_buf_1 _13845_ (.A(_08019_),
    .X(_08020_));
 sg13g2_xnor2_1 _13846_ (.Y(_08021_),
    .A(_07772_),
    .B(_08020_));
 sg13g2_nor2_1 _13847_ (.A(net252),
    .B(_08021_),
    .Y(_00019_));
 sg13g2_nand2_1 _13848_ (.Y(_08022_),
    .A(_07772_),
    .B(_08020_));
 sg13g2_xor2_1 _13849_ (.B(_08022_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ),
    .X(_08023_));
 sg13g2_nor2_1 _13850_ (.A(net252),
    .B(_08023_),
    .Y(_00020_));
 sg13g2_and3_1 _13851_ (.X(_08024_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ),
    .B(_07772_),
    .C(_08020_));
 sg13g2_buf_1 _13852_ (.A(_08024_),
    .X(_08025_));
 sg13g2_xnor2_1 _13853_ (.Y(_08026_),
    .A(_07775_),
    .B(_08025_));
 sg13g2_nor2_1 _13854_ (.A(_08008_),
    .B(_08026_),
    .Y(_00021_));
 sg13g2_nand2_1 _13855_ (.Y(_08027_),
    .A(_07775_),
    .B(_08025_));
 sg13g2_xor2_1 _13856_ (.B(_08027_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .X(_08028_));
 sg13g2_nor2_1 _13857_ (.A(net252),
    .B(_08028_),
    .Y(_00022_));
 sg13g2_inv_1 _13858_ (.Y(_08029_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ));
 sg13g2_nand3_1 _13859_ (.B(_07775_),
    .C(_08025_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .Y(_08030_));
 sg13g2_xnor2_1 _13860_ (.Y(_08031_),
    .A(_08029_),
    .B(_08030_));
 sg13g2_nor2_1 _13861_ (.A(net252),
    .B(_08031_),
    .Y(_00023_));
 sg13g2_nor2_2 _13862_ (.A(_08029_),
    .B(_08030_),
    .Y(_08032_));
 sg13g2_xnor2_1 _13863_ (.Y(_08033_),
    .A(_07782_),
    .B(_08032_));
 sg13g2_nor2_1 _13864_ (.A(_08008_),
    .B(_08033_),
    .Y(_00024_));
 sg13g2_nand2_1 _13865_ (.Y(_08034_),
    .A(_07782_),
    .B(_08032_));
 sg13g2_xor2_1 _13866_ (.B(_08034_),
    .A(_07778_),
    .X(_08035_));
 sg13g2_nor2_1 _13867_ (.A(net252),
    .B(_08035_),
    .Y(_00025_));
 sg13g2_and3_1 _13868_ (.X(_08036_),
    .A(_07778_),
    .B(_07782_),
    .C(_08032_));
 sg13g2_xnor2_1 _13869_ (.Y(_08037_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .B(_08036_));
 sg13g2_nor2_1 _13870_ (.A(_07962_),
    .B(_08037_),
    .Y(_00027_));
 sg13g2_nand4_1 _13871_ (.B(_07778_),
    .C(_07782_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .Y(_08038_),
    .D(_08032_));
 sg13g2_xor2_1 _13872_ (.B(_08038_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ),
    .X(_08039_));
 sg13g2_nor2_1 _13873_ (.A(_07962_),
    .B(_08039_),
    .Y(_00028_));
 sg13g2_buf_2 _13874_ (.A(\top_ihp.wb_uart.uart_tx.state[0] ),
    .X(_08040_));
 sg13g2_inv_1 _13875_ (.Y(_08041_),
    .A(_08040_));
 sg13g2_buf_1 _13876_ (.A(\top_ihp.wb_uart.uart_tx.state[1] ),
    .X(_08042_));
 sg13g2_buf_2 _13877_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[0] ),
    .X(_08043_));
 sg13g2_buf_2 _13878_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[1] ),
    .X(_08044_));
 sg13g2_buf_2 _13879_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ),
    .X(_08045_));
 sg13g2_nor4_1 _13880_ (.A(_08045_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ),
    .Y(_08046_));
 sg13g2_buf_1 _13881_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ),
    .X(_08047_));
 sg13g2_buf_1 _13882_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ),
    .X(_08048_));
 sg13g2_buf_1 _13883_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[23] ),
    .X(_08049_));
 sg13g2_nor4_1 _13884_ (.A(_08047_),
    .B(_08048_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .D(_08049_),
    .Y(_08050_));
 sg13g2_buf_1 _13885_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ),
    .X(_08051_));
 sg13g2_buf_1 _13886_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ),
    .X(_08052_));
 sg13g2_buf_1 _13887_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[28] ),
    .X(_08053_));
 sg13g2_nor4_1 _13888_ (.A(_08051_),
    .B(_08052_),
    .C(_08053_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ),
    .Y(_08054_));
 sg13g2_buf_8 _13889_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[0] ),
    .X(_08055_));
 sg13g2_buf_8 _13890_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[1] ),
    .X(_08056_));
 sg13g2_inv_1 _13891_ (.Y(_08057_),
    .A(_08056_));
 sg13g2_buf_1 _13892_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[24] ),
    .X(_08058_));
 sg13g2_nor4_1 _13893_ (.A(_08055_),
    .B(_08057_),
    .C(_08058_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .Y(_08059_));
 sg13g2_nand4_1 _13894_ (.B(_08050_),
    .C(_08054_),
    .A(_08046_),
    .Y(_08060_),
    .D(_08059_));
 sg13g2_buf_1 _13895_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[9] ),
    .X(_08061_));
 sg13g2_inv_1 _13896_ (.Y(_08062_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ));
 sg13g2_buf_1 _13897_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .X(_08063_));
 sg13g2_buf_1 _13898_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ),
    .X(_08064_));
 sg13g2_nor4_1 _13899_ (.A(_08061_),
    .B(_08062_),
    .C(_08063_),
    .D(_08064_),
    .Y(_08065_));
 sg13g2_buf_8 _13900_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ),
    .X(_08066_));
 sg13g2_buf_1 _13901_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[6] ),
    .X(_08067_));
 sg13g2_inv_1 _13902_ (.Y(_08068_),
    .A(_08067_));
 sg13g2_nor4_1 _13903_ (.A(_08066_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .D(_08068_),
    .Y(_08069_));
 sg13g2_buf_1 _13904_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ),
    .X(_08070_));
 sg13g2_buf_1 _13905_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ),
    .X(_08071_));
 sg13g2_buf_2 _13906_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ),
    .X(_08072_));
 sg13g2_nor4_1 _13907_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ),
    .B(_08070_),
    .C(_08071_),
    .D(_08072_),
    .Y(_08073_));
 sg13g2_buf_1 _13908_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[3] ),
    .X(_08074_));
 sg13g2_nand2_1 _13909_ (.Y(_08075_),
    .A(_08074_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_nor3_1 _13910_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ),
    .C(_08075_),
    .Y(_08076_));
 sg13g2_nand4_1 _13911_ (.B(_08069_),
    .C(_08073_),
    .A(_08065_),
    .Y(_08077_),
    .D(_08076_));
 sg13g2_nor2_1 _13912_ (.A(_08060_),
    .B(_08077_),
    .Y(_08078_));
 sg13g2_buf_1 _13913_ (.A(_08078_),
    .X(_08079_));
 sg13g2_nand4_1 _13914_ (.B(_08044_),
    .C(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .A(_08043_),
    .Y(_08080_),
    .D(_08079_));
 sg13g2_nor2_1 _13915_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ),
    .B(_08080_),
    .Y(_08081_));
 sg13g2_a21o_1 _13916_ (.A2(_07920_),
    .A1(_07840_),
    .B1(_07673_),
    .X(_08082_));
 sg13g2_buf_2 _13917_ (.A(_08082_),
    .X(_08083_));
 sg13g2_nor2_1 _13918_ (.A(net1024),
    .B(_08083_),
    .Y(_08084_));
 sg13g2_a21oi_1 _13919_ (.A1(net1024),
    .A2(_08081_),
    .Y(_08085_),
    .B1(_08084_));
 sg13g2_nand2_1 _13920_ (.Y(_08086_),
    .A(_08040_),
    .B(_08079_));
 sg13g2_inv_1 _13921_ (.Y(_08087_),
    .A(_08086_));
 sg13g2_a21oi_1 _13922_ (.A1(_08041_),
    .A2(_08085_),
    .Y(\top_ihp.wb_uart.uart_tx.next_state[0] ),
    .B1(_08087_));
 sg13g2_xnor2_1 _13923_ (.Y(\top_ihp.wb_uart.uart_tx.next_state[1] ),
    .A(net1024),
    .B(_08086_));
 sg13g2_o21ai_1 _13924_ (.B1(_08079_),
    .Y(_08088_),
    .A1(net1024),
    .A2(_08040_));
 sg13g2_or3_1 _13925_ (.A(_08042_),
    .B(_08040_),
    .C(_08083_),
    .X(_08089_));
 sg13g2_buf_2 _13926_ (.A(_08089_),
    .X(_08090_));
 sg13g2_nand2_1 _13927_ (.Y(_08091_),
    .A(_08088_),
    .B(net551));
 sg13g2_buf_8 _13928_ (.A(_08091_),
    .X(_08092_));
 sg13g2_buf_1 _13929_ (.A(_08092_),
    .X(_08093_));
 sg13g2_nor2_1 _13930_ (.A(_08055_),
    .B(net151),
    .Y(_00036_));
 sg13g2_xnor2_1 _13931_ (.Y(_08094_),
    .A(_08055_),
    .B(_08056_));
 sg13g2_nor2_1 _13932_ (.A(net151),
    .B(_08094_),
    .Y(_00047_));
 sg13g2_nand2_1 _13933_ (.Y(_08095_),
    .A(_08055_),
    .B(_08056_));
 sg13g2_xor2_1 _13934_ (.B(_08095_),
    .A(_08066_),
    .X(_08096_));
 sg13g2_nor2_1 _13935_ (.A(net151),
    .B(_08096_),
    .Y(_00058_));
 sg13g2_nand3_1 _13936_ (.B(_08056_),
    .C(_08066_),
    .A(_08055_),
    .Y(_08097_));
 sg13g2_buf_2 _13937_ (.A(_08097_),
    .X(_08098_));
 sg13g2_xor2_1 _13938_ (.B(_08098_),
    .A(_08074_),
    .X(_08099_));
 sg13g2_nor2_1 _13939_ (.A(net151),
    .B(_08099_),
    .Y(_00061_));
 sg13g2_nand4_1 _13940_ (.B(_08056_),
    .C(_08066_),
    .A(_08055_),
    .Y(_08100_),
    .D(_08074_));
 sg13g2_xor2_1 _13941_ (.B(_08100_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ),
    .X(_08101_));
 sg13g2_nor2_1 _13942_ (.A(net151),
    .B(_08101_),
    .Y(_00062_));
 sg13g2_nor2_1 _13943_ (.A(_08075_),
    .B(_08098_),
    .Y(_08102_));
 sg13g2_xnor2_1 _13944_ (.Y(_08103_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .B(_08102_));
 sg13g2_nor2_1 _13945_ (.A(_08093_),
    .B(_08103_),
    .Y(_00063_));
 sg13g2_nand3_1 _13946_ (.B(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ),
    .A(_08074_),
    .Y(_08104_));
 sg13g2_buf_1 _13947_ (.A(_08104_),
    .X(_08105_));
 sg13g2_nor2_1 _13948_ (.A(_08098_),
    .B(_08105_),
    .Y(_08106_));
 sg13g2_xnor2_1 _13949_ (.Y(_08107_),
    .A(_08067_),
    .B(_08106_));
 sg13g2_nor2_1 _13950_ (.A(net151),
    .B(_08107_),
    .Y(_00064_));
 sg13g2_nand2_1 _13951_ (.Y(_08108_),
    .A(_08067_),
    .B(_08106_));
 sg13g2_xor2_1 _13952_ (.B(_08108_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .X(_08109_));
 sg13g2_nor2_1 _13953_ (.A(_08093_),
    .B(_08109_),
    .Y(_00065_));
 sg13g2_nand2_1 _13954_ (.Y(_08110_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .B(_08067_));
 sg13g2_nor3_1 _13955_ (.A(_08098_),
    .B(_08105_),
    .C(_08110_),
    .Y(_08111_));
 sg13g2_xnor2_1 _13956_ (.Y(_08112_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ),
    .B(_08111_));
 sg13g2_nor2_1 _13957_ (.A(net151),
    .B(_08112_),
    .Y(_00066_));
 sg13g2_nor4_2 _13958_ (.A(_08062_),
    .B(_08098_),
    .C(_08105_),
    .Y(_08113_),
    .D(_08110_));
 sg13g2_xnor2_1 _13959_ (.Y(_08114_),
    .A(_08061_),
    .B(_08113_));
 sg13g2_nor2_1 _13960_ (.A(net151),
    .B(_08114_),
    .Y(_00067_));
 sg13g2_buf_1 _13961_ (.A(_08092_),
    .X(_08115_));
 sg13g2_and2_1 _13962_ (.A(_08061_),
    .B(_08113_),
    .X(_08116_));
 sg13g2_xnor2_1 _13963_ (.Y(_08117_),
    .A(_08063_),
    .B(_08116_));
 sg13g2_nor2_1 _13964_ (.A(net150),
    .B(_08117_),
    .Y(_00037_));
 sg13g2_nand2_1 _13965_ (.Y(_08118_),
    .A(_08063_),
    .B(_08116_));
 sg13g2_xor2_1 _13966_ (.B(_08118_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ),
    .X(_08119_));
 sg13g2_nor2_1 _13967_ (.A(net150),
    .B(_08119_),
    .Y(_00038_));
 sg13g2_and4_1 _13968_ (.A(_08061_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ),
    .C(_08063_),
    .D(_08113_),
    .X(_08120_));
 sg13g2_buf_1 _13969_ (.A(_08120_),
    .X(_08121_));
 sg13g2_xnor2_1 _13970_ (.Y(_08122_),
    .A(_08070_),
    .B(_08121_));
 sg13g2_nor2_1 _13971_ (.A(net150),
    .B(_08122_),
    .Y(_00039_));
 sg13g2_nand2_1 _13972_ (.Y(_08123_),
    .A(_08070_),
    .B(_08121_));
 sg13g2_xor2_1 _13973_ (.B(_08123_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ),
    .X(_08124_));
 sg13g2_nor2_1 _13974_ (.A(net150),
    .B(_08124_),
    .Y(_00040_));
 sg13g2_and3_1 _13975_ (.X(_08125_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ),
    .B(_08070_),
    .C(_08121_));
 sg13g2_buf_1 _13976_ (.A(_08125_),
    .X(_08126_));
 sg13g2_xnor2_1 _13977_ (.Y(_08127_),
    .A(_08072_),
    .B(_08126_));
 sg13g2_nor2_1 _13978_ (.A(net150),
    .B(_08127_),
    .Y(_00041_));
 sg13g2_nand2_1 _13979_ (.Y(_08128_),
    .A(_08072_),
    .B(_08126_));
 sg13g2_xor2_1 _13980_ (.B(_08128_),
    .A(_08071_),
    .X(_08129_));
 sg13g2_nor2_1 _13981_ (.A(net150),
    .B(_08129_),
    .Y(_00042_));
 sg13g2_nand3_1 _13982_ (.B(_08072_),
    .C(_08126_),
    .A(_08071_),
    .Y(_08130_));
 sg13g2_xor2_1 _13983_ (.B(_08130_),
    .A(_08064_),
    .X(_08131_));
 sg13g2_nor2_1 _13984_ (.A(_08115_),
    .B(_08131_),
    .Y(_00043_));
 sg13g2_nand4_1 _13985_ (.B(_08072_),
    .C(_08064_),
    .A(_08071_),
    .Y(_08132_),
    .D(_08126_));
 sg13g2_xor2_1 _13986_ (.B(_08132_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ),
    .X(_08133_));
 sg13g2_nor2_1 _13987_ (.A(net150),
    .B(_08133_),
    .Y(_00044_));
 sg13g2_and4_1 _13988_ (.A(_08071_),
    .B(_08072_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ),
    .D(_08064_),
    .X(_08134_));
 sg13g2_and2_1 _13989_ (.A(_08126_),
    .B(_08134_),
    .X(_08135_));
 sg13g2_buf_8 _13990_ (.A(_08135_),
    .X(_08136_));
 sg13g2_xnor2_1 _13991_ (.Y(_08137_),
    .A(_08047_),
    .B(_08136_));
 sg13g2_nor2_1 _13992_ (.A(net150),
    .B(_08137_),
    .Y(_00045_));
 sg13g2_nand2_1 _13993_ (.Y(_08138_),
    .A(_08047_),
    .B(_08136_));
 sg13g2_xor2_1 _13994_ (.B(_08138_),
    .A(_08045_),
    .X(_08139_));
 sg13g2_nor2_1 _13995_ (.A(_08115_),
    .B(_08139_),
    .Y(_00046_));
 sg13g2_buf_1 _13996_ (.A(_08092_),
    .X(_08140_));
 sg13g2_nand3_1 _13997_ (.B(_08047_),
    .C(_08136_),
    .A(_08045_),
    .Y(_08141_));
 sg13g2_xor2_1 _13998_ (.B(_08141_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .X(_08142_));
 sg13g2_nor2_1 _13999_ (.A(_08140_),
    .B(_08142_),
    .Y(_00048_));
 sg13g2_and4_1 _14000_ (.A(_08045_),
    .B(_08047_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .D(_08136_),
    .X(_08143_));
 sg13g2_buf_1 _14001_ (.A(_08143_),
    .X(_08144_));
 sg13g2_xnor2_1 _14002_ (.Y(_08145_),
    .A(_08048_),
    .B(_08144_));
 sg13g2_nor2_1 _14003_ (.A(net149),
    .B(_08145_),
    .Y(_00049_));
 sg13g2_nand2_1 _14004_ (.Y(_08146_),
    .A(_08048_),
    .B(_08144_));
 sg13g2_xor2_1 _14005_ (.B(_08146_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .X(_08147_));
 sg13g2_nor2_1 _14006_ (.A(_08140_),
    .B(_08147_),
    .Y(_00050_));
 sg13g2_and3_1 _14007_ (.X(_08148_),
    .A(_08048_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .C(_08144_));
 sg13g2_buf_1 _14008_ (.A(_08148_),
    .X(_08149_));
 sg13g2_xnor2_1 _14009_ (.Y(_08150_),
    .A(_08049_),
    .B(_08149_));
 sg13g2_nor2_1 _14010_ (.A(net149),
    .B(_08150_),
    .Y(_00051_));
 sg13g2_nand2_1 _14011_ (.Y(_08151_),
    .A(_08049_),
    .B(_08149_));
 sg13g2_xor2_1 _14012_ (.B(_08151_),
    .A(_08058_),
    .X(_08152_));
 sg13g2_nor2_1 _14013_ (.A(net149),
    .B(_08152_),
    .Y(_00052_));
 sg13g2_nand3_1 _14014_ (.B(_08058_),
    .C(_08149_),
    .A(_08049_),
    .Y(_08153_));
 sg13g2_xor2_1 _14015_ (.B(_08153_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ),
    .X(_08154_));
 sg13g2_nor2_1 _14016_ (.A(net149),
    .B(_08154_),
    .Y(_00053_));
 sg13g2_and4_1 _14017_ (.A(_08049_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ),
    .C(_08058_),
    .D(_08149_),
    .X(_08155_));
 sg13g2_buf_1 _14018_ (.A(_08155_),
    .X(_08156_));
 sg13g2_xnor2_1 _14019_ (.Y(_08157_),
    .A(_08051_),
    .B(_08156_));
 sg13g2_nor2_1 _14020_ (.A(net149),
    .B(_08157_),
    .Y(_00054_));
 sg13g2_nand2_1 _14021_ (.Y(_08158_),
    .A(_08051_),
    .B(_08156_));
 sg13g2_xor2_1 _14022_ (.B(_08158_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ),
    .X(_08159_));
 sg13g2_nor2_1 _14023_ (.A(net149),
    .B(_08159_),
    .Y(_00055_));
 sg13g2_and3_1 _14024_ (.X(_08160_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ),
    .B(_08051_),
    .C(_08156_));
 sg13g2_buf_1 _14025_ (.A(_08160_),
    .X(_08161_));
 sg13g2_xnor2_1 _14026_ (.Y(_08162_),
    .A(_08053_),
    .B(_08161_));
 sg13g2_nor2_1 _14027_ (.A(net149),
    .B(_08162_),
    .Y(_00056_));
 sg13g2_nand2_1 _14028_ (.Y(_08163_),
    .A(_08053_),
    .B(_08161_));
 sg13g2_xor2_1 _14029_ (.B(_08163_),
    .A(_08052_),
    .X(_08164_));
 sg13g2_nor2_1 _14030_ (.A(net149),
    .B(_08164_),
    .Y(_00057_));
 sg13g2_nand3_1 _14031_ (.B(_08053_),
    .C(_08161_),
    .A(_08052_),
    .Y(_08165_));
 sg13g2_xor2_1 _14032_ (.B(_08165_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .X(_08166_));
 sg13g2_nor2_1 _14033_ (.A(_08092_),
    .B(_08166_),
    .Y(_00059_));
 sg13g2_nand4_1 _14034_ (.B(_08053_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .A(_08052_),
    .Y(_08167_),
    .D(_08161_));
 sg13g2_xor2_1 _14035_ (.B(_08167_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ),
    .X(_08168_));
 sg13g2_nor2_1 _14036_ (.A(_08092_),
    .B(_08168_),
    .Y(_00060_));
 sg13g2_buf_1 _14037_ (.A(net984),
    .X(_08169_));
 sg13g2_o21ai_1 _14038_ (.B1(net940),
    .Y(_08170_),
    .A1(_07474_),
    .A2(_07438_));
 sg13g2_nor2b_1 _14039_ (.A(_07475_),
    .B_N(_07474_),
    .Y(_08171_));
 sg13g2_a22oi_1 _14040_ (.Y(_08172_),
    .B1(_08171_),
    .B2(net807),
    .A2(_08170_),
    .A1(_07475_));
 sg13g2_buf_2 _14041_ (.A(_08172_),
    .X(_08173_));
 sg13g2_inv_1 _14042_ (.Y(\top_ihp.oisc.wb_adr_o[0] ),
    .A(_08173_));
 sg13g2_xnor2_1 _14043_ (.Y(_08174_),
    .A(_07477_),
    .B(_07848_));
 sg13g2_a21o_1 _14044_ (.A2(_08174_),
    .A1(net807),
    .B1(net982),
    .X(_08175_));
 sg13g2_nor2_1 _14045_ (.A(net1041),
    .B(_08174_),
    .Y(_08176_));
 sg13g2_a22oi_1 _14046_ (.Y(_08177_),
    .B1(_08176_),
    .B2(net807),
    .A2(_08175_),
    .A1(net1041));
 sg13g2_buf_2 _14047_ (.A(_08177_),
    .X(_08178_));
 sg13g2_inv_1 _14048_ (.Y(\top_ihp.oisc.wb_adr_o[1] ),
    .A(_08178_));
 sg13g2_buf_2 _14049_ (.A(\top_ihp.wb_imem.state[1] ),
    .X(_08179_));
 sg13g2_buf_1 _14050_ (.A(\top_ihp.wb_emem.last_bit ),
    .X(_08180_));
 sg13g2_buf_2 _14051_ (.A(\top_ihp.wb_emem.state[2] ),
    .X(_08181_));
 sg13g2_buf_2 _14052_ (.A(\top_ihp.wb_emem.state[3] ),
    .X(_08182_));
 sg13g2_nor2_1 _14053_ (.A(_08181_),
    .B(_08182_),
    .Y(_08183_));
 sg13g2_buf_2 _14054_ (.A(_08183_),
    .X(_08184_));
 sg13g2_buf_1 _14055_ (.A(\top_ihp.wb_emem.state[1] ),
    .X(_08185_));
 sg13g2_buf_1 _14056_ (.A(\top_ihp.wb_emem.state[0] ),
    .X(_08186_));
 sg13g2_and2_1 _14057_ (.A(_08185_),
    .B(net1013),
    .X(_08187_));
 sg13g2_buf_2 _14058_ (.A(_08187_),
    .X(_08188_));
 sg13g2_nand3_1 _14059_ (.B(_08184_),
    .C(_08188_),
    .A(_08180_),
    .Y(_08189_));
 sg13g2_buf_2 _14060_ (.A(_08189_),
    .X(_08190_));
 sg13g2_buf_2 _14061_ (.A(\top_ihp.wb_ack_spi ),
    .X(_08191_));
 sg13g2_and2_1 _14062_ (.A(_08191_),
    .B(\top_ihp.wb_dati_spi[15] ),
    .X(_08192_));
 sg13g2_inv_1 _14063_ (.Y(_08193_),
    .A(_08180_));
 sg13g2_buf_1 _14064_ (.A(_08193_),
    .X(_08194_));
 sg13g2_inv_1 _14065_ (.Y(_08195_),
    .A(\top_ihp.wb_dati_ram[15] ));
 sg13g2_or2_1 _14066_ (.X(_08196_),
    .B(_08182_),
    .A(_08181_));
 sg13g2_buf_2 _14067_ (.A(_08196_),
    .X(_08197_));
 sg13g2_nand2_1 _14068_ (.Y(_08198_),
    .A(_08185_),
    .B(net1013));
 sg13g2_buf_1 _14069_ (.A(_08198_),
    .X(_08199_));
 sg13g2_buf_1 _14070_ (.A(_08199_),
    .X(_08200_));
 sg13g2_nor4_1 _14071_ (.A(net981),
    .B(_08195_),
    .C(_08197_),
    .D(net903),
    .Y(_08201_));
 sg13g2_a221oi_1 _14072_ (.B2(_08192_),
    .C1(_08201_),
    .B1(_08190_),
    .A1(_08179_),
    .Y(_08202_),
    .A2(net878));
 sg13g2_buf_1 _14073_ (.A(_08202_),
    .X(_08203_));
 sg13g2_nand3_1 _14074_ (.B(_07744_),
    .C(_07754_),
    .A(_08179_),
    .Y(_08204_));
 sg13g2_buf_2 _14075_ (.A(_08204_),
    .X(_08205_));
 sg13g2_buf_8 _14076_ (.A(_08205_),
    .X(_08206_));
 sg13g2_and2_1 _14077_ (.A(_00072_),
    .B(_00071_),
    .X(_08207_));
 sg13g2_buf_1 _14078_ (.A(_08207_),
    .X(_08208_));
 sg13g2_o21ai_1 _14079_ (.B1(_08208_),
    .Y(_08209_),
    .A1(\top_ihp.wb_dati_rom[15] ),
    .A2(net862));
 sg13g2_or2_1 _14080_ (.X(_08210_),
    .B(_08209_),
    .A(_08203_));
 sg13g2_buf_1 _14081_ (.A(_08191_),
    .X(_08211_));
 sg13g2_and3_1 _14082_ (.X(_08212_),
    .A(_08179_),
    .B(_07744_),
    .C(_07754_));
 sg13g2_buf_8 _14083_ (.A(_08212_),
    .X(_08213_));
 sg13g2_nor3_1 _14084_ (.A(_08193_),
    .B(_08197_),
    .C(_08199_),
    .Y(_08214_));
 sg13g2_buf_1 _14085_ (.A(\top_ihp.wb_ack_uart ),
    .X(_08215_));
 sg13g2_buf_1 _14086_ (.A(\top_ihp.wb_ack_gpio ),
    .X(_08216_));
 sg13g2_or2_1 _14087_ (.X(_08217_),
    .B(_08216_),
    .A(_08215_));
 sg13g2_buf_1 _14088_ (.A(_08217_),
    .X(_08218_));
 sg13g2_or4_1 _14089_ (.A(_08211_),
    .B(_08213_),
    .C(_08214_),
    .D(net980),
    .X(_08219_));
 sg13g2_buf_8 _14090_ (.A(_08219_),
    .X(_08220_));
 sg13g2_nand2_1 _14091_ (.Y(_08221_),
    .A(net1017),
    .B(net845));
 sg13g2_buf_1 _14092_ (.A(_08221_),
    .X(_08222_));
 sg13g2_buf_1 _14093_ (.A(net805),
    .X(_08223_));
 sg13g2_buf_1 _14094_ (.A(net776),
    .X(_08224_));
 sg13g2_buf_1 _14095_ (.A(net805),
    .X(_08225_));
 sg13g2_nand2_1 _14096_ (.Y(_08226_),
    .A(\top_ihp.oisc.decoder.instruction[15] ),
    .B(net775));
 sg13g2_o21ai_1 _14097_ (.B1(_08226_),
    .Y(_00107_),
    .A1(_08210_),
    .A2(net738));
 sg13g2_buf_1 _14098_ (.A(\top_ihp.oisc.micro_op[9] ),
    .X(_08227_));
 sg13g2_buf_1 _14099_ (.A(\top_ihp.oisc.micro_state[1] ),
    .X(_08228_));
 sg13g2_and2_1 _14100_ (.A(_08228_),
    .B(net1016),
    .X(_08229_));
 sg13g2_buf_1 _14101_ (.A(_08229_),
    .X(_08230_));
 sg13g2_nand2_1 _14102_ (.Y(_08231_),
    .A(_08227_),
    .B(net939));
 sg13g2_inv_1 _14103_ (.Y(\top_ihp.oisc.reg_rb[1] ),
    .A(_08231_));
 sg13g2_buf_1 _14104_ (.A(\top_ihp.oisc.micro_op[8] ),
    .X(_08232_));
 sg13g2_nand2_1 _14105_ (.Y(_08233_),
    .A(_08232_),
    .B(net939));
 sg13g2_inv_1 _14106_ (.Y(\top_ihp.oisc.reg_rb[0] ),
    .A(_08233_));
 sg13g2_nand2_1 _14107_ (.Y(_08234_),
    .A(\top_ihp.oisc.micro_op[11] ),
    .B(_08230_));
 sg13g2_buf_2 _14108_ (.A(_08234_),
    .X(_08235_));
 sg13g2_inv_1 _14109_ (.Y(\top_ihp.oisc.reg_rb[3] ),
    .A(_08235_));
 sg13g2_nand2_1 _14110_ (.Y(_08236_),
    .A(_07428_),
    .B(_07433_));
 sg13g2_buf_2 _14111_ (.A(_08236_),
    .X(_08237_));
 sg13g2_buf_2 _14112_ (.A(\top_ihp.oisc.micro_op[10] ),
    .X(_08238_));
 sg13g2_nand2_1 _14113_ (.Y(_08239_),
    .A(_08238_),
    .B(net939));
 sg13g2_o21ai_1 _14114_ (.B1(_08239_),
    .Y(_08240_),
    .A1(_08237_),
    .A2(net939));
 sg13g2_buf_1 _14115_ (.A(_08240_),
    .X(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_buf_2 _14116_ (.A(\top_ihp.oisc.state[6] ),
    .X(_08241_));
 sg13g2_nor4_1 _14117_ (.A(_08191_),
    .B(_08213_),
    .C(_08214_),
    .D(net980),
    .Y(_08242_));
 sg13g2_buf_2 _14118_ (.A(_08242_),
    .X(_08243_));
 sg13g2_buf_8 _14119_ (.A(_08243_),
    .X(_08244_));
 sg13g2_o21ai_1 _14120_ (.B1(_08244_),
    .Y(_08245_),
    .A1(net982),
    .A2(_08241_));
 sg13g2_buf_1 _14121_ (.A(_08245_),
    .X(_08246_));
 sg13g2_buf_1 _14122_ (.A(net1016),
    .X(_08247_));
 sg13g2_nor2_1 _14123_ (.A(net979),
    .B(_00076_),
    .Y(_08248_));
 sg13g2_and2_1 _14124_ (.A(_07423_),
    .B(_08237_),
    .X(_08249_));
 sg13g2_buf_1 _14125_ (.A(_08249_),
    .X(_08250_));
 sg13g2_a21o_1 _14126_ (.A2(_08248_),
    .A1(net774),
    .B1(_08250_),
    .X(_00002_));
 sg13g2_xor2_1 _14127_ (.B(\top_ihp.wb_spi.spi_clk_cnt[0] ),
    .A(\top_ihp.spi_clk_o ),
    .X(_00140_));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_nand2_1 _14129_ (.Y(_08251_),
    .A(net1016),
    .B(\top_ihp.oisc.micro_state[0] ));
 sg13g2_and2_1 _14130_ (.A(_08237_),
    .B(_08251_),
    .X(_08252_));
 sg13g2_buf_1 _14131_ (.A(_08252_),
    .X(_08253_));
 sg13g2_buf_1 _14132_ (.A(_08253_),
    .X(_08254_));
 sg13g2_buf_1 _14133_ (.A(\top_ihp.oisc.micro_pc[7] ),
    .X(_08255_));
 sg13g2_inv_1 _14134_ (.Y(_08256_),
    .A(_08255_));
 sg13g2_buf_1 _14135_ (.A(_08256_),
    .X(_08257_));
 sg13g2_buf_1 _14136_ (.A(\top_ihp.oisc.micro_pc[6] ),
    .X(_08258_));
 sg13g2_inv_1 _14137_ (.Y(_08259_),
    .A(net1023));
 sg13g2_buf_1 _14138_ (.A(_08259_),
    .X(_08260_));
 sg13g2_buf_1 _14139_ (.A(_00085_),
    .X(_08261_));
 sg13g2_buf_1 _14140_ (.A(net1022),
    .X(_08262_));
 sg13g2_buf_2 _14141_ (.A(_00083_),
    .X(_08263_));
 sg13g2_buf_2 _14142_ (.A(\top_ihp.oisc.micro_pc[0] ),
    .X(_08264_));
 sg13g2_buf_1 _14143_ (.A(_08264_),
    .X(_08265_));
 sg13g2_buf_1 _14144_ (.A(net1010),
    .X(_08266_));
 sg13g2_buf_1 _14145_ (.A(net976),
    .X(_08267_));
 sg13g2_buf_1 _14146_ (.A(_08267_),
    .X(_08268_));
 sg13g2_buf_1 _14147_ (.A(\top_ihp.oisc.micro_pc[1] ),
    .X(_08269_));
 sg13g2_buf_1 _14148_ (.A(net1021),
    .X(_08270_));
 sg13g2_buf_1 _14149_ (.A(net1009),
    .X(_08271_));
 sg13g2_buf_1 _14150_ (.A(net975),
    .X(_08272_));
 sg13g2_buf_1 _14151_ (.A(net937),
    .X(_08273_));
 sg13g2_buf_1 _14152_ (.A(_00086_),
    .X(_08274_));
 sg13g2_buf_1 _14153_ (.A(\top_ihp.oisc.micro_pc[4] ),
    .X(_08275_));
 sg13g2_inv_1 _14154_ (.Y(_08276_),
    .A(_08275_));
 sg13g2_buf_1 _14155_ (.A(_08276_),
    .X(_08277_));
 sg13g2_nand2_1 _14156_ (.Y(_08278_),
    .A(_08274_),
    .B(_08277_));
 sg13g2_buf_1 _14157_ (.A(\top_ihp.oisc.micro_pc[2] ),
    .X(_08279_));
 sg13g2_inv_1 _14158_ (.Y(_08280_),
    .A(_08279_));
 sg13g2_buf_1 _14159_ (.A(_08275_),
    .X(_08281_));
 sg13g2_nand2_1 _14160_ (.Y(_08282_),
    .A(_08280_),
    .B(net1008));
 sg13g2_buf_1 _14161_ (.A(_08282_),
    .X(_08283_));
 sg13g2_o21ai_1 _14162_ (.B1(net936),
    .Y(_08284_),
    .A1(_08273_),
    .A2(_08278_));
 sg13g2_inv_1 _14163_ (.Y(_08285_),
    .A(net1021));
 sg13g2_buf_1 _14164_ (.A(_08285_),
    .X(_08286_));
 sg13g2_nor2_1 _14165_ (.A(net973),
    .B(net936),
    .Y(_08287_));
 sg13g2_a21oi_1 _14166_ (.A1(net902),
    .A2(_08284_),
    .Y(_08288_),
    .B1(_08287_));
 sg13g2_nor3_1 _14167_ (.A(net1011),
    .B(_08263_),
    .C(_08288_),
    .Y(_08289_));
 sg13g2_buf_1 _14168_ (.A(net1010),
    .X(_08290_));
 sg13g2_buf_1 _14169_ (.A(_08280_),
    .X(_08291_));
 sg13g2_nor2_1 _14170_ (.A(net972),
    .B(net971),
    .Y(_08292_));
 sg13g2_buf_2 _14171_ (.A(\top_ihp.oisc.micro_pc[3] ),
    .X(_08293_));
 sg13g2_inv_1 _14172_ (.Y(_08294_),
    .A(_08293_));
 sg13g2_buf_1 _14173_ (.A(_08294_),
    .X(_08295_));
 sg13g2_nor2_1 _14174_ (.A(_08276_),
    .B(net970),
    .Y(_08296_));
 sg13g2_buf_2 _14175_ (.A(_08296_),
    .X(_08297_));
 sg13g2_inv_1 _14176_ (.Y(_08298_),
    .A(net1020));
 sg13g2_buf_1 _14177_ (.A(_08298_),
    .X(_08299_));
 sg13g2_buf_1 _14178_ (.A(net974),
    .X(_08300_));
 sg13g2_nand2_1 _14179_ (.Y(_08301_),
    .A(net969),
    .B(net935));
 sg13g2_buf_1 _14180_ (.A(_08279_),
    .X(_08302_));
 sg13g2_nor2_1 _14181_ (.A(net1007),
    .B(_08276_),
    .Y(_08303_));
 sg13g2_buf_1 _14182_ (.A(_08303_),
    .X(_08304_));
 sg13g2_buf_1 _14183_ (.A(_08274_),
    .X(_08305_));
 sg13g2_buf_1 _14184_ (.A(net1008),
    .X(_08306_));
 sg13g2_nor2_2 _14185_ (.A(_08305_),
    .B(net968),
    .Y(_08307_));
 sg13g2_inv_1 _14186_ (.Y(_08308_),
    .A(_08264_));
 sg13g2_buf_1 _14187_ (.A(_08308_),
    .X(_08309_));
 sg13g2_buf_1 _14188_ (.A(net967),
    .X(_08310_));
 sg13g2_o21ai_1 _14189_ (.B1(_08310_),
    .Y(_08311_),
    .A1(net934),
    .A2(_08307_));
 sg13g2_o21ai_1 _14190_ (.B1(_08311_),
    .Y(_08312_),
    .A1(net901),
    .A2(_08301_));
 sg13g2_buf_1 _14191_ (.A(_08295_),
    .X(_08313_));
 sg13g2_buf_1 _14192_ (.A(net932),
    .X(_08314_));
 sg13g2_buf_1 _14193_ (.A(\top_ihp.oisc.micro_pc[5] ),
    .X(_08315_));
 sg13g2_buf_1 _14194_ (.A(_08315_),
    .X(_08316_));
 sg13g2_buf_1 _14195_ (.A(_08316_),
    .X(_08317_));
 sg13g2_buf_1 _14196_ (.A(net966),
    .X(_08318_));
 sg13g2_a221oi_1 _14197_ (.B2(net900),
    .C1(net931),
    .B1(_08312_),
    .A1(_08292_),
    .Y(_08319_),
    .A2(_08297_));
 sg13g2_buf_1 _14198_ (.A(net935),
    .X(_08320_));
 sg13g2_buf_1 _14199_ (.A(net971),
    .X(_08321_));
 sg13g2_buf_1 _14200_ (.A(net972),
    .X(_08322_));
 sg13g2_nor2_1 _14201_ (.A(net1009),
    .B(_08313_),
    .Y(_08323_));
 sg13g2_buf_1 _14202_ (.A(_08293_),
    .X(_08324_));
 sg13g2_nor2_2 _14203_ (.A(_08286_),
    .B(net1004),
    .Y(_08325_));
 sg13g2_nor2_1 _14204_ (.A(_08323_),
    .B(_08325_),
    .Y(_08326_));
 sg13g2_buf_1 _14205_ (.A(net1004),
    .X(_08327_));
 sg13g2_nand2_1 _14206_ (.Y(_08328_),
    .A(_08286_),
    .B(net965));
 sg13g2_nor2_1 _14207_ (.A(net976),
    .B(_08328_),
    .Y(_08329_));
 sg13g2_a21oi_1 _14208_ (.A1(_08322_),
    .A2(_08326_),
    .Y(_08330_),
    .B1(_08329_));
 sg13g2_nor2_1 _14209_ (.A(net1007),
    .B(net970),
    .Y(_08331_));
 sg13g2_buf_1 _14210_ (.A(_08331_),
    .X(_08332_));
 sg13g2_nor2_1 _14211_ (.A(_08264_),
    .B(net973),
    .Y(_08333_));
 sg13g2_buf_1 _14212_ (.A(_08333_),
    .X(_08334_));
 sg13g2_nand2_1 _14213_ (.Y(_08335_),
    .A(net898),
    .B(net897));
 sg13g2_o21ai_1 _14214_ (.B1(_08335_),
    .Y(_08336_),
    .A1(net930),
    .A2(_08330_));
 sg13g2_nor2_1 _14215_ (.A(net967),
    .B(net1021),
    .Y(_08337_));
 sg13g2_buf_2 _14216_ (.A(_08337_),
    .X(_08338_));
 sg13g2_nand2_1 _14217_ (.Y(_08339_),
    .A(net1007),
    .B(net1008));
 sg13g2_buf_2 _14218_ (.A(_08339_),
    .X(_08340_));
 sg13g2_nor2_1 _14219_ (.A(net1011),
    .B(_08340_),
    .Y(_08341_));
 sg13g2_inv_2 _14220_ (.Y(_08342_),
    .A(_08315_));
 sg13g2_buf_1 _14221_ (.A(_08342_),
    .X(_08343_));
 sg13g2_buf_1 _14222_ (.A(_08343_),
    .X(_08344_));
 sg13g2_a221oi_1 _14223_ (.B2(_08341_),
    .C1(net928),
    .B1(_08338_),
    .A1(net899),
    .Y(_08345_),
    .A2(_08336_));
 sg13g2_nor3_1 _14224_ (.A(net977),
    .B(_08319_),
    .C(_08345_),
    .Y(_08346_));
 sg13g2_a21oi_1 _14225_ (.A1(_08260_),
    .A2(_08289_),
    .Y(_08347_),
    .B1(_08346_));
 sg13g2_buf_1 _14226_ (.A(net968),
    .X(_08348_));
 sg13g2_nor2_1 _14227_ (.A(_08264_),
    .B(net1021),
    .Y(_08349_));
 sg13g2_buf_1 _14228_ (.A(_08349_),
    .X(_08350_));
 sg13g2_nor2_1 _14229_ (.A(_08280_),
    .B(_08293_),
    .Y(_08351_));
 sg13g2_buf_2 _14230_ (.A(_08351_),
    .X(_08352_));
 sg13g2_nand2_1 _14231_ (.Y(_08353_),
    .A(net963),
    .B(_08352_));
 sg13g2_nand2_1 _14232_ (.Y(_08354_),
    .A(net972),
    .B(_08331_));
 sg13g2_nand3_1 _14233_ (.B(_08353_),
    .C(_08354_),
    .A(net927),
    .Y(_08355_));
 sg13g2_nand2_1 _14234_ (.Y(_08356_),
    .A(net967),
    .B(net1021));
 sg13g2_buf_2 _14235_ (.A(_08356_),
    .X(_08357_));
 sg13g2_nor3_2 _14236_ (.A(net1006),
    .B(net964),
    .C(_08357_),
    .Y(_08358_));
 sg13g2_inv_1 _14237_ (.Y(_08359_),
    .A(net1022));
 sg13g2_a22oi_1 _14238_ (.Y(_08360_),
    .B1(_08358_),
    .B2(_08359_),
    .A2(_08355_),
    .A1(_08344_));
 sg13g2_nor3_1 _14239_ (.A(net1006),
    .B(net1005),
    .C(_08357_),
    .Y(_08361_));
 sg13g2_nand2_1 _14240_ (.Y(_08362_),
    .A(net1010),
    .B(net1009));
 sg13g2_buf_1 _14241_ (.A(_08362_),
    .X(_08363_));
 sg13g2_buf_1 _14242_ (.A(_08363_),
    .X(_08364_));
 sg13g2_nor2_1 _14243_ (.A(_08278_),
    .B(net896),
    .Y(_08365_));
 sg13g2_buf_1 _14244_ (.A(net1023),
    .X(_08366_));
 sg13g2_a221oi_1 _14245_ (.B2(net931),
    .C1(net1003),
    .B1(_08365_),
    .A1(_08355_),
    .Y(_08367_),
    .A2(_08361_));
 sg13g2_o21ai_1 _14246_ (.B1(_08367_),
    .Y(_08368_),
    .A1(net899),
    .A2(_08360_));
 sg13g2_buf_1 _14247_ (.A(_08350_),
    .X(_08369_));
 sg13g2_nor2_1 _14248_ (.A(net1007),
    .B(_08275_),
    .Y(_08370_));
 sg13g2_buf_2 _14249_ (.A(_08370_),
    .X(_08371_));
 sg13g2_buf_1 _14250_ (.A(net1007),
    .X(_08372_));
 sg13g2_nand2_2 _14251_ (.Y(_08373_),
    .A(net962),
    .B(net974));
 sg13g2_o21ai_1 _14252_ (.B1(net936),
    .Y(_08374_),
    .A1(_08273_),
    .A2(_08373_));
 sg13g2_a22oi_1 _14253_ (.Y(_08375_),
    .B1(_08374_),
    .B2(net902),
    .A2(_08371_),
    .A1(net926));
 sg13g2_and2_1 _14254_ (.A(_08264_),
    .B(net1021),
    .X(_08376_));
 sg13g2_buf_1 _14255_ (.A(_08376_),
    .X(_08377_));
 sg13g2_nor2_2 _14256_ (.A(_08298_),
    .B(net1004),
    .Y(_08378_));
 sg13g2_nand2_1 _14257_ (.Y(_08379_),
    .A(_08263_),
    .B(net1023));
 sg13g2_a21oi_1 _14258_ (.A1(net961),
    .A2(_08378_),
    .Y(_08380_),
    .B1(_08379_));
 sg13g2_o21ai_1 _14259_ (.B1(_08380_),
    .Y(_08381_),
    .A1(_08314_),
    .A2(_08375_));
 sg13g2_a21oi_1 _14260_ (.A1(_08368_),
    .A2(_08381_),
    .Y(_08382_),
    .B1(net978));
 sg13g2_a21oi_1 _14261_ (.A1(net978),
    .A2(_08347_),
    .Y(_08383_),
    .B1(_08382_));
 sg13g2_buf_1 _14262_ (.A(_08253_),
    .X(_08384_));
 sg13g2_nand2_1 _14263_ (.Y(_08385_),
    .A(_07425_),
    .B(net843));
 sg13g2_o21ai_1 _14264_ (.B1(_08385_),
    .Y(_00269_),
    .A1(net844),
    .A2(_08383_));
 sg13g2_buf_1 _14265_ (.A(net927),
    .X(_08386_));
 sg13g2_nor2_1 _14266_ (.A(net973),
    .B(net1020),
    .Y(_08387_));
 sg13g2_nor3_1 _14267_ (.A(net1009),
    .B(_08302_),
    .C(net1008),
    .Y(_08388_));
 sg13g2_a21o_1 _14268_ (.A2(_08387_),
    .A1(net895),
    .B1(_08388_),
    .X(_08389_));
 sg13g2_buf_1 _14269_ (.A(net965),
    .X(_08390_));
 sg13g2_buf_1 _14270_ (.A(net925),
    .X(_08391_));
 sg13g2_a22oi_1 _14271_ (.Y(_08392_),
    .B1(_08389_),
    .B2(net894),
    .A2(_08325_),
    .A1(_08304_));
 sg13g2_nor2_1 _14272_ (.A(_08275_),
    .B(_08293_),
    .Y(_08393_));
 sg13g2_buf_1 _14273_ (.A(_08393_),
    .X(_08394_));
 sg13g2_nand2_2 _14274_ (.Y(_08395_),
    .A(net1021),
    .B(net1007));
 sg13g2_inv_1 _14275_ (.Y(_08396_),
    .A(_08395_));
 sg13g2_nor2_1 _14276_ (.A(net973),
    .B(_08279_),
    .Y(_08397_));
 sg13g2_buf_2 _14277_ (.A(_08397_),
    .X(_08398_));
 sg13g2_a22oi_1 _14278_ (.Y(_08399_),
    .B1(_08398_),
    .B2(_08290_),
    .A2(net963),
    .A1(net962));
 sg13g2_nor2_2 _14279_ (.A(net1008),
    .B(net970),
    .Y(_08400_));
 sg13g2_nor2_1 _14280_ (.A(net974),
    .B(net1004),
    .Y(_08401_));
 sg13g2_buf_1 _14281_ (.A(_08401_),
    .X(_08402_));
 sg13g2_nor2_1 _14282_ (.A(_08400_),
    .B(_08402_),
    .Y(_08403_));
 sg13g2_nand3b_1 _14283_ (.B(_08403_),
    .C(net1005),
    .Y(_08404_),
    .A_N(_08399_));
 sg13g2_nor2_2 _14284_ (.A(_08277_),
    .B(_08342_),
    .Y(_08405_));
 sg13g2_nor2_1 _14285_ (.A(net1020),
    .B(_08293_),
    .Y(_08406_));
 sg13g2_buf_1 _14286_ (.A(_08406_),
    .X(_08407_));
 sg13g2_nand3_1 _14287_ (.B(_08405_),
    .C(_08407_),
    .A(net961),
    .Y(_08408_));
 sg13g2_nand3_1 _14288_ (.B(_08404_),
    .C(_08408_),
    .A(net1023),
    .Y(_08409_));
 sg13g2_a21oi_1 _14289_ (.A1(net960),
    .A2(_08396_),
    .Y(_08410_),
    .B1(_08409_));
 sg13g2_o21ai_1 _14290_ (.B1(_08410_),
    .Y(_08411_),
    .A1(net902),
    .A2(_08392_));
 sg13g2_inv_1 _14291_ (.Y(_08412_),
    .A(_08409_));
 sg13g2_nand2_1 _14292_ (.Y(_08413_),
    .A(net974),
    .B(net1004));
 sg13g2_buf_1 _14293_ (.A(_08413_),
    .X(_08414_));
 sg13g2_nor2_1 _14294_ (.A(net1022),
    .B(net935),
    .Y(_08415_));
 sg13g2_nor3_1 _14295_ (.A(net933),
    .B(net960),
    .C(_08415_),
    .Y(_08416_));
 sg13g2_a21oi_1 _14296_ (.A1(net933),
    .A2(_08414_),
    .Y(_08417_),
    .B1(_08416_));
 sg13g2_buf_1 _14297_ (.A(_00088_),
    .X(_08418_));
 sg13g2_nor2b_1 _14298_ (.A(net894),
    .B_N(_08418_),
    .Y(_08419_));
 sg13g2_nor2_1 _14299_ (.A(net971),
    .B(net968),
    .Y(_08420_));
 sg13g2_a221oi_1 _14300_ (.B2(_08420_),
    .C1(net1003),
    .B1(_08419_),
    .A1(_08398_),
    .Y(_08421_),
    .A2(_08417_));
 sg13g2_buf_1 _14301_ (.A(net1005),
    .X(_08422_));
 sg13g2_buf_1 _14302_ (.A(net959),
    .X(_08423_));
 sg13g2_o21ai_1 _14303_ (.B1(net924),
    .Y(_08424_),
    .A1(_08412_),
    .A2(_08421_));
 sg13g2_a221oi_1 _14304_ (.B2(_08407_),
    .C1(net899),
    .B1(net926),
    .A1(net894),
    .Y(_08425_),
    .A2(_08418_));
 sg13g2_buf_1 _14305_ (.A(net895),
    .X(_08426_));
 sg13g2_buf_1 _14306_ (.A(net975),
    .X(_08427_));
 sg13g2_nand2_1 _14307_ (.Y(_08428_),
    .A(net923),
    .B(_08407_));
 sg13g2_buf_1 _14308_ (.A(net933),
    .X(_08429_));
 sg13g2_a21oi_1 _14309_ (.A1(_08328_),
    .A2(_08428_),
    .Y(_08430_),
    .B1(net893));
 sg13g2_nor2_1 _14310_ (.A(net876),
    .B(_08430_),
    .Y(_08431_));
 sg13g2_nor2_1 _14311_ (.A(_08316_),
    .B(net1023),
    .Y(_08432_));
 sg13g2_o21ai_1 _14312_ (.B1(_08432_),
    .Y(_08433_),
    .A1(_08425_),
    .A2(_08431_));
 sg13g2_nand3_1 _14313_ (.B(_08424_),
    .C(_08433_),
    .A(_08411_),
    .Y(_08434_));
 sg13g2_buf_1 _14314_ (.A(_08258_),
    .X(_08435_));
 sg13g2_buf_1 _14315_ (.A(net895),
    .X(_08436_));
 sg13g2_nand3_1 _14316_ (.B(_08359_),
    .C(net897),
    .A(net969),
    .Y(_08437_));
 sg13g2_nor2_1 _14317_ (.A(net1007),
    .B(net1004),
    .Y(_08438_));
 sg13g2_buf_1 _14318_ (.A(_08438_),
    .X(_08439_));
 sg13g2_nand3_1 _14319_ (.B(net961),
    .C(_08439_),
    .A(net966),
    .Y(_08440_));
 sg13g2_o21ai_1 _14320_ (.B1(_08440_),
    .Y(_08441_),
    .A1(net966),
    .A2(_08437_));
 sg13g2_buf_1 _14321_ (.A(_08348_),
    .X(_08442_));
 sg13g2_nor2_2 _14322_ (.A(net1021),
    .B(_08280_),
    .Y(_08443_));
 sg13g2_nor2_2 _14323_ (.A(_08443_),
    .B(_08398_),
    .Y(_08444_));
 sg13g2_nand2_1 _14324_ (.Y(_08445_),
    .A(_08265_),
    .B(net932));
 sg13g2_nand2_1 _14325_ (.Y(_08446_),
    .A(_08332_),
    .B(net963));
 sg13g2_o21ai_1 _14326_ (.B1(_08446_),
    .Y(_08447_),
    .A1(_08444_),
    .A2(_08445_));
 sg13g2_nand2_1 _14327_ (.Y(_08448_),
    .A(net966),
    .B(_08447_));
 sg13g2_buf_1 _14328_ (.A(net923),
    .X(_08449_));
 sg13g2_nor2_1 _14329_ (.A(_08372_),
    .B(net1005),
    .Y(_08450_));
 sg13g2_nand3_1 _14330_ (.B(net1011),
    .C(_08450_),
    .A(net891),
    .Y(_08451_));
 sg13g2_nand3_1 _14331_ (.B(_08448_),
    .C(_08451_),
    .A(net892),
    .Y(_08452_));
 sg13g2_o21ai_1 _14332_ (.B1(_08452_),
    .Y(_08453_),
    .A1(net875),
    .A2(_08441_));
 sg13g2_nand2_2 _14333_ (.Y(_08454_),
    .A(_08264_),
    .B(net973));
 sg13g2_nand2_1 _14334_ (.Y(_08455_),
    .A(_08270_),
    .B(net974));
 sg13g2_buf_2 _14335_ (.A(_08455_),
    .X(_08456_));
 sg13g2_o21ai_1 _14336_ (.B1(_08456_),
    .Y(_08457_),
    .A1(_08272_),
    .A2(_08283_));
 sg13g2_nand2_1 _14337_ (.Y(_08458_),
    .A(net893),
    .B(_08457_));
 sg13g2_o21ai_1 _14338_ (.B1(_08458_),
    .Y(_08459_),
    .A1(_08454_),
    .A2(_08278_));
 sg13g2_nand4_1 _14339_ (.B(_08263_),
    .C(net1003),
    .A(net1011),
    .Y(_08460_),
    .D(_08459_));
 sg13g2_o21ai_1 _14340_ (.B1(_08460_),
    .Y(_08461_),
    .A1(net1002),
    .A2(_08453_));
 sg13g2_nor2_1 _14341_ (.A(net978),
    .B(_08461_),
    .Y(_08462_));
 sg13g2_a21oi_1 _14342_ (.A1(net978),
    .A2(_08434_),
    .Y(_08463_),
    .B1(_08462_));
 sg13g2_mux2_1 _14343_ (.A0(_08463_),
    .A1(_08238_),
    .S(net843),
    .X(_00270_));
 sg13g2_buf_1 _14344_ (.A(_08255_),
    .X(_08464_));
 sg13g2_buf_1 _14345_ (.A(_08464_),
    .X(_08465_));
 sg13g2_buf_1 _14346_ (.A(net1003),
    .X(_08466_));
 sg13g2_nand2_1 _14347_ (.Y(_08467_),
    .A(_08291_),
    .B(_08327_));
 sg13g2_nand2_1 _14348_ (.Y(_08468_),
    .A(net1007),
    .B(_08293_));
 sg13g2_buf_2 _14349_ (.A(_08468_),
    .X(_08469_));
 sg13g2_o21ai_1 _14350_ (.B1(_08428_),
    .Y(_08470_),
    .A1(net891),
    .A2(_08469_));
 sg13g2_nand2_1 _14351_ (.Y(_08471_),
    .A(_08429_),
    .B(_08470_));
 sg13g2_o21ai_1 _14352_ (.B1(_08471_),
    .Y(_08472_),
    .A1(_08467_),
    .A2(net896));
 sg13g2_nor2_2 _14353_ (.A(_08281_),
    .B(_08342_),
    .Y(_08473_));
 sg13g2_nor3_1 _14354_ (.A(net1006),
    .B(net1022),
    .C(_08363_),
    .Y(_08474_));
 sg13g2_buf_1 _14355_ (.A(_00084_),
    .X(_08475_));
 sg13g2_nor2_1 _14356_ (.A(net1005),
    .B(_08475_),
    .Y(_08476_));
 sg13g2_a22oi_1 _14357_ (.Y(_08477_),
    .B1(_08474_),
    .B2(_08476_),
    .A2(_08473_),
    .A1(_08472_));
 sg13g2_inv_1 _14358_ (.Y(_08478_),
    .A(_08475_));
 sg13g2_nand4_1 _14359_ (.B(_08435_),
    .C(_08478_),
    .A(net1011),
    .Y(_08479_),
    .D(_08358_));
 sg13g2_o21ai_1 _14360_ (.B1(_08479_),
    .Y(_08480_),
    .A1(net957),
    .A2(_08477_));
 sg13g2_a22oi_1 _14361_ (.Y(_08481_),
    .B1(net961),
    .B2(net934),
    .A2(net926),
    .A1(_08307_));
 sg13g2_nor3_1 _14362_ (.A(_08262_),
    .B(_08318_),
    .C(_08481_),
    .Y(_08482_));
 sg13g2_nor2_1 _14363_ (.A(net1009),
    .B(_08298_),
    .Y(_08483_));
 sg13g2_nor3_1 _14364_ (.A(_08265_),
    .B(_08387_),
    .C(_08483_),
    .Y(_08484_));
 sg13g2_a21oi_1 _14365_ (.A1(net1006),
    .A2(_08338_),
    .Y(_08485_),
    .B1(_08484_));
 sg13g2_o21ai_1 _14366_ (.B1(_08405_),
    .Y(_08486_),
    .A1(_08262_),
    .A2(_08485_));
 sg13g2_nand2_1 _14367_ (.Y(_08487_),
    .A(_08280_),
    .B(net970));
 sg13g2_buf_1 _14368_ (.A(_08487_),
    .X(_08488_));
 sg13g2_o21ai_1 _14369_ (.B1(net935),
    .Y(_08489_),
    .A1(_08357_),
    .A2(_08488_));
 sg13g2_nand2_1 _14370_ (.Y(_08490_),
    .A(net966),
    .B(_08489_));
 sg13g2_nor2_2 _14371_ (.A(net1020),
    .B(net970),
    .Y(_08491_));
 sg13g2_nand4_1 _14372_ (.B(_08475_),
    .C(_08338_),
    .A(net928),
    .Y(_08492_),
    .D(_08491_));
 sg13g2_a21oi_1 _14373_ (.A1(_08490_),
    .A2(_08492_),
    .Y(_08493_),
    .B1(net1002));
 sg13g2_a22oi_1 _14374_ (.Y(_08494_),
    .B1(_08486_),
    .B2(_08493_),
    .A2(_08482_),
    .A1(net957));
 sg13g2_nand2_1 _14375_ (.Y(_08495_),
    .A(net958),
    .B(_08494_));
 sg13g2_o21ai_1 _14376_ (.B1(_08495_),
    .Y(_08496_),
    .A1(net958),
    .A2(_08480_));
 sg13g2_nand2_1 _14377_ (.Y(_08497_),
    .A(\top_ihp.oisc.micro_op[11] ),
    .B(net843));
 sg13g2_o21ai_1 _14378_ (.B1(_08497_),
    .Y(_00271_),
    .A1(net844),
    .A2(_08496_));
 sg13g2_a21oi_1 _14379_ (.A1(_08357_),
    .A2(_08454_),
    .Y(_08498_),
    .B1(_08299_));
 sg13g2_nor2_1 _14380_ (.A(net923),
    .B(_08488_),
    .Y(_08499_));
 sg13g2_a21oi_1 _14381_ (.A1(_08390_),
    .A2(_08498_),
    .Y(_08500_),
    .B1(_08499_));
 sg13g2_nand2_1 _14382_ (.Y(_08501_),
    .A(net965),
    .B(_08418_));
 sg13g2_nor2_1 _14383_ (.A(net930),
    .B(_08501_),
    .Y(_08502_));
 sg13g2_nand2_1 _14384_ (.Y(_08503_),
    .A(_08298_),
    .B(net970));
 sg13g2_buf_1 _14385_ (.A(_08503_),
    .X(_08504_));
 sg13g2_nand2_1 _14386_ (.Y(_08505_),
    .A(net967),
    .B(net973));
 sg13g2_buf_1 _14387_ (.A(_08505_),
    .X(_08506_));
 sg13g2_a21oi_1 _14388_ (.A1(_08467_),
    .A2(_08504_),
    .Y(_08507_),
    .B1(_08506_));
 sg13g2_nor3_1 _14389_ (.A(_08386_),
    .B(_08502_),
    .C(_08507_),
    .Y(_08508_));
 sg13g2_a21oi_1 _14390_ (.A1(net876),
    .A2(_08500_),
    .Y(_08509_),
    .B1(_08508_));
 sg13g2_buf_1 _14391_ (.A(net973),
    .X(_08510_));
 sg13g2_nor2_2 _14392_ (.A(net1022),
    .B(net1008),
    .Y(_08511_));
 sg13g2_nor2_1 _14393_ (.A(net967),
    .B(net1006),
    .Y(_08512_));
 sg13g2_a22oi_1 _14394_ (.Y(_08513_),
    .B1(_08511_),
    .B2(_08512_),
    .A2(net934),
    .A1(net1022));
 sg13g2_nor2_1 _14395_ (.A(net971),
    .B(net935),
    .Y(_08514_));
 sg13g2_nand3_1 _14396_ (.B(net1022),
    .C(_08514_),
    .A(net933),
    .Y(_08515_));
 sg13g2_o21ai_1 _14397_ (.B1(_08515_),
    .Y(_08516_),
    .A1(_08510_),
    .A2(_08513_));
 sg13g2_and2_1 _14398_ (.A(_08344_),
    .B(_08516_),
    .X(_08517_));
 sg13g2_a21oi_1 _14399_ (.A1(net924),
    .A2(_08509_),
    .Y(_08518_),
    .B1(_08517_));
 sg13g2_nand2_1 _14400_ (.Y(_08519_),
    .A(net965),
    .B(_08371_));
 sg13g2_nor3_1 _14401_ (.A(net971),
    .B(net974),
    .C(net932),
    .Y(_08520_));
 sg13g2_nor3_1 _14402_ (.A(net976),
    .B(_08352_),
    .C(_08371_),
    .Y(_08521_));
 sg13g2_buf_1 _14403_ (.A(net891),
    .X(_08522_));
 sg13g2_o21ai_1 _14404_ (.B1(net874),
    .Y(_08523_),
    .A1(_08520_),
    .A2(_08521_));
 sg13g2_o21ai_1 _14405_ (.B1(_08523_),
    .Y(_08524_),
    .A1(net890),
    .A2(_08519_));
 sg13g2_a21oi_1 _14406_ (.A1(_08263_),
    .A2(_08524_),
    .Y(_08525_),
    .B1(net977));
 sg13g2_a21oi_1 _14407_ (.A1(net977),
    .A2(_08518_),
    .Y(_08526_),
    .B1(_08525_));
 sg13g2_nand2_1 _14408_ (.Y(_08527_),
    .A(net1020),
    .B(net970));
 sg13g2_o21ai_1 _14409_ (.B1(_08527_),
    .Y(_08528_),
    .A1(net976),
    .A2(_08469_));
 sg13g2_buf_1 _14410_ (.A(_00087_),
    .X(_08529_));
 sg13g2_nand2_1 _14411_ (.Y(_08530_),
    .A(net932),
    .B(_08529_));
 sg13g2_nand3_1 _14412_ (.B(_08354_),
    .C(_08530_),
    .A(net937),
    .Y(_08531_));
 sg13g2_o21ai_1 _14413_ (.B1(_08531_),
    .Y(_08532_),
    .A1(net891),
    .A2(_08528_));
 sg13g2_nand2_2 _14414_ (.Y(_08533_),
    .A(_08302_),
    .B(net970));
 sg13g2_nand2_1 _14415_ (.Y(_08534_),
    .A(net1009),
    .B(_08491_));
 sg13g2_a21oi_1 _14416_ (.A1(_08533_),
    .A2(_08534_),
    .Y(_08535_),
    .B1(net929));
 sg13g2_nor3_1 _14417_ (.A(net927),
    .B(_08499_),
    .C(_08535_),
    .Y(_08536_));
 sg13g2_a21o_1 _14418_ (.A2(_08532_),
    .A1(net892),
    .B1(_08536_),
    .X(_08537_));
 sg13g2_buf_1 _14419_ (.A(net1020),
    .X(_08538_));
 sg13g2_nor2_1 _14420_ (.A(_08309_),
    .B(_08313_),
    .Y(_08539_));
 sg13g2_a21oi_1 _14421_ (.A1(net1000),
    .A2(_08539_),
    .Y(_08540_),
    .B1(_08439_));
 sg13g2_nand2_1 _14422_ (.Y(_08541_),
    .A(net1008),
    .B(net932));
 sg13g2_buf_1 _14423_ (.A(_08541_),
    .X(_08542_));
 sg13g2_nand2_1 _14424_ (.Y(_08543_),
    .A(_08414_),
    .B(_08542_));
 sg13g2_nor2_1 _14425_ (.A(net897),
    .B(_08543_),
    .Y(_08544_));
 sg13g2_o21ai_1 _14426_ (.B1(_08544_),
    .Y(_08545_),
    .A1(net874),
    .A2(_08540_));
 sg13g2_a21oi_1 _14427_ (.A1(net937),
    .A2(_08504_),
    .Y(_08546_),
    .B1(net898));
 sg13g2_nor2_1 _14428_ (.A(net929),
    .B(_08483_),
    .Y(_08547_));
 sg13g2_a22oi_1 _14429_ (.Y(_08548_),
    .B1(_08547_),
    .B2(_08428_),
    .A2(_08546_),
    .A1(net938));
 sg13g2_nand2_1 _14430_ (.Y(_08549_),
    .A(_08398_),
    .B(net960));
 sg13g2_o21ai_1 _14431_ (.B1(net922),
    .Y(_08550_),
    .A1(net925),
    .A2(_08307_));
 sg13g2_buf_1 _14432_ (.A(net929),
    .X(_08551_));
 sg13g2_a21oi_1 _14433_ (.A1(_08549_),
    .A2(_08550_),
    .Y(_08552_),
    .B1(net889));
 sg13g2_a21oi_1 _14434_ (.A1(net892),
    .A2(_08548_),
    .Y(_08553_),
    .B1(_08552_));
 sg13g2_nand2_1 _14435_ (.Y(_08554_),
    .A(net976),
    .B(_08371_));
 sg13g2_nor2_1 _14436_ (.A(net1010),
    .B(net932),
    .Y(_08555_));
 sg13g2_o21ai_1 _14437_ (.B1(_08555_),
    .Y(_08556_),
    .A1(_08304_),
    .A2(_08420_));
 sg13g2_o21ai_1 _14438_ (.B1(_08556_),
    .Y(_08557_),
    .A1(net969),
    .A2(_08554_));
 sg13g2_nor2_1 _14439_ (.A(net967),
    .B(net971),
    .Y(_08558_));
 sg13g2_nand2_1 _14440_ (.Y(_08559_),
    .A(net1010),
    .B(_08281_));
 sg13g2_o21ai_1 _14441_ (.B1(_08559_),
    .Y(_08560_),
    .A1(net972),
    .A2(_08278_));
 sg13g2_a22oi_1 _14442_ (.Y(_08561_),
    .B1(_08560_),
    .B2(_08272_),
    .A2(_08558_),
    .A1(_08301_));
 sg13g2_a221oi_1 _14443_ (.B2(net933),
    .C1(net925),
    .B1(_08396_),
    .A1(net930),
    .Y(_08562_),
    .A2(_08338_));
 sg13g2_a21oi_1 _14444_ (.A1(net925),
    .A2(_08561_),
    .Y(_08563_),
    .B1(_08562_));
 sg13g2_a221oi_1 _14445_ (.B2(net922),
    .C1(_08563_),
    .B1(_08557_),
    .A1(net961),
    .Y(_08564_),
    .A2(_08420_));
 sg13g2_mux4_1 _14446_ (.S0(net1003),
    .A0(_08537_),
    .A1(_08545_),
    .A2(_08553_),
    .A3(_08564_),
    .S1(net928),
    .X(_08565_));
 sg13g2_nand2_1 _14447_ (.Y(_08566_),
    .A(net978),
    .B(_08565_));
 sg13g2_o21ai_1 _14448_ (.B1(_08566_),
    .Y(_08567_),
    .A1(net978),
    .A2(_08526_));
 sg13g2_nand2_1 _14449_ (.Y(_08568_),
    .A(\top_ihp.oisc.micro_op[12] ),
    .B(net843));
 sg13g2_o21ai_1 _14450_ (.B1(_08568_),
    .Y(_00272_),
    .A1(net844),
    .A2(_08567_));
 sg13g2_buf_1 _14451_ (.A(net962),
    .X(_08569_));
 sg13g2_nor2_1 _14452_ (.A(net921),
    .B(_08357_),
    .Y(_08570_));
 sg13g2_and2_1 _14453_ (.A(_08543_),
    .B(_08570_),
    .X(_08571_));
 sg13g2_a21o_1 _14454_ (.A2(_08544_),
    .A1(net969),
    .B1(_08571_),
    .X(_08572_));
 sg13g2_nor2_1 _14455_ (.A(net968),
    .B(_08378_),
    .Y(_08573_));
 sg13g2_nor3_1 _14456_ (.A(net933),
    .B(net898),
    .C(_08573_),
    .Y(_08574_));
 sg13g2_nor3_1 _14457_ (.A(net901),
    .B(_08521_),
    .C(_08574_),
    .Y(_08575_));
 sg13g2_o21ai_1 _14458_ (.B1(_08519_),
    .Y(_08576_),
    .A1(net930),
    .A2(_08542_));
 sg13g2_a21oi_1 _14459_ (.A1(net894),
    .A2(_08340_),
    .Y(_08577_),
    .B1(net896));
 sg13g2_nor4_1 _14460_ (.A(net959),
    .B(_08575_),
    .C(_08576_),
    .D(_08577_),
    .Y(_08578_));
 sg13g2_a21oi_1 _14461_ (.A1(net924),
    .A2(_08572_),
    .Y(_08579_),
    .B1(_08578_));
 sg13g2_nand2_1 _14462_ (.Y(_08580_),
    .A(net1009),
    .B(net1004));
 sg13g2_o21ai_1 _14463_ (.B1(_08580_),
    .Y(_08581_),
    .A1(net923),
    .A2(_08504_));
 sg13g2_nand2_1 _14464_ (.Y(_08582_),
    .A(net938),
    .B(_08581_));
 sg13g2_o21ai_1 _14465_ (.B1(net893),
    .Y(_08583_),
    .A1(_08323_),
    .A2(_08398_));
 sg13g2_nand3_1 _14466_ (.B(_08582_),
    .C(_08583_),
    .A(_08426_),
    .Y(_08584_));
 sg13g2_nor2_1 _14467_ (.A(net1022),
    .B(net921),
    .Y(_08585_));
 sg13g2_nand2_1 _14468_ (.Y(_08586_),
    .A(net897),
    .B(_08585_));
 sg13g2_nand2_1 _14469_ (.Y(_08587_),
    .A(net899),
    .B(_08586_));
 sg13g2_nand4_1 _14470_ (.B(net1001),
    .C(_08584_),
    .A(_08263_),
    .Y(_08588_),
    .D(_08587_));
 sg13g2_o21ai_1 _14471_ (.B1(_08588_),
    .Y(_08589_),
    .A1(net1001),
    .A2(_08579_));
 sg13g2_nor2_2 _14472_ (.A(net962),
    .B(_08454_),
    .Y(_08590_));
 sg13g2_a21oi_1 _14473_ (.A1(_08569_),
    .A2(_08418_),
    .Y(_08591_),
    .B1(_08590_));
 sg13g2_nand2b_1 _14474_ (.Y(_08592_),
    .B(net967),
    .A_N(_08580_));
 sg13g2_o21ai_1 _14475_ (.B1(_08592_),
    .Y(_08593_),
    .A1(_08390_),
    .A2(_08591_));
 sg13g2_o21ai_1 _14476_ (.B1(net935),
    .Y(_08594_),
    .A1(_08261_),
    .A2(net961));
 sg13g2_o21ai_1 _14477_ (.B1(_08594_),
    .Y(_08595_),
    .A1(net899),
    .A2(_08593_));
 sg13g2_a21oi_1 _14478_ (.A1(_08427_),
    .A2(_08402_),
    .Y(_08596_),
    .B1(_08323_));
 sg13g2_nand2_1 _14479_ (.Y(_08597_),
    .A(net897),
    .B(net960));
 sg13g2_o21ai_1 _14480_ (.B1(_08597_),
    .Y(_08598_),
    .A1(net933),
    .A2(_08596_));
 sg13g2_nand2_1 _14481_ (.Y(_08599_),
    .A(_08530_),
    .B(_08592_));
 sg13g2_a221oi_1 _14482_ (.B2(_08514_),
    .C1(net959),
    .B1(_08599_),
    .A1(net930),
    .Y(_08600_),
    .A2(_08598_));
 sg13g2_a21oi_1 _14483_ (.A1(_08318_),
    .A2(_08595_),
    .Y(_08601_),
    .B1(_08600_));
 sg13g2_nand2_2 _14484_ (.Y(_08602_),
    .A(_08324_),
    .B(_08342_));
 sg13g2_nor2_1 _14485_ (.A(net930),
    .B(_08602_),
    .Y(_08603_));
 sg13g2_o21ai_1 _14486_ (.B1(net902),
    .Y(_08604_),
    .A1(_08398_),
    .A2(_08603_));
 sg13g2_buf_1 _14487_ (.A(_08569_),
    .X(_08605_));
 sg13g2_nor3_1 _14488_ (.A(_08605_),
    .B(net890),
    .C(_08602_),
    .Y(_08606_));
 sg13g2_nor2_1 _14489_ (.A(_08473_),
    .B(_08606_),
    .Y(_08607_));
 sg13g2_nor2_1 _14490_ (.A(net925),
    .B(net964),
    .Y(_08608_));
 sg13g2_o21ai_1 _14491_ (.B1(net874),
    .Y(_08609_),
    .A1(_08603_),
    .A2(_08608_));
 sg13g2_nand3_1 _14492_ (.B(_08607_),
    .C(_08609_),
    .A(_08604_),
    .Y(_08610_));
 sg13g2_nor2_1 _14493_ (.A(net923),
    .B(_08342_),
    .Y(_08611_));
 sg13g2_nand2_2 _14494_ (.Y(_08612_),
    .A(_08299_),
    .B(net965));
 sg13g2_o21ai_1 _14495_ (.B1(_08488_),
    .Y(_08613_),
    .A1(net938),
    .A2(_08612_));
 sg13g2_a21oi_1 _14496_ (.A1(_08611_),
    .A2(_08613_),
    .Y(_08614_),
    .B1(net876));
 sg13g2_nor2_1 _14497_ (.A(_08255_),
    .B(_08614_),
    .Y(_08615_));
 sg13g2_a22oi_1 _14498_ (.Y(_08616_),
    .B1(_08610_),
    .B2(_08615_),
    .A2(_08601_),
    .A1(net1001));
 sg13g2_nor2_1 _14499_ (.A(_08466_),
    .B(_08616_),
    .Y(_08617_));
 sg13g2_a21oi_1 _14500_ (.A1(net957),
    .A2(_08589_),
    .Y(_08618_),
    .B1(_08617_));
 sg13g2_nand2_1 _14501_ (.Y(_08619_),
    .A(\top_ihp.oisc.micro_op[13] ),
    .B(_08384_));
 sg13g2_o21ai_1 _14502_ (.B1(_08619_),
    .Y(_00273_),
    .A1(net844),
    .A2(_08618_));
 sg13g2_nand2_1 _14503_ (.Y(_08620_),
    .A(net1020),
    .B(_08400_));
 sg13g2_o21ai_1 _14504_ (.B1(_08620_),
    .Y(_08621_),
    .A1(net1000),
    .A2(_08542_));
 sg13g2_buf_1 _14505_ (.A(net972),
    .X(_08622_));
 sg13g2_a22oi_1 _14506_ (.Y(_08623_),
    .B1(net960),
    .B2(net921),
    .A2(_08297_),
    .A1(net969));
 sg13g2_nand2_1 _14507_ (.Y(_08624_),
    .A(net920),
    .B(_08623_));
 sg13g2_o21ai_1 _14508_ (.B1(_08624_),
    .Y(_08625_),
    .A1(net889),
    .A2(_08621_));
 sg13g2_a221oi_1 _14509_ (.B2(_08340_),
    .C1(net901),
    .B1(_08539_),
    .A1(_08292_),
    .Y(_08626_),
    .A2(_08394_));
 sg13g2_a21oi_1 _14510_ (.A1(net874),
    .A2(_08625_),
    .Y(_08627_),
    .B1(_08626_));
 sg13g2_nor3_1 _14511_ (.A(net972),
    .B(_08443_),
    .C(_08398_),
    .Y(_08628_));
 sg13g2_a21oi_1 _14512_ (.A1(_08322_),
    .A2(_08395_),
    .Y(_08629_),
    .B1(_08628_));
 sg13g2_a221oi_1 _14513_ (.B2(net900),
    .C1(net895),
    .B1(_08629_),
    .A1(net926),
    .Y(_08630_),
    .A2(_08491_));
 sg13g2_nor2_1 _14514_ (.A(net1010),
    .B(_08327_),
    .Y(_08631_));
 sg13g2_a21oi_1 _14515_ (.A1(_08266_),
    .A2(_08332_),
    .Y(_08632_),
    .B1(_08631_));
 sg13g2_nor2_1 _14516_ (.A(_08449_),
    .B(_08632_),
    .Y(_08633_));
 sg13g2_nor3_1 _14517_ (.A(_08320_),
    .B(_08502_),
    .C(_08633_),
    .Y(_08634_));
 sg13g2_nor3_1 _14518_ (.A(net1003),
    .B(_08630_),
    .C(_08634_),
    .Y(_08635_));
 sg13g2_a21oi_1 _14519_ (.A1(net1002),
    .A2(_08627_),
    .Y(_08636_),
    .B1(_08635_));
 sg13g2_nor2_2 _14520_ (.A(net975),
    .B(net962),
    .Y(_08637_));
 sg13g2_nor2_1 _14521_ (.A(net938),
    .B(_08637_),
    .Y(_08638_));
 sg13g2_a21oi_1 _14522_ (.A1(net874),
    .A2(_08352_),
    .Y(_08639_),
    .B1(_08638_));
 sg13g2_a21o_1 _14523_ (.A2(net934),
    .A1(net920),
    .B1(_08292_),
    .X(_08640_));
 sg13g2_nand3_1 _14524_ (.B(_08359_),
    .C(_08640_),
    .A(net922),
    .Y(_08641_));
 sg13g2_o21ai_1 _14525_ (.B1(_08641_),
    .Y(_08642_),
    .A1(net876),
    .A2(_08639_));
 sg13g2_nor2_1 _14526_ (.A(net928),
    .B(_08366_),
    .Y(_08643_));
 sg13g2_nand3_1 _14527_ (.B(net961),
    .C(_08373_),
    .A(net936),
    .Y(_08644_));
 sg13g2_o21ai_1 _14528_ (.B1(_08644_),
    .Y(_08645_),
    .A1(net936),
    .A2(net890));
 sg13g2_nand2_1 _14529_ (.Y(_08646_),
    .A(net1006),
    .B(net965));
 sg13g2_nor3_1 _14530_ (.A(net897),
    .B(_08338_),
    .C(_08646_),
    .Y(_08647_));
 sg13g2_a22oi_1 _14531_ (.Y(_08648_),
    .B1(_08647_),
    .B2(_08405_),
    .A2(_08645_),
    .A1(_08608_));
 sg13g2_nor2_1 _14532_ (.A(_08260_),
    .B(_08648_),
    .Y(_08649_));
 sg13g2_a21oi_1 _14533_ (.A1(_08642_),
    .A2(_08643_),
    .Y(_08650_),
    .B1(_08649_));
 sg13g2_o21ai_1 _14534_ (.B1(_08650_),
    .Y(_08651_),
    .A1(_08423_),
    .A2(_08636_));
 sg13g2_a22oi_1 _14535_ (.Y(_08652_),
    .B1(_08373_),
    .B2(_08378_),
    .A2(_08533_),
    .A1(_08307_));
 sg13g2_buf_1 _14536_ (.A(net962),
    .X(_08653_));
 sg13g2_nand2_1 _14537_ (.Y(_08654_),
    .A(net919),
    .B(net960));
 sg13g2_nand2_1 _14538_ (.Y(_08655_),
    .A(net971),
    .B(_08297_));
 sg13g2_o21ai_1 _14539_ (.B1(net1000),
    .Y(_08656_),
    .A1(net934),
    .A2(_08352_));
 sg13g2_nand3_1 _14540_ (.B(_08655_),
    .C(_08656_),
    .A(_08654_),
    .Y(_08657_));
 sg13g2_nand2_1 _14541_ (.Y(_08658_),
    .A(net926),
    .B(_08657_));
 sg13g2_o21ai_1 _14542_ (.B1(_08658_),
    .Y(_08659_),
    .A1(net896),
    .A2(_08652_));
 sg13g2_nor2_1 _14543_ (.A(net922),
    .B(_08488_),
    .Y(_08660_));
 sg13g2_nor2_1 _14544_ (.A(net891),
    .B(_08612_),
    .Y(_08661_));
 sg13g2_nor2_1 _14545_ (.A(_08267_),
    .B(_08300_),
    .Y(_08662_));
 sg13g2_o21ai_1 _14546_ (.B1(_08662_),
    .Y(_08663_),
    .A1(_08660_),
    .A2(_08661_));
 sg13g2_a21oi_1 _14547_ (.A1(_08445_),
    .A2(_08469_),
    .Y(_08664_),
    .B1(_08456_));
 sg13g2_nor2_1 _14548_ (.A(net1023),
    .B(_08664_),
    .Y(_08665_));
 sg13g2_nor2_1 _14549_ (.A(net975),
    .B(_08445_),
    .Y(_08666_));
 sg13g2_o21ai_1 _14550_ (.B1(net919),
    .Y(_08667_),
    .A1(_08555_),
    .A2(_08666_));
 sg13g2_o21ai_1 _14551_ (.B1(_08667_),
    .Y(_08668_),
    .A1(net888),
    .A2(_08530_));
 sg13g2_nand2_1 _14552_ (.Y(_08669_),
    .A(net895),
    .B(_08437_));
 sg13g2_o21ai_1 _14553_ (.B1(_08669_),
    .Y(_08670_),
    .A1(_08442_),
    .A2(_08668_));
 sg13g2_a22oi_1 _14554_ (.Y(_08671_),
    .B1(_08670_),
    .B2(net1002),
    .A2(_08665_),
    .A1(_08663_));
 sg13g2_a22oi_1 _14555_ (.Y(_08672_),
    .B1(_08671_),
    .B2(net928),
    .A2(_08659_),
    .A1(_08643_));
 sg13g2_nand2_1 _14556_ (.Y(_08673_),
    .A(net958),
    .B(_08672_));
 sg13g2_o21ai_1 _14557_ (.B1(_08673_),
    .Y(_08674_),
    .A1(net958),
    .A2(_08651_));
 sg13g2_nand2_1 _14558_ (.Y(_08675_),
    .A(\top_ihp.oisc.micro_op[14] ),
    .B(_08384_));
 sg13g2_o21ai_1 _14559_ (.B1(_08675_),
    .Y(_00274_),
    .A1(_08254_),
    .A2(_08674_));
 sg13g2_nor2_1 _14560_ (.A(net964),
    .B(_08539_),
    .Y(_08676_));
 sg13g2_nand2_1 _14561_ (.Y(_08677_),
    .A(net932),
    .B(net1005));
 sg13g2_o21ai_1 _14562_ (.B1(_08602_),
    .Y(_08678_),
    .A1(net927),
    .A2(_08677_));
 sg13g2_nand2_1 _14563_ (.Y(_08679_),
    .A(net926),
    .B(_08678_));
 sg13g2_o21ai_1 _14564_ (.B1(_08679_),
    .Y(_08680_),
    .A1(_08456_),
    .A2(_08676_));
 sg13g2_o21ai_1 _14565_ (.B1(_08646_),
    .Y(_08681_),
    .A1(net937),
    .A2(_08504_));
 sg13g2_a22oi_1 _14566_ (.Y(_08682_),
    .B1(_08681_),
    .B2(_08551_),
    .A2(_08439_),
    .A1(net963));
 sg13g2_nand2_2 _14567_ (.Y(_08683_),
    .A(net965),
    .B(net1005));
 sg13g2_inv_1 _14568_ (.Y(_08684_),
    .A(_08683_));
 sg13g2_a22oi_1 _14569_ (.Y(_08685_),
    .B1(_08684_),
    .B2(_08538_),
    .A2(_08450_),
    .A1(net929));
 sg13g2_nand2b_1 _14570_ (.Y(_08686_),
    .B(net901),
    .A_N(_08685_));
 sg13g2_o21ai_1 _14571_ (.B1(_08686_),
    .Y(_08687_),
    .A1(net928),
    .A2(_08682_));
 sg13g2_nand2_1 _14572_ (.Y(_08688_),
    .A(net923),
    .B(_08602_));
 sg13g2_a21oi_1 _14573_ (.A1(_08677_),
    .A2(_08688_),
    .Y(_08689_),
    .B1(_08554_));
 sg13g2_a221oi_1 _14574_ (.B2(net875),
    .C1(_08689_),
    .B1(_08687_),
    .A1(net888),
    .Y(_08690_),
    .A2(_08680_));
 sg13g2_o21ai_1 _14575_ (.B1(net919),
    .Y(_08691_),
    .A1(_08400_),
    .A2(_08415_));
 sg13g2_o21ai_1 _14576_ (.B1(_08691_),
    .Y(_08692_),
    .A1(net901),
    .A2(_08414_));
 sg13g2_nand2_1 _14577_ (.Y(_08693_),
    .A(net967),
    .B(net935));
 sg13g2_nand2_1 _14578_ (.Y(_08694_),
    .A(_08559_),
    .B(_08693_));
 sg13g2_a22oi_1 _14579_ (.Y(_08695_),
    .B1(_08694_),
    .B2(_08660_),
    .A2(_08692_),
    .A1(net893));
 sg13g2_or2_1 _14580_ (.X(_08696_),
    .B(_08695_),
    .A(_08379_));
 sg13g2_o21ai_1 _14581_ (.B1(_08696_),
    .Y(_08697_),
    .A1(net957),
    .A2(_08690_));
 sg13g2_nor2_1 _14582_ (.A(_08309_),
    .B(net962),
    .Y(_08698_));
 sg13g2_o21ai_1 _14583_ (.B1(net936),
    .Y(_08699_),
    .A1(_08291_),
    .A2(_08402_));
 sg13g2_a22oi_1 _14584_ (.Y(_08700_),
    .B1(_08699_),
    .B2(_08310_),
    .A2(_08698_),
    .A1(_08394_));
 sg13g2_o21ai_1 _14585_ (.B1(_08542_),
    .Y(_08701_),
    .A1(net922),
    .A2(_08414_));
 sg13g2_nand3_1 _14586_ (.B(net919),
    .C(_08701_),
    .A(net938),
    .Y(_08702_));
 sg13g2_o21ai_1 _14587_ (.B1(_08702_),
    .Y(_08703_),
    .A1(net901),
    .A2(_08700_));
 sg13g2_inv_1 _14588_ (.Y(_08704_),
    .A(_08703_));
 sg13g2_nand2_1 _14589_ (.Y(_08705_),
    .A(net937),
    .B(_08533_));
 sg13g2_nand2_1 _14590_ (.Y(_08706_),
    .A(net919),
    .B(net896));
 sg13g2_a22oi_1 _14591_ (.Y(_08707_),
    .B1(_08706_),
    .B2(_08491_),
    .A2(_08705_),
    .A1(net893));
 sg13g2_a22oi_1 _14592_ (.Y(_08708_),
    .B1(_08707_),
    .B2(net899),
    .A2(_08341_),
    .A1(net893));
 sg13g2_nor2_1 _14593_ (.A(net1000),
    .B(net896),
    .Y(_08709_));
 sg13g2_a22oi_1 _14594_ (.Y(_08710_),
    .B1(_08576_),
    .B2(net893),
    .A2(_08709_),
    .A1(_08297_));
 sg13g2_nor2_1 _14595_ (.A(net1009),
    .B(_08527_),
    .Y(_08711_));
 sg13g2_a21oi_1 _14596_ (.A1(net937),
    .A2(net925),
    .Y(_08712_),
    .B1(_08711_));
 sg13g2_nand2_1 _14597_ (.Y(_08713_),
    .A(net975),
    .B(_08378_));
 sg13g2_nor2_1 _14598_ (.A(net929),
    .B(_08443_),
    .Y(_08714_));
 sg13g2_a22oi_1 _14599_ (.Y(_08715_),
    .B1(_08713_),
    .B2(_08714_),
    .A2(_08712_),
    .A1(net938));
 sg13g2_o21ai_1 _14600_ (.B1(net969),
    .Y(_08716_),
    .A1(_08303_),
    .A2(_08352_));
 sg13g2_nand2_1 _14601_ (.Y(_08717_),
    .A(_08655_),
    .B(_08716_));
 sg13g2_nor3_1 _14602_ (.A(net976),
    .B(net919),
    .C(_08542_),
    .Y(_08718_));
 sg13g2_a21o_1 _14603_ (.A2(_08717_),
    .A1(net938),
    .B1(_08718_),
    .X(_08719_));
 sg13g2_a22oi_1 _14604_ (.Y(_08720_),
    .B1(_08719_),
    .B2(net922),
    .A2(_08715_),
    .A1(net899));
 sg13g2_mux4_1 _14605_ (.S0(net977),
    .A0(_08704_),
    .A1(_08708_),
    .A2(_08710_),
    .A3(_08720_),
    .S1(net928),
    .X(_08721_));
 sg13g2_nor2_1 _14606_ (.A(net1001),
    .B(_08721_),
    .Y(_08722_));
 sg13g2_a21oi_1 _14607_ (.A1(net958),
    .A2(_08697_),
    .Y(_08723_),
    .B1(_08722_));
 sg13g2_nand2_1 _14608_ (.Y(_08724_),
    .A(\top_ihp.oisc.micro_op[15] ),
    .B(net843));
 sg13g2_o21ai_1 _14609_ (.B1(_08724_),
    .Y(_00275_),
    .A1(_08254_),
    .A2(_08723_));
 sg13g2_a22oi_1 _14610_ (.Y(_08725_),
    .B1(_08372_),
    .B2(net963),
    .A2(net1006),
    .A1(_08271_));
 sg13g2_o21ai_1 _14611_ (.B1(net972),
    .Y(_08726_),
    .A1(net1006),
    .A2(_08396_));
 sg13g2_nand2_1 _14612_ (.Y(_08727_),
    .A(_08725_),
    .B(_08726_));
 sg13g2_a22oi_1 _14613_ (.Y(_08728_),
    .B1(_08727_),
    .B2(net925),
    .A2(_08407_),
    .A1(_08350_));
 sg13g2_nor2_1 _14614_ (.A(_08320_),
    .B(_08728_),
    .Y(_08729_));
 sg13g2_a21oi_1 _14615_ (.A1(_08511_),
    .A2(_08590_),
    .Y(_08730_),
    .B1(_08729_));
 sg13g2_nand2_1 _14616_ (.Y(_08731_),
    .A(net973),
    .B(_08491_));
 sg13g2_o21ai_1 _14617_ (.B1(_08731_),
    .Y(_08732_),
    .A1(net1004),
    .A2(_08444_));
 sg13g2_nand2_1 _14618_ (.Y(_08733_),
    .A(net974),
    .B(_08732_));
 sg13g2_o21ai_1 _14619_ (.B1(_08733_),
    .Y(_08734_),
    .A1(net975),
    .A2(net936));
 sg13g2_a21oi_1 _14620_ (.A1(_08622_),
    .A2(_08734_),
    .Y(_08735_),
    .B1(_08317_));
 sg13g2_a21oi_1 _14621_ (.A1(_08423_),
    .A2(_08730_),
    .Y(_08736_),
    .B1(_08735_));
 sg13g2_nand2_1 _14622_ (.Y(_08737_),
    .A(_08340_),
    .B(_08519_));
 sg13g2_a22oi_1 _14623_ (.Y(_08738_),
    .B1(_08737_),
    .B2(net891),
    .A2(_08637_),
    .A1(_08402_));
 sg13g2_nor2_1 _14624_ (.A(net889),
    .B(_08738_),
    .Y(_08739_));
 sg13g2_a22oi_1 _14625_ (.Y(_08740_),
    .B1(_08693_),
    .B2(net919),
    .A2(_08456_),
    .A1(net920));
 sg13g2_o21ai_1 _14626_ (.B1(_08443_),
    .Y(_08741_),
    .A1(net920),
    .A2(net960));
 sg13g2_o21ai_1 _14627_ (.B1(_08741_),
    .Y(_08742_),
    .A1(net900),
    .A2(_08740_));
 sg13g2_o21ai_1 _14628_ (.B1(net928),
    .Y(_08743_),
    .A1(_08739_),
    .A2(_08742_));
 sg13g2_nand2_1 _14629_ (.Y(_08744_),
    .A(net1010),
    .B(_08407_));
 sg13g2_o21ai_1 _14630_ (.B1(_08744_),
    .Y(_08745_),
    .A1(_08290_),
    .A2(_08467_));
 sg13g2_a21oi_1 _14631_ (.A1(net891),
    .A2(_08745_),
    .Y(_08746_),
    .B1(_08300_));
 sg13g2_nor2_1 _14632_ (.A(_08490_),
    .B(_08746_),
    .Y(_08747_));
 sg13g2_nor4_2 _14633_ (.A(net968),
    .B(net964),
    .C(_08363_),
    .Y(_08748_),
    .D(_08612_));
 sg13g2_nor2_1 _14634_ (.A(_08747_),
    .B(_08748_),
    .Y(_08749_));
 sg13g2_a21oi_1 _14635_ (.A1(_08743_),
    .A2(_08749_),
    .Y(_08750_),
    .B1(net977));
 sg13g2_a21oi_1 _14636_ (.A1(net977),
    .A2(_08736_),
    .Y(_08751_),
    .B1(_08750_));
 sg13g2_nand2_1 _14637_ (.Y(_08752_),
    .A(net892),
    .B(_08582_));
 sg13g2_a21oi_1 _14638_ (.A1(_08488_),
    .A2(_08646_),
    .Y(_08753_),
    .B1(net890));
 sg13g2_a21oi_1 _14639_ (.A1(_08369_),
    .A2(_08585_),
    .Y(_08754_),
    .B1(net895));
 sg13g2_nor2_1 _14640_ (.A(_08422_),
    .B(_08754_),
    .Y(_08755_));
 sg13g2_o21ai_1 _14641_ (.B1(_08755_),
    .Y(_08756_),
    .A1(_08752_),
    .A2(_08753_));
 sg13g2_nor2_1 _14642_ (.A(net919),
    .B(net964),
    .Y(_08757_));
 sg13g2_xnor2_1 _14643_ (.Y(_08758_),
    .A(_08551_),
    .B(_08757_));
 sg13g2_nor2_1 _14644_ (.A(_08391_),
    .B(_08456_),
    .Y(_08759_));
 sg13g2_a21o_1 _14645_ (.A2(_08529_),
    .A1(net921),
    .B1(net925),
    .X(_08760_));
 sg13g2_o21ai_1 _14646_ (.B1(_08358_),
    .Y(_08761_),
    .A1(_08590_),
    .A2(_08760_));
 sg13g2_nand3_1 _14647_ (.B(_08529_),
    .C(_08352_),
    .A(net966),
    .Y(_08762_));
 sg13g2_nand3_1 _14648_ (.B(_08698_),
    .C(_08688_),
    .A(_08328_),
    .Y(_08763_));
 sg13g2_nand3_1 _14649_ (.B(_08762_),
    .C(_08763_),
    .A(_08761_),
    .Y(_08764_));
 sg13g2_a221oi_1 _14650_ (.B2(net875),
    .C1(net1002),
    .B1(_08764_),
    .A1(_08758_),
    .Y(_08765_),
    .A2(_08759_));
 sg13g2_a21oi_1 _14651_ (.A1(net957),
    .A2(_08756_),
    .Y(_08766_),
    .B1(_08765_));
 sg13g2_nor2_1 _14652_ (.A(_08257_),
    .B(_08766_),
    .Y(_08767_));
 sg13g2_a21oi_1 _14653_ (.A1(_08257_),
    .A2(_08751_),
    .Y(_08768_),
    .B1(_08767_));
 sg13g2_mux2_1 _14654_ (.A0(_08768_),
    .A1(_07424_),
    .S(net843),
    .X(_00276_));
 sg13g2_inv_1 _14655_ (.Y(_08769_),
    .A(_08326_));
 sg13g2_a22oi_1 _14656_ (.Y(_08770_),
    .B1(_08769_),
    .B2(_08512_),
    .A2(_08334_),
    .A1(net898));
 sg13g2_nor2_1 _14657_ (.A(_08454_),
    .B(_08504_),
    .Y(_08771_));
 sg13g2_nor4_1 _14658_ (.A(_08386_),
    .B(_08502_),
    .C(_08570_),
    .D(_08771_),
    .Y(_08772_));
 sg13g2_a21oi_1 _14659_ (.A1(net876),
    .A2(_08770_),
    .Y(_08773_),
    .B1(_08772_));
 sg13g2_a21oi_1 _14660_ (.A1(_08542_),
    .A2(_08620_),
    .Y(_08774_),
    .B1(net923));
 sg13g2_a21o_1 _14661_ (.A2(_08396_),
    .A1(_08297_),
    .B1(_08774_),
    .X(_08775_));
 sg13g2_a21o_1 _14662_ (.A2(_08469_),
    .A1(net927),
    .B1(_08573_),
    .X(_08776_));
 sg13g2_a22oi_1 _14663_ (.Y(_08777_),
    .B1(_08776_),
    .B2(net897),
    .A2(_08775_),
    .A1(net889));
 sg13g2_nor2_1 _14664_ (.A(net931),
    .B(_08777_),
    .Y(_08778_));
 sg13g2_a21oi_1 _14665_ (.A1(net924),
    .A2(_08773_),
    .Y(_08779_),
    .B1(_08778_));
 sg13g2_a21oi_1 _14666_ (.A1(net969),
    .A2(net960),
    .Y(_08780_),
    .B1(_08520_));
 sg13g2_nand2_1 _14667_ (.Y(_08781_),
    .A(net1008),
    .B(net963));
 sg13g2_a21oi_1 _14668_ (.A1(_08504_),
    .A2(_08469_),
    .Y(_08782_),
    .B1(_08781_));
 sg13g2_nor2_1 _14669_ (.A(_08342_),
    .B(_08782_),
    .Y(_08783_));
 sg13g2_o21ai_1 _14670_ (.B1(_08783_),
    .Y(_08784_),
    .A1(_08363_),
    .A2(_08780_));
 sg13g2_nand2_1 _14671_ (.Y(_08785_),
    .A(_08259_),
    .B(_08784_));
 sg13g2_or2_1 _14672_ (.X(_08786_),
    .B(_08785_),
    .A(_08735_));
 sg13g2_buf_1 _14673_ (.A(_08786_),
    .X(_08787_));
 sg13g2_o21ai_1 _14674_ (.B1(_08787_),
    .Y(_08788_),
    .A1(net977),
    .A2(_08779_));
 sg13g2_nand2_1 _14675_ (.Y(_08789_),
    .A(net920),
    .B(_08325_));
 sg13g2_o21ai_1 _14676_ (.B1(_08789_),
    .Y(_08790_),
    .A1(net1011),
    .A2(net890));
 sg13g2_xnor2_1 _14677_ (.Y(_08791_),
    .A(net929),
    .B(_08444_));
 sg13g2_o21ai_1 _14678_ (.B1(_08539_),
    .Y(_08792_),
    .A1(_08387_),
    .A2(_08637_));
 sg13g2_o21ai_1 _14679_ (.B1(_08792_),
    .Y(_08793_),
    .A1(net894),
    .A2(_08791_));
 sg13g2_a22oi_1 _14680_ (.Y(_08794_),
    .B1(_08793_),
    .B2(net875),
    .A2(_08790_),
    .A1(_08371_));
 sg13g2_or2_1 _14681_ (.X(_08795_),
    .B(_08794_),
    .A(_08379_));
 sg13g2_a22oi_1 _14682_ (.Y(_08796_),
    .B1(_08402_),
    .B2(_08637_),
    .A2(_08400_),
    .A1(net937));
 sg13g2_a21oi_1 _14683_ (.A1(_08403_),
    .A2(_08387_),
    .Y(_08797_),
    .B1(net938));
 sg13g2_a21oi_1 _14684_ (.A1(net889),
    .A2(_08796_),
    .Y(_08798_),
    .B1(_08797_));
 sg13g2_nand2_1 _14685_ (.Y(_08799_),
    .A(_08301_),
    .B(_08340_));
 sg13g2_a22oi_1 _14686_ (.Y(_08800_),
    .B1(_08631_),
    .B2(_08799_),
    .A2(net934),
    .A1(net920));
 sg13g2_nor3_1 _14687_ (.A(net874),
    .B(net959),
    .C(_08800_),
    .Y(_08801_));
 sg13g2_a21oi_1 _14688_ (.A1(net959),
    .A2(_08798_),
    .Y(_08802_),
    .B1(_08801_));
 sg13g2_or2_1 _14689_ (.X(_08803_),
    .B(_08802_),
    .A(_08435_));
 sg13g2_nand3_1 _14690_ (.B(_08795_),
    .C(_08803_),
    .A(net1001),
    .Y(_08804_));
 sg13g2_o21ai_1 _14691_ (.B1(_08804_),
    .Y(_08805_),
    .A1(net958),
    .A2(_08788_));
 sg13g2_nand2_1 _14692_ (.Y(_08806_),
    .A(_07430_),
    .B(net843));
 sg13g2_o21ai_1 _14693_ (.B1(_08806_),
    .Y(_00277_),
    .A1(net844),
    .A2(_08805_));
 sg13g2_o21ai_1 _14694_ (.B1(_08534_),
    .Y(_08807_),
    .A1(net975),
    .A2(_08533_));
 sg13g2_a22oi_1 _14695_ (.Y(_08808_),
    .B1(_08807_),
    .B2(net976),
    .A2(_08352_),
    .A1(net897));
 sg13g2_inv_1 _14696_ (.Y(_08809_),
    .A(_08808_));
 sg13g2_a22oi_1 _14697_ (.Y(_08810_),
    .B1(_08809_),
    .B2(_08348_),
    .A2(_08511_),
    .A1(_08498_));
 sg13g2_nor2_1 _14698_ (.A(net959),
    .B(_08810_),
    .Y(_08811_));
 sg13g2_o21ai_1 _14699_ (.B1(net1002),
    .Y(_08812_),
    .A1(_08747_),
    .A2(_08811_));
 sg13g2_nand2_1 _14700_ (.Y(_08813_),
    .A(_08787_),
    .B(_08812_));
 sg13g2_nor3_1 _14701_ (.A(_08538_),
    .B(net927),
    .C(_08357_),
    .Y(_08814_));
 sg13g2_a21oi_1 _14702_ (.A1(net892),
    .A2(_08590_),
    .Y(_08815_),
    .B1(_08814_));
 sg13g2_and2_1 _14703_ (.A(_08338_),
    .B(_08476_),
    .X(_08816_));
 sg13g2_a21oi_1 _14704_ (.A1(_08439_),
    .A2(_08816_),
    .Y(_08817_),
    .B1(_08748_));
 sg13g2_o21ai_1 _14705_ (.B1(_08817_),
    .Y(_08818_),
    .A1(_08677_),
    .A2(_08815_));
 sg13g2_nor2_1 _14706_ (.A(_08653_),
    .B(net890),
    .Y(_08819_));
 sg13g2_a21o_1 _14707_ (.A2(_08819_),
    .A1(net1011),
    .B1(_08474_),
    .X(_08820_));
 sg13g2_nor2_1 _14708_ (.A(_08475_),
    .B(_08379_),
    .Y(_08821_));
 sg13g2_a22oi_1 _14709_ (.Y(_08822_),
    .B1(_08820_),
    .B2(_08821_),
    .A2(_08818_),
    .A1(net977));
 sg13g2_nand2_1 _14710_ (.Y(_08823_),
    .A(net1001),
    .B(_08822_));
 sg13g2_o21ai_1 _14711_ (.B1(_08823_),
    .Y(_08824_),
    .A1(_08465_),
    .A2(_08813_));
 sg13g2_nand2_1 _14712_ (.Y(_08825_),
    .A(_07429_),
    .B(_08253_));
 sg13g2_o21ai_1 _14713_ (.B1(_08825_),
    .Y(_00278_),
    .A1(net844),
    .A2(_08824_));
 sg13g2_inv_1 _14714_ (.Y(_08826_),
    .A(_07426_));
 sg13g2_nor3_1 _14715_ (.A(net895),
    .B(_08454_),
    .C(_08612_),
    .Y(_08827_));
 sg13g2_a21oi_1 _14716_ (.A1(net876),
    .A2(_08820_),
    .Y(_08828_),
    .B1(_08827_));
 sg13g2_nand2_1 _14717_ (.Y(_08829_),
    .A(net1010),
    .B(net971));
 sg13g2_nor2_1 _14718_ (.A(_08270_),
    .B(net974),
    .Y(_08830_));
 sg13g2_a21oi_1 _14719_ (.A1(_08271_),
    .A2(_08473_),
    .Y(_08831_),
    .B1(_08830_));
 sg13g2_nand3_1 _14720_ (.B(_08333_),
    .C(_08473_),
    .A(net962),
    .Y(_08832_));
 sg13g2_o21ai_1 _14721_ (.B1(_08832_),
    .Y(_08833_),
    .A1(_08829_),
    .A2(_08831_));
 sg13g2_a221oi_1 _14722_ (.B2(net900),
    .C1(_08748_),
    .B1(_08833_),
    .A1(_08361_),
    .Y(_08834_),
    .A2(_08511_));
 sg13g2_or2_1 _14723_ (.X(_08835_),
    .B(_08834_),
    .A(net1003));
 sg13g2_o21ai_1 _14724_ (.B1(_08835_),
    .Y(_08836_),
    .A1(_08379_),
    .A2(_08828_));
 sg13g2_a21o_1 _14725_ (.A2(_08836_),
    .A1(net1001),
    .B1(_08253_),
    .X(_08837_));
 sg13g2_a21oi_1 _14726_ (.A1(net875),
    .A2(_08586_),
    .Y(_08838_),
    .B1(_08490_));
 sg13g2_o21ai_1 _14727_ (.B1(_08466_),
    .Y(_08839_),
    .A1(_08811_),
    .A2(_08838_));
 sg13g2_a21oi_1 _14728_ (.A1(_08787_),
    .A2(_08839_),
    .Y(_08840_),
    .B1(net958));
 sg13g2_nor2_1 _14729_ (.A(_08837_),
    .B(_08840_),
    .Y(_08841_));
 sg13g2_a21oi_1 _14730_ (.A1(_08826_),
    .A2(_08251_),
    .Y(_00279_),
    .B1(_08841_));
 sg13g2_inv_1 _14731_ (.Y(_08842_),
    .A(_07431_));
 sg13g2_a21oi_1 _14732_ (.A1(net978),
    .A2(_08813_),
    .Y(_08843_),
    .B1(_08837_));
 sg13g2_a21oi_1 _14733_ (.A1(_08842_),
    .A2(net844),
    .Y(_00280_),
    .B1(_08843_));
 sg13g2_o21ai_1 _14734_ (.B1(_08533_),
    .Y(_08844_),
    .A1(_08407_),
    .A2(_08829_));
 sg13g2_nand3_1 _14735_ (.B(net965),
    .C(_08529_),
    .A(net921),
    .Y(_08845_));
 sg13g2_o21ai_1 _14736_ (.B1(_08845_),
    .Y(_08846_),
    .A1(net890),
    .A2(_08527_));
 sg13g2_a21oi_1 _14737_ (.A1(net901),
    .A2(_08844_),
    .Y(_08847_),
    .B1(_08846_));
 sg13g2_nand2_1 _14738_ (.Y(_08848_),
    .A(_08427_),
    .B(_08439_));
 sg13g2_o21ai_1 _14739_ (.B1(_08848_),
    .Y(_08849_),
    .A1(net937),
    .A2(net1000));
 sg13g2_a21oi_1 _14740_ (.A1(net893),
    .A2(_08849_),
    .Y(_08850_),
    .B1(net895));
 sg13g2_a21oi_1 _14741_ (.A1(net876),
    .A2(_08847_),
    .Y(_08851_),
    .B1(_08850_));
 sg13g2_nand3b_1 _14742_ (.B(net972),
    .C(_08456_),
    .Y(_08852_),
    .A_N(_08830_));
 sg13g2_o21ai_1 _14743_ (.B1(_08852_),
    .Y(_08853_),
    .A1(net929),
    .A2(_08456_));
 sg13g2_a221oi_1 _14744_ (.B2(net888),
    .C1(net900),
    .B1(_08853_),
    .A1(net927),
    .Y(_08854_),
    .A2(net963));
 sg13g2_a21oi_1 _14745_ (.A1(net923),
    .A2(net968),
    .Y(_08855_),
    .B1(_08388_));
 sg13g2_nor2_1 _14746_ (.A(net920),
    .B(_08855_),
    .Y(_08856_));
 sg13g2_a21oi_1 _14747_ (.A1(net921),
    .A2(_08418_),
    .Y(_08857_),
    .B1(net927));
 sg13g2_a21oi_1 _14748_ (.A1(net1000),
    .A2(_08338_),
    .Y(_08858_),
    .B1(net935));
 sg13g2_nor2_1 _14749_ (.A(_08857_),
    .B(_08858_),
    .Y(_08859_));
 sg13g2_nor3_1 _14750_ (.A(net894),
    .B(_08856_),
    .C(_08859_),
    .Y(_08860_));
 sg13g2_o21ai_1 _14751_ (.B1(net931),
    .Y(_08861_),
    .A1(_08854_),
    .A2(_08860_));
 sg13g2_o21ai_1 _14752_ (.B1(_08861_),
    .Y(_08862_),
    .A1(net931),
    .A2(_08851_));
 sg13g2_o21ai_1 _14753_ (.B1(_08373_),
    .Y(_08863_),
    .A1(net929),
    .A2(net936));
 sg13g2_a21oi_1 _14754_ (.A1(net921),
    .A2(_08405_),
    .Y(_08864_),
    .B1(_08371_));
 sg13g2_nand2_1 _14755_ (.Y(_08865_),
    .A(_08321_),
    .B(_08473_));
 sg13g2_o21ai_1 _14756_ (.B1(_08865_),
    .Y(_08866_),
    .A1(net933),
    .A2(_08864_));
 sg13g2_a22oi_1 _14757_ (.Y(_08867_),
    .B1(_08866_),
    .B2(net874),
    .A2(_08863_),
    .A1(_08611_));
 sg13g2_a21oi_1 _14758_ (.A1(_08266_),
    .A2(_08444_),
    .Y(_08868_),
    .B1(_08555_));
 sg13g2_o21ai_1 _14759_ (.B1(_08446_),
    .Y(_08869_),
    .A1(net966),
    .A2(_08868_));
 sg13g2_o21ai_1 _14760_ (.B1(_08405_),
    .Y(_08870_),
    .A1(_08321_),
    .A2(_08418_));
 sg13g2_nor3_1 _14761_ (.A(net900),
    .B(_08590_),
    .C(_08870_),
    .Y(_08871_));
 sg13g2_a21oi_1 _14762_ (.A1(net899),
    .A2(_08869_),
    .Y(_08872_),
    .B1(_08871_));
 sg13g2_o21ai_1 _14763_ (.B1(_08872_),
    .Y(_08873_),
    .A1(net894),
    .A2(_08867_));
 sg13g2_a21o_1 _14764_ (.A2(net898),
    .A1(net922),
    .B1(_08325_),
    .X(_08874_));
 sg13g2_nand4_1 _14765_ (.B(net964),
    .C(net1023),
    .A(net892),
    .Y(_08875_),
    .D(_08848_));
 sg13g2_a221oi_1 _14766_ (.B2(net902),
    .C1(_08875_),
    .B1(_08874_),
    .A1(_08292_),
    .Y(_08876_),
    .A2(_08326_));
 sg13g2_a21oi_1 _14767_ (.A1(net1002),
    .A2(_08873_),
    .Y(_08877_),
    .B1(_08876_));
 sg13g2_o21ai_1 _14768_ (.B1(_08877_),
    .Y(_08878_),
    .A1(net957),
    .A2(_08862_));
 sg13g2_nor2_1 _14769_ (.A(_08314_),
    .B(_08485_),
    .Y(_08879_));
 sg13g2_a21oi_1 _14770_ (.A1(net926),
    .A2(_08439_),
    .Y(_08880_),
    .B1(_08879_));
 sg13g2_nand2_1 _14771_ (.Y(_08881_),
    .A(_08328_),
    .B(_08848_));
 sg13g2_a21oi_1 _14772_ (.A1(net889),
    .A2(_08881_),
    .Y(_08882_),
    .B1(_08442_));
 sg13g2_a22oi_1 _14773_ (.Y(_08883_),
    .B1(_08599_),
    .B2(net888),
    .A2(net898),
    .A1(net922));
 sg13g2_a221oi_1 _14774_ (.B2(_08883_),
    .C1(_08366_),
    .B1(_08882_),
    .A1(_08426_),
    .Y(_08884_),
    .A2(_08880_));
 sg13g2_nand3_1 _14775_ (.B(net968),
    .C(_08488_),
    .A(_08298_),
    .Y(_08885_));
 sg13g2_o21ai_1 _14776_ (.B1(_08885_),
    .Y(_08886_),
    .A1(net934),
    .A2(_08527_));
 sg13g2_nand3_1 _14777_ (.B(net968),
    .C(net890),
    .A(net1020),
    .Y(_08887_));
 sg13g2_o21ai_1 _14778_ (.B1(_08887_),
    .Y(_08888_),
    .A1(net934),
    .A2(_08363_));
 sg13g2_a22oi_1 _14779_ (.Y(_08889_),
    .B1(_08888_),
    .B2(net932),
    .A2(_08886_),
    .A1(net963));
 sg13g2_o21ai_1 _14780_ (.B1(_08889_),
    .Y(_08890_),
    .A1(_08414_),
    .A2(_08395_));
 sg13g2_o21ai_1 _14781_ (.B1(net921),
    .Y(_08891_),
    .A1(_08297_),
    .A2(_08511_));
 sg13g2_nor2b_1 _14782_ (.A(_08287_),
    .B_N(_08891_),
    .Y(_08892_));
 sg13g2_nor3_1 _14783_ (.A(net889),
    .B(_08259_),
    .C(_08892_),
    .Y(_08893_));
 sg13g2_a21oi_1 _14784_ (.A1(_08259_),
    .A2(_08890_),
    .Y(_08894_),
    .B1(_08893_));
 sg13g2_nor2_1 _14785_ (.A(net931),
    .B(_08894_),
    .Y(_08895_));
 sg13g2_a21oi_1 _14786_ (.A1(net924),
    .A2(_08884_),
    .Y(_08896_),
    .B1(_08895_));
 sg13g2_nand2_1 _14787_ (.Y(_08897_),
    .A(net1001),
    .B(_08896_));
 sg13g2_o21ai_1 _14788_ (.B1(_08897_),
    .Y(_08898_),
    .A1(net958),
    .A2(_08878_));
 sg13g2_nand2_1 _14789_ (.Y(_08899_),
    .A(_08232_),
    .B(_08253_));
 sg13g2_o21ai_1 _14790_ (.B1(_08899_),
    .Y(_00281_),
    .A1(net844),
    .A2(_08898_));
 sg13g2_nor2_1 _14791_ (.A(net930),
    .B(net1005),
    .Y(_08900_));
 sg13g2_a21o_1 _14792_ (.A2(_08900_),
    .A1(net901),
    .B1(_08499_),
    .X(_08901_));
 sg13g2_a22oi_1 _14793_ (.Y(_08902_),
    .B1(_08901_),
    .B2(net902),
    .A2(_08900_),
    .A1(net926));
 sg13g2_nor2_1 _14794_ (.A(_08305_),
    .B(net964),
    .Y(_08903_));
 sg13g2_o21ai_1 _14795_ (.B1(_08449_),
    .Y(_08904_),
    .A1(net898),
    .A2(_08903_));
 sg13g2_a21oi_1 _14796_ (.A1(_08683_),
    .A2(_08904_),
    .Y(_08905_),
    .B1(net889));
 sg13g2_nand3_1 _14797_ (.B(net964),
    .C(_08631_),
    .A(net1000),
    .Y(_08906_));
 sg13g2_a21oi_1 _14798_ (.A1(_08683_),
    .A2(_08906_),
    .Y(_08907_),
    .B1(net874));
 sg13g2_nor3_1 _14799_ (.A(net894),
    .B(_08422_),
    .C(net896),
    .Y(_08908_));
 sg13g2_nor4_1 _14800_ (.A(net876),
    .B(_08905_),
    .C(_08907_),
    .D(_08908_),
    .Y(_08909_));
 sg13g2_a21oi_1 _14801_ (.A1(_08436_),
    .A2(_08902_),
    .Y(_08910_),
    .B1(_08909_));
 sg13g2_nor2_1 _14802_ (.A(net888),
    .B(_08323_),
    .Y(_08911_));
 sg13g2_a22oi_1 _14803_ (.Y(_08912_),
    .B1(_08789_),
    .B2(_08911_),
    .A2(_08530_),
    .A1(net888));
 sg13g2_a21o_1 _14804_ (.A2(_08331_),
    .A1(net975),
    .B1(_08711_),
    .X(_08913_));
 sg13g2_nand3_1 _14805_ (.B(_08731_),
    .C(_08713_),
    .A(net976),
    .Y(_08914_));
 sg13g2_o21ai_1 _14806_ (.B1(_08914_),
    .Y(_08915_),
    .A1(net920),
    .A2(_08913_));
 sg13g2_nor2_1 _14807_ (.A(net892),
    .B(_08915_),
    .Y(_08916_));
 sg13g2_a21oi_1 _14808_ (.A1(net875),
    .A2(_08912_),
    .Y(_08917_),
    .B1(_08916_));
 sg13g2_a21oi_1 _14809_ (.A1(net891),
    .A2(_08414_),
    .Y(_08918_),
    .B1(_08402_));
 sg13g2_nand2_1 _14810_ (.Y(_08919_),
    .A(_08443_),
    .B(_08403_));
 sg13g2_o21ai_1 _14811_ (.B1(_08919_),
    .Y(_08920_),
    .A1(net888),
    .A2(_08918_));
 sg13g2_a221oi_1 _14812_ (.B2(net902),
    .C1(net931),
    .B1(_08920_),
    .A1(_08334_),
    .Y(_08921_),
    .A2(_08514_));
 sg13g2_a21oi_1 _14813_ (.A1(net924),
    .A2(_08917_),
    .Y(_08922_),
    .B1(_08921_));
 sg13g2_o21ai_1 _14814_ (.B1(_08662_),
    .Y(_08923_),
    .A1(_08398_),
    .A2(_08661_));
 sg13g2_nand3_1 _14815_ (.B(_08377_),
    .C(_08371_),
    .A(_08359_),
    .Y(_08924_));
 sg13g2_a21oi_1 _14816_ (.A1(_08923_),
    .A2(_08924_),
    .Y(_08925_),
    .B1(net924));
 sg13g2_a221oi_1 _14817_ (.B2(net888),
    .C1(_08325_),
    .B1(_08501_),
    .A1(net898),
    .Y(_08926_),
    .A2(_08338_));
 sg13g2_nand2_1 _14818_ (.Y(_08927_),
    .A(net959),
    .B(_08915_));
 sg13g2_o21ai_1 _14819_ (.B1(_08927_),
    .Y(_08928_),
    .A1(net931),
    .A2(_08926_));
 sg13g2_nor2_1 _14820_ (.A(_08395_),
    .B(_08602_),
    .Y(_08929_));
 sg13g2_a21oi_1 _14821_ (.A1(net969),
    .A2(_08611_),
    .Y(_08930_),
    .B1(_08450_));
 sg13g2_nor2_1 _14822_ (.A(_08653_),
    .B(_08683_),
    .Y(_08931_));
 sg13g2_o21ai_1 _14823_ (.B1(_08369_),
    .Y(_08932_),
    .A1(_08900_),
    .A2(_08931_));
 sg13g2_o21ai_1 _14824_ (.B1(_08932_),
    .Y(_08933_),
    .A1(_08445_),
    .A2(_08930_));
 sg13g2_nor3_1 _14825_ (.A(net875),
    .B(_08929_),
    .C(_08933_),
    .Y(_08934_));
 sg13g2_a21oi_1 _14826_ (.A1(_08436_),
    .A2(_08928_),
    .Y(_08935_),
    .B1(_08934_));
 sg13g2_mux4_1 _14827_ (.S0(net978),
    .A0(_08910_),
    .A1(_08922_),
    .A2(_08925_),
    .A3(_08935_),
    .S1(net957),
    .X(_08936_));
 sg13g2_mux2_1 _14828_ (.A0(_08936_),
    .A1(_08227_),
    .S(net843),
    .X(_00282_));
 sg13g2_nand2_1 _14829_ (.Y(_08937_),
    .A(net1016),
    .B(\top_ihp.oisc.micro_state[2] ));
 sg13g2_nand2_1 _14830_ (.Y(_08938_),
    .A(_00074_),
    .B(_08937_));
 sg13g2_buf_1 _14831_ (.A(net1089),
    .X(_08939_));
 sg13g2_o21ai_1 _14832_ (.B1(_08939_),
    .Y(_08940_),
    .A1(_07436_),
    .A2(_08938_));
 sg13g2_buf_2 _14833_ (.A(_08940_),
    .X(_08941_));
 sg13g2_buf_1 _14834_ (.A(_08941_),
    .X(_08942_));
 sg13g2_buf_2 _14835_ (.A(\top_ihp.oisc.state[3] ),
    .X(_08943_));
 sg13g2_buf_1 _14836_ (.A(_08943_),
    .X(_08944_));
 sg13g2_inv_1 _14837_ (.Y(_08945_),
    .A(_07425_));
 sg13g2_buf_2 _14838_ (.A(\top_ihp.oisc.op_a[31] ),
    .X(_08946_));
 sg13g2_nor2b_1 _14839_ (.A(\top_ihp.oisc.op_b[31] ),
    .B_N(_08946_),
    .Y(_08947_));
 sg13g2_xnor2_1 _14840_ (.Y(_08948_),
    .A(\top_ihp.oisc.op_b[31] ),
    .B(_08946_));
 sg13g2_nor3_1 _14841_ (.A(_07720_),
    .B(_07844_),
    .C(_07916_),
    .Y(_08949_));
 sg13g2_and2_1 _14842_ (.A(_08948_),
    .B(_08949_),
    .X(_08950_));
 sg13g2_buf_1 _14843_ (.A(_08950_),
    .X(_08951_));
 sg13g2_nor2b_1 _14844_ (.A(_07699_),
    .B_N(_08951_),
    .Y(_08952_));
 sg13g2_and3_1 _14845_ (.X(_08953_),
    .A(_07598_),
    .B(_07611_),
    .C(_08952_));
 sg13g2_nand2b_1 _14846_ (.Y(_08954_),
    .B(net1026),
    .A_N(_07726_));
 sg13g2_nor2b_1 _14847_ (.A(net1026),
    .B_N(_07726_),
    .Y(_08955_));
 sg13g2_a21oi_1 _14848_ (.A1(_07719_),
    .A2(_08954_),
    .Y(_08956_),
    .B1(_08955_));
 sg13g2_nor2b_1 _14849_ (.A(_08956_),
    .B_N(_08948_),
    .Y(_08957_));
 sg13g2_a21o_1 _14850_ (.A2(_08951_),
    .A1(_07718_),
    .B1(_08957_),
    .X(_08958_));
 sg13g2_nor3_1 _14851_ (.A(_08947_),
    .B(_08953_),
    .C(_08958_),
    .Y(_08959_));
 sg13g2_xor2_1 _14852_ (.B(net1044),
    .A(_07444_),
    .X(_08960_));
 sg13g2_xnor2_1 _14853_ (.Y(_08961_),
    .A(net1037),
    .B(_07485_));
 sg13g2_nand3_1 _14854_ (.B(_07479_),
    .C(_08961_),
    .A(_07476_),
    .Y(_08962_));
 sg13g2_nor4_1 _14855_ (.A(_08960_),
    .B(_07493_),
    .C(_07480_),
    .D(_08962_),
    .Y(_08963_));
 sg13g2_or4_1 _14856_ (.A(_07464_),
    .B(_07603_),
    .C(_07607_),
    .D(_07608_),
    .X(_08964_));
 sg13g2_buf_1 _14857_ (.A(_08964_),
    .X(_08965_));
 sg13g2_nor4_1 _14858_ (.A(_08965_),
    .B(_07499_),
    .C(_08171_),
    .D(_08947_),
    .Y(_08966_));
 sg13g2_and4_1 _14859_ (.A(_07853_),
    .B(_07556_),
    .C(_08963_),
    .D(_08966_),
    .X(_08967_));
 sg13g2_nand3b_1 _14860_ (.B(_08951_),
    .C(_08967_),
    .Y(_08968_),
    .A_N(_07843_));
 sg13g2_buf_1 _14861_ (.A(_08968_),
    .X(_08969_));
 sg13g2_nand2b_1 _14862_ (.Y(_08970_),
    .B(_08969_),
    .A_N(_08959_));
 sg13g2_buf_2 _14863_ (.A(_08970_),
    .X(_08971_));
 sg13g2_nand2_1 _14864_ (.Y(_08972_),
    .A(_08945_),
    .B(_08971_));
 sg13g2_nor3_1 _14865_ (.A(_08943_),
    .B(net879),
    .C(_08937_),
    .Y(_08973_));
 sg13g2_buf_1 _14866_ (.A(_08973_),
    .X(_08974_));
 sg13g2_and2_1 _14867_ (.A(_08429_),
    .B(net842),
    .X(_08975_));
 sg13g2_a22oi_1 _14868_ (.Y(_08976_),
    .B1(_08972_),
    .B2(_08975_),
    .A2(\top_ihp.oisc.decoder.decoded[0] ),
    .A1(net999));
 sg13g2_and3_1 _14869_ (.X(_08977_),
    .A(_08945_),
    .B(_08971_),
    .C(net842));
 sg13g2_o21ai_1 _14870_ (.B1(_08268_),
    .Y(_08978_),
    .A1(_08941_),
    .A2(_08977_));
 sg13g2_o21ai_1 _14871_ (.B1(_08978_),
    .Y(_00283_),
    .A1(net822),
    .A2(_08976_));
 sg13g2_nand3b_1 _14872_ (.B(net842),
    .C(_08510_),
    .Y(_08979_),
    .A_N(_08941_));
 sg13g2_nand2_1 _14873_ (.Y(_08980_),
    .A(_08522_),
    .B(net842));
 sg13g2_or2_1 _14874_ (.X(_08981_),
    .B(_08958_),
    .A(_08953_));
 sg13g2_buf_1 _14875_ (.A(_08981_),
    .X(_08982_));
 sg13g2_nand3_1 _14876_ (.B(_07425_),
    .C(_08622_),
    .A(_07424_),
    .Y(_08983_));
 sg13g2_nand2_1 _14877_ (.Y(_08984_),
    .A(_07424_),
    .B(_08983_));
 sg13g2_nor3_1 _14878_ (.A(_08947_),
    .B(_08982_),
    .C(_08984_),
    .Y(_08985_));
 sg13g2_nand2_1 _14879_ (.Y(_08986_),
    .A(_08268_),
    .B(_08969_));
 sg13g2_nor2_1 _14880_ (.A(_08959_),
    .B(_08986_),
    .Y(_08987_));
 sg13g2_nand3_1 _14881_ (.B(net902),
    .C(_08983_),
    .A(_07425_),
    .Y(_08988_));
 sg13g2_o21ai_1 _14882_ (.B1(_08988_),
    .Y(_08989_),
    .A1(_08969_),
    .A2(_08984_));
 sg13g2_nor3_1 _14883_ (.A(_08985_),
    .B(_08987_),
    .C(_08989_),
    .Y(_08990_));
 sg13g2_mux2_1 _14884_ (.A0(_08979_),
    .A1(_08980_),
    .S(_08990_),
    .X(_08991_));
 sg13g2_inv_1 _14885_ (.Y(_08992_),
    .A(_08943_));
 sg13g2_inv_1 _14886_ (.Y(_08993_),
    .A(\top_ihp.oisc.decoder.decoded[1] ));
 sg13g2_nor3_1 _14887_ (.A(_08992_),
    .B(_08993_),
    .C(_08941_),
    .Y(_08994_));
 sg13g2_a21oi_1 _14888_ (.A1(_08522_),
    .A2(_08941_),
    .Y(_08995_),
    .B1(_08994_));
 sg13g2_nand2_1 _14889_ (.Y(_00284_),
    .A(_08991_),
    .B(_08995_));
 sg13g2_xnor2_1 _14890_ (.Y(_08996_),
    .A(net1000),
    .B(_08377_));
 sg13g2_a21o_1 _14891_ (.A2(_08264_),
    .A1(_07425_),
    .B1(_08269_),
    .X(_08997_));
 sg13g2_a22oi_1 _14892_ (.Y(_08998_),
    .B1(_08997_),
    .B2(_07424_),
    .A2(net961),
    .A1(_07425_));
 sg13g2_xor2_1 _14893_ (.B(_08605_),
    .A(_07430_),
    .X(_08999_));
 sg13g2_xnor2_1 _14894_ (.Y(_09000_),
    .A(_08998_),
    .B(_08999_));
 sg13g2_mux2_1 _14895_ (.A0(_08996_),
    .A1(_09000_),
    .S(_08971_),
    .X(_09001_));
 sg13g2_a221oi_1 _14896_ (.B2(_09001_),
    .C1(_08941_),
    .B1(net842),
    .A1(net999),
    .Y(_09002_),
    .A2(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_a21oi_1 _14897_ (.A1(net930),
    .A2(net822),
    .Y(_00285_),
    .B1(_09002_));
 sg13g2_nor2_1 _14898_ (.A(_08529_),
    .B(_08395_),
    .Y(_09003_));
 sg13g2_xnor2_1 _14899_ (.Y(_09004_),
    .A(net1011),
    .B(_09003_));
 sg13g2_nand2_1 _14900_ (.Y(_09005_),
    .A(_07430_),
    .B(_08279_));
 sg13g2_nor2_1 _14901_ (.A(_07430_),
    .B(_08279_),
    .Y(_09006_));
 sg13g2_a21oi_2 _14902_ (.B1(_09006_),
    .Y(_09007_),
    .A2(_09005_),
    .A1(_08998_));
 sg13g2_xnor2_1 _14903_ (.Y(_09008_),
    .A(_07429_),
    .B(_08391_));
 sg13g2_xnor2_1 _14904_ (.Y(_09009_),
    .A(_09007_),
    .B(_09008_));
 sg13g2_mux2_1 _14905_ (.A0(_09004_),
    .A1(_09009_),
    .S(_08971_),
    .X(_09010_));
 sg13g2_a221oi_1 _14906_ (.B2(_09010_),
    .C1(_08941_),
    .B1(net842),
    .A1(net999),
    .Y(_09011_),
    .A2(\top_ihp.oisc.decoder.decoded[3] ));
 sg13g2_a21oi_1 _14907_ (.A1(net900),
    .A2(net822),
    .Y(_00286_),
    .B1(_09011_));
 sg13g2_nor2_1 _14908_ (.A(_08364_),
    .B(_08469_),
    .Y(_09012_));
 sg13g2_xnor2_1 _14909_ (.Y(_09013_),
    .A(_08475_),
    .B(_09012_));
 sg13g2_nand2_1 _14910_ (.Y(_09014_),
    .A(_08324_),
    .B(_09007_));
 sg13g2_o21ai_1 _14911_ (.B1(_07429_),
    .Y(_09015_),
    .A1(_08293_),
    .A2(_09007_));
 sg13g2_nand2_1 _14912_ (.Y(_09016_),
    .A(_09014_),
    .B(_09015_));
 sg13g2_xnor2_1 _14913_ (.Y(_09017_),
    .A(_07426_),
    .B(net892));
 sg13g2_xnor2_1 _14914_ (.Y(_09018_),
    .A(_09016_),
    .B(_09017_));
 sg13g2_mux2_1 _14915_ (.A0(_09013_),
    .A1(_09018_),
    .S(_08971_),
    .X(_09019_));
 sg13g2_a22oi_1 _14916_ (.Y(_09020_),
    .B1(net842),
    .B2(_09019_),
    .A2(\top_ihp.oisc.decoder.decoded[4] ),
    .A1(net999));
 sg13g2_nand2_1 _14917_ (.Y(_09021_),
    .A(net875),
    .B(net822));
 sg13g2_o21ai_1 _14918_ (.B1(_09021_),
    .Y(_00287_),
    .A1(net822),
    .A2(_09020_));
 sg13g2_nor3_1 _14919_ (.A(net900),
    .B(_08340_),
    .C(net896),
    .Y(_09022_));
 sg13g2_xnor2_1 _14920_ (.Y(_09023_),
    .A(_08263_),
    .B(_09022_));
 sg13g2_nor2_1 _14921_ (.A(_08306_),
    .B(_09016_),
    .Y(_09024_));
 sg13g2_a21oi_1 _14922_ (.A1(_08306_),
    .A2(_09016_),
    .Y(_09025_),
    .B1(_07426_));
 sg13g2_nor2_2 _14923_ (.A(_09024_),
    .B(_09025_),
    .Y(_09026_));
 sg13g2_nand2_1 _14924_ (.Y(_09027_),
    .A(_07431_),
    .B(_08343_));
 sg13g2_nand2_1 _14925_ (.Y(_09028_),
    .A(_08842_),
    .B(_08317_));
 sg13g2_and2_1 _14926_ (.A(_09027_),
    .B(_09028_),
    .X(_09029_));
 sg13g2_xnor2_1 _14927_ (.Y(_09030_),
    .A(_09026_),
    .B(_09029_));
 sg13g2_mux2_1 _14928_ (.A0(_09023_),
    .A1(_09030_),
    .S(_08971_),
    .X(_09031_));
 sg13g2_a22oi_1 _14929_ (.Y(_09032_),
    .B1(net842),
    .B2(_09031_),
    .A2(\top_ihp.oisc.decoder.decoded[5] ),
    .A1(net999));
 sg13g2_nand2_1 _14930_ (.Y(_09033_),
    .A(net924),
    .B(net822));
 sg13g2_o21ai_1 _14931_ (.B1(_09033_),
    .Y(_00288_),
    .A1(net822),
    .A2(_09032_));
 sg13g2_nor3_1 _14932_ (.A(_08340_),
    .B(_08364_),
    .C(_08683_),
    .Y(_09034_));
 sg13g2_xnor2_1 _14933_ (.Y(_09035_),
    .A(_00082_),
    .B(_09034_));
 sg13g2_mux2_1 _14934_ (.A0(_09027_),
    .A1(_09028_),
    .S(_09026_),
    .X(_09036_));
 sg13g2_xnor2_1 _14935_ (.Y(_09037_),
    .A(net1002),
    .B(_09036_));
 sg13g2_mux2_1 _14936_ (.A0(_09035_),
    .A1(_09037_),
    .S(_08971_),
    .X(_09038_));
 sg13g2_a22oi_1 _14937_ (.Y(_09039_),
    .B1(_08974_),
    .B2(_09038_),
    .A2(\top_ihp.oisc.decoder.decoded[6] ),
    .A1(net999));
 sg13g2_nand2_1 _14938_ (.Y(_09040_),
    .A(net957),
    .B(net822));
 sg13g2_o21ai_1 _14939_ (.B1(_09040_),
    .Y(_00289_),
    .A1(_08942_),
    .A2(_09039_));
 sg13g2_nand4_1 _14940_ (.B(net1003),
    .C(_08297_),
    .A(net959),
    .Y(_09041_),
    .D(_09003_));
 sg13g2_xor2_1 _14941_ (.B(_09041_),
    .A(_00081_),
    .X(_09042_));
 sg13g2_nand2_1 _14942_ (.Y(_09043_),
    .A(_07431_),
    .B(_08432_));
 sg13g2_nand3_1 _14943_ (.B(net966),
    .C(net1023),
    .A(_08842_),
    .Y(_09044_));
 sg13g2_mux2_1 _14944_ (.A0(_09043_),
    .A1(_09044_),
    .S(_09026_),
    .X(_09045_));
 sg13g2_xnor2_1 _14945_ (.Y(_09046_),
    .A(_08464_),
    .B(_09045_));
 sg13g2_mux2_1 _14946_ (.A0(_09042_),
    .A1(_09046_),
    .S(_08971_),
    .X(_09047_));
 sg13g2_a22oi_1 _14947_ (.Y(_09048_),
    .B1(_08974_),
    .B2(_09047_),
    .A2(\top_ihp.oisc.decoder.decoded[7] ),
    .A1(net999));
 sg13g2_nand2_1 _14948_ (.Y(_09049_),
    .A(_08465_),
    .B(_08941_));
 sg13g2_o21ai_1 _14949_ (.B1(_09049_),
    .Y(_00290_),
    .A1(_08942_),
    .A2(_09048_));
 sg13g2_inv_1 _14950_ (.Y(_09050_),
    .A(\top_ihp.oisc.micro_state[2] ));
 sg13g2_mux2_1 _14951_ (.A0(_13204_),
    .A1(_09050_),
    .S(net979),
    .X(_00291_));
 sg13g2_nand2b_1 _14952_ (.Y(_09051_),
    .B(_08228_),
    .A_N(net979));
 sg13g2_o21ai_1 _14953_ (.B1(_09051_),
    .Y(_00292_),
    .A1(net879),
    .A2(_08251_));
 sg13g2_nand2_1 _14954_ (.Y(_09052_),
    .A(_08237_),
    .B(net939));
 sg13g2_o21ai_1 _14955_ (.B1(_09052_),
    .Y(_00293_),
    .A1(net979),
    .A2(_09050_));
 sg13g2_inv_1 _14956_ (.Y(_09053_),
    .A(\top_ihp.oisc.regs[0][0] ));
 sg13g2_buf_1 _14957_ (.A(\top_ihp.oisc.state[4] ),
    .X(_09054_));
 sg13g2_buf_1 _14958_ (.A(\top_ihp.oisc.decoder.instruction[8] ),
    .X(_09055_));
 sg13g2_nand2_1 _14959_ (.Y(_09056_),
    .A(_07420_),
    .B(_08241_));
 sg13g2_buf_1 _14960_ (.A(_09056_),
    .X(_09057_));
 sg13g2_buf_1 _14961_ (.A(\top_ihp.oisc.decoder.decoded[12] ),
    .X(_09058_));
 sg13g2_nand4_1 _14962_ (.B(_09058_),
    .C(_07428_),
    .A(net1016),
    .Y(_09059_),
    .D(_07433_));
 sg13g2_buf_1 _14963_ (.A(\top_ihp.oisc.decoder.decoded[14] ),
    .X(_09060_));
 sg13g2_buf_1 _14964_ (.A(\top_ihp.oisc.decoder.decoded[13] ),
    .X(_09061_));
 sg13g2_xor2_1 _14965_ (.B(_09061_),
    .A(_09060_),
    .X(_09062_));
 sg13g2_buf_2 _14966_ (.A(_00073_),
    .X(_09063_));
 sg13g2_a22oi_1 _14967_ (.Y(_09064_),
    .B1(_09062_),
    .B2(_09063_),
    .A2(_09059_),
    .A1(_09057_));
 sg13g2_buf_1 _14968_ (.A(_09064_),
    .X(_09065_));
 sg13g2_a221oi_1 _14969_ (.B2(_09058_),
    .C1(_08937_),
    .B1(net879),
    .A1(_07420_),
    .Y(_09066_),
    .A2(_08241_));
 sg13g2_buf_2 _14970_ (.A(_09066_),
    .X(_09067_));
 sg13g2_a22oi_1 _14971_ (.Y(_09068_),
    .B1(_09067_),
    .B2(\top_ihp.oisc.micro_res_addr[1] ),
    .A2(_09065_),
    .A1(_09055_));
 sg13g2_nand2b_1 _14972_ (.Y(_09069_),
    .B(_00074_),
    .A_N(_09068_));
 sg13g2_buf_1 _14973_ (.A(\top_ihp.oisc.state[2] ),
    .X(_09070_));
 sg13g2_buf_1 _14974_ (.A(_09070_),
    .X(_09071_));
 sg13g2_inv_1 _14975_ (.Y(_09072_),
    .A(net998));
 sg13g2_o21ai_1 _14976_ (.B1(_09072_),
    .Y(_09073_),
    .A1(net1019),
    .A2(_09069_));
 sg13g2_buf_1 _14977_ (.A(\top_ihp.oisc.decoder.instruction[7] ),
    .X(_09074_));
 sg13g2_a22oi_1 _14978_ (.Y(_09075_),
    .B1(_09067_),
    .B2(\top_ihp.oisc.micro_res_addr[0] ),
    .A2(_09065_),
    .A1(_09074_));
 sg13g2_nand2_1 _14979_ (.Y(_09076_),
    .A(_09072_),
    .B(_08992_));
 sg13g2_buf_1 _14980_ (.A(_09076_),
    .X(_09077_));
 sg13g2_nor2_1 _14981_ (.A(net1019),
    .B(_09077_),
    .Y(_09078_));
 sg13g2_nand2b_1 _14982_ (.Y(_09079_),
    .B(_09078_),
    .A_N(_09075_));
 sg13g2_buf_1 _14983_ (.A(_09079_),
    .X(_09080_));
 sg13g2_nand2b_1 _14984_ (.Y(_09081_),
    .B(_09080_),
    .A_N(_09073_));
 sg13g2_buf_2 _14985_ (.A(_09081_),
    .X(_09082_));
 sg13g2_buf_2 _14986_ (.A(_00075_),
    .X(_09083_));
 sg13g2_nor2_1 _14987_ (.A(_08943_),
    .B(net1019),
    .Y(_09084_));
 sg13g2_nand2_1 _14988_ (.Y(_09085_),
    .A(_09083_),
    .B(_09084_));
 sg13g2_nor2_1 _14989_ (.A(_09067_),
    .B(_09085_),
    .Y(_09086_));
 sg13g2_buf_1 _14990_ (.A(\top_ihp.oisc.decoder.instruction[11] ),
    .X(_09087_));
 sg13g2_nand4_1 _14991_ (.B(_09087_),
    .C(_09065_),
    .A(_09083_),
    .Y(_09088_),
    .D(_09084_));
 sg13g2_buf_2 _14992_ (.A(\top_ihp.oisc.state[0] ),
    .X(_09089_));
 sg13g2_buf_1 _14993_ (.A(_09089_),
    .X(_09090_));
 sg13g2_a21oi_1 _14994_ (.A1(_09058_),
    .A2(_08241_),
    .Y(_09091_),
    .B1(net997));
 sg13g2_nand3_1 _14995_ (.B(_09078_),
    .C(_09091_),
    .A(_08937_),
    .Y(_09092_));
 sg13g2_nand2_1 _14996_ (.Y(_09093_),
    .A(_09088_),
    .B(_09092_));
 sg13g2_nor2_1 _14997_ (.A(_09086_),
    .B(_09093_),
    .Y(_09094_));
 sg13g2_buf_2 _14998_ (.A(_09094_),
    .X(_09095_));
 sg13g2_buf_1 _14999_ (.A(\top_ihp.oisc.decoder.instruction[10] ),
    .X(_09096_));
 sg13g2_a22oi_1 _15000_ (.Y(_09097_),
    .B1(_09067_),
    .B2(\top_ihp.oisc.micro_res_addr[3] ),
    .A2(_09065_),
    .A1(_09096_));
 sg13g2_inv_1 _15001_ (.Y(_09098_),
    .A(_09097_));
 sg13g2_buf_1 _15002_ (.A(\top_ihp.oisc.decoder.instruction[9] ),
    .X(_09099_));
 sg13g2_nand2_1 _15003_ (.Y(_09100_),
    .A(_09099_),
    .B(_09065_));
 sg13g2_nand2_1 _15004_ (.Y(_09101_),
    .A(\top_ihp.oisc.micro_res_addr[2] ),
    .B(_09067_));
 sg13g2_nand3_1 _15005_ (.B(_09100_),
    .C(_09101_),
    .A(_09084_),
    .Y(_09102_));
 sg13g2_o21ai_1 _15006_ (.B1(_09083_),
    .Y(_09103_),
    .A1(_09098_),
    .A2(_09102_));
 sg13g2_buf_2 _15007_ (.A(_09103_),
    .X(_09104_));
 sg13g2_and2_1 _15008_ (.A(_09095_),
    .B(net737),
    .X(_09105_));
 sg13g2_buf_2 _15009_ (.A(_09105_),
    .X(_09106_));
 sg13g2_nor2b_1 _15010_ (.A(_09082_),
    .B_N(_09106_),
    .Y(_09107_));
 sg13g2_buf_1 _15011_ (.A(_09107_),
    .X(_09108_));
 sg13g2_buf_1 _15012_ (.A(_09061_),
    .X(_09109_));
 sg13g2_buf_1 _15013_ (.A(net996),
    .X(_09110_));
 sg13g2_buf_1 _15014_ (.A(_09063_),
    .X(_09111_));
 sg13g2_and3_1 _15015_ (.X(_09112_),
    .A(net956),
    .B(net995),
    .C(_09074_));
 sg13g2_nand3b_1 _15016_ (.B(\top_ihp.oisc.decoder.decoded[15] ),
    .C(net956),
    .Y(_09113_),
    .A_N(net995));
 sg13g2_inv_2 _15017_ (.Y(_09114_),
    .A(net996));
 sg13g2_nand2_1 _15018_ (.Y(_09115_),
    .A(_09114_),
    .B(_09063_));
 sg13g2_inv_1 _15019_ (.Y(_09116_),
    .A(\top_ihp.oisc.decoder.instruction[20] ));
 sg13g2_a21oi_1 _15020_ (.A1(_09113_),
    .A2(_09115_),
    .Y(_09117_),
    .B1(_09116_));
 sg13g2_buf_1 _15021_ (.A(_09060_),
    .X(_09118_));
 sg13g2_inv_1 _15022_ (.Y(_09119_),
    .A(net994));
 sg13g2_o21ai_1 _15023_ (.B1(_09119_),
    .Y(_09120_),
    .A1(_09112_),
    .A2(_09117_));
 sg13g2_inv_1 _15024_ (.Y(_09121_),
    .A(net1019));
 sg13g2_buf_1 _15025_ (.A(_09121_),
    .X(_09122_));
 sg13g2_buf_1 _15026_ (.A(_09077_),
    .X(_09123_));
 sg13g2_nor2_1 _15027_ (.A(net955),
    .B(net873),
    .Y(_09124_));
 sg13g2_buf_2 _15028_ (.A(\top_ihp.oisc.mem_addr_lowbits[0] ),
    .X(_09125_));
 sg13g2_nor2b_1 _15029_ (.A(_07822_),
    .B_N(_09125_),
    .Y(_09126_));
 sg13g2_buf_1 _15030_ (.A(_09126_),
    .X(_09127_));
 sg13g2_and2_1 _15031_ (.A(_08191_),
    .B(\top_ihp.wb_dati_spi[16] ),
    .X(_09128_));
 sg13g2_inv_1 _15032_ (.Y(_09129_),
    .A(\top_ihp.wb_dati_ram[16] ));
 sg13g2_nor4_1 _15033_ (.A(_08194_),
    .B(_09129_),
    .C(_08197_),
    .D(_08199_),
    .Y(_09130_));
 sg13g2_a221oi_1 _15034_ (.B2(_09128_),
    .C1(_09130_),
    .B1(_08190_),
    .A1(_08179_),
    .Y(_09131_),
    .A2(net878));
 sg13g2_nor2_1 _15035_ (.A(_07677_),
    .B(_08215_),
    .Y(_09132_));
 sg13g2_o21ai_1 _15036_ (.B1(_09132_),
    .Y(_09133_),
    .A1(\top_ihp.wb_dati_rom[16] ),
    .A2(_08205_));
 sg13g2_nor2_1 _15037_ (.A(_09131_),
    .B(_09133_),
    .Y(_09134_));
 sg13g2_buf_1 _15038_ (.A(_07823_),
    .X(_09135_));
 sg13g2_buf_1 _15039_ (.A(\top_ihp.oisc.mem_addr_lowbits[1] ),
    .X(_09136_));
 sg13g2_inv_1 _15040_ (.Y(_09137_),
    .A(net1018));
 sg13g2_buf_1 _15041_ (.A(_09137_),
    .X(_09138_));
 sg13g2_nor2_1 _15042_ (.A(net993),
    .B(_09138_),
    .Y(_09139_));
 sg13g2_buf_2 _15043_ (.A(_09139_),
    .X(_09140_));
 sg13g2_buf_1 _15044_ (.A(_08214_),
    .X(_09141_));
 sg13g2_nand2_1 _15045_ (.Y(_09142_),
    .A(\top_ihp.wb_dati_ram[0] ),
    .B(_09141_));
 sg13g2_buf_1 _15046_ (.A(net1012),
    .X(_09143_));
 sg13g2_buf_1 _15047_ (.A(net953),
    .X(_09144_));
 sg13g2_buf_2 _15048_ (.A(_08190_),
    .X(_09145_));
 sg13g2_buf_1 _15049_ (.A(net861),
    .X(_09146_));
 sg13g2_nand3_1 _15050_ (.B(\top_ihp.wb_dati_spi[0] ),
    .C(net841),
    .A(net918),
    .Y(_09147_));
 sg13g2_a21oi_1 _15051_ (.A1(_09142_),
    .A2(_09147_),
    .Y(_09148_),
    .B1(_08213_));
 sg13g2_a21oi_1 _15052_ (.A1(\top_ihp.wb_dati_rom[0] ),
    .A2(_08213_),
    .Y(_09149_),
    .B1(_09148_));
 sg13g2_nand2_1 _15053_ (.Y(_09150_),
    .A(_08216_),
    .B(\top_ihp.wb_dati_gpio[0] ));
 sg13g2_o21ai_1 _15054_ (.B1(_09150_),
    .Y(_09151_),
    .A1(_08216_),
    .A2(_09149_));
 sg13g2_buf_1 _15055_ (.A(_08215_),
    .X(_09152_));
 sg13g2_mux2_1 _15056_ (.A0(_09151_),
    .A1(\top_ihp.wb_dati_uart[0] ),
    .S(net992),
    .X(_09153_));
 sg13g2_a22oi_1 _15057_ (.Y(_09154_),
    .B1(_09153_),
    .B2(net954),
    .A2(_09140_),
    .A1(_09134_));
 sg13g2_or2_1 _15058_ (.X(_09155_),
    .B(_09154_),
    .A(_09127_));
 sg13g2_buf_1 _15059_ (.A(_09135_),
    .X(_09156_));
 sg13g2_buf_1 _15060_ (.A(net952),
    .X(_09157_));
 sg13g2_nor2_1 _15061_ (.A(_07822_),
    .B(net993),
    .Y(_09158_));
 sg13g2_nand2_1 _15062_ (.Y(_09159_),
    .A(_09125_),
    .B(_09158_));
 sg13g2_buf_2 _15063_ (.A(_09159_),
    .X(_09160_));
 sg13g2_buf_1 _15064_ (.A(net1018),
    .X(_09161_));
 sg13g2_nand2_1 _15065_ (.Y(_09162_),
    .A(_00072_),
    .B(_00071_));
 sg13g2_buf_1 _15066_ (.A(_09162_),
    .X(_09163_));
 sg13g2_buf_1 _15067_ (.A(net990),
    .X(_09164_));
 sg13g2_buf_1 _15068_ (.A(_08206_),
    .X(_09165_));
 sg13g2_buf_1 _15069_ (.A(net840),
    .X(_09166_));
 sg13g2_nor2_1 _15070_ (.A(\top_ihp.wb_dati_rom[24] ),
    .B(net821),
    .Y(_09167_));
 sg13g2_buf_1 _15071_ (.A(_08179_),
    .X(_09168_));
 sg13g2_buf_1 _15072_ (.A(net950),
    .X(_09169_));
 sg13g2_and3_1 _15073_ (.X(_09170_),
    .A(net918),
    .B(\top_ihp.wb_dati_spi[24] ),
    .C(net841));
 sg13g2_a221oi_1 _15074_ (.B2(\top_ihp.wb_dati_ram[24] ),
    .C1(_09170_),
    .B1(net872),
    .A1(_09169_),
    .Y(_09171_),
    .A2(net846));
 sg13g2_nor3_2 _15075_ (.A(net951),
    .B(_09167_),
    .C(_09171_),
    .Y(_09172_));
 sg13g2_nor2_1 _15076_ (.A(\top_ihp.wb_dati_rom[8] ),
    .B(net821),
    .Y(_09173_));
 sg13g2_buf_1 _15077_ (.A(net861),
    .X(_09174_));
 sg13g2_and3_1 _15078_ (.X(_09175_),
    .A(net918),
    .B(\top_ihp.wb_dati_spi[8] ),
    .C(net839));
 sg13g2_a221oi_1 _15079_ (.B2(\top_ihp.wb_dati_ram[8] ),
    .C1(_09175_),
    .B1(net872),
    .A1(net916),
    .Y(_09176_),
    .A2(net846));
 sg13g2_nor3_2 _15080_ (.A(net990),
    .B(_09173_),
    .C(_09176_),
    .Y(_09177_));
 sg13g2_and2_1 _15081_ (.A(net954),
    .B(_09177_),
    .X(_09178_));
 sg13g2_a21oi_1 _15082_ (.A1(_09161_),
    .A2(_09172_),
    .Y(_09179_),
    .B1(_09178_));
 sg13g2_buf_1 _15083_ (.A(_09057_),
    .X(_09180_));
 sg13g2_buf_1 _15084_ (.A(net915),
    .X(_09181_));
 sg13g2_nor2_1 _15085_ (.A(net998),
    .B(_08943_),
    .Y(_09182_));
 sg13g2_buf_1 _15086_ (.A(_09182_),
    .X(_09183_));
 sg13g2_nand2_1 _15087_ (.Y(_09184_),
    .A(_09121_),
    .B(_09183_));
 sg13g2_nor2_1 _15088_ (.A(net887),
    .B(_09184_),
    .Y(_09185_));
 sg13g2_o21ai_1 _15089_ (.B1(_09185_),
    .Y(_09186_),
    .A1(_09160_),
    .A2(_09179_));
 sg13g2_a21oi_1 _15090_ (.A1(net917),
    .A2(_09153_),
    .Y(_09187_),
    .B1(_09186_));
 sg13g2_buf_1 _15091_ (.A(_09183_),
    .X(_09188_));
 sg13g2_buf_1 _15092_ (.A(net1019),
    .X(_09189_));
 sg13g2_and2_1 _15093_ (.A(_07420_),
    .B(_08241_),
    .X(_09190_));
 sg13g2_buf_2 _15094_ (.A(_09190_),
    .X(_09191_));
 sg13g2_nor2_1 _15095_ (.A(net989),
    .B(_09191_),
    .Y(_09192_));
 sg13g2_nand3_1 _15096_ (.B(_07475_),
    .C(_09183_),
    .A(_07474_),
    .Y(_09193_));
 sg13g2_o21ai_1 _15097_ (.B1(_09193_),
    .Y(_09194_),
    .A1(_07474_),
    .A2(_07475_));
 sg13g2_nand2_1 _15098_ (.Y(_09195_),
    .A(_09192_),
    .B(_09194_));
 sg13g2_o21ai_1 _15099_ (.B1(_09195_),
    .Y(_09196_),
    .A1(_07475_),
    .A2(net886));
 sg13g2_a221oi_1 _15100_ (.B2(_09187_),
    .C1(_09196_),
    .B1(_09155_),
    .A1(_09120_),
    .Y(_09197_),
    .A2(_09124_));
 sg13g2_buf_1 _15101_ (.A(_09197_),
    .X(_09198_));
 sg13g2_buf_2 _15102_ (.A(_09198_),
    .X(_09199_));
 sg13g2_nand2_1 _15103_ (.Y(_09200_),
    .A(net412),
    .B(_09108_));
 sg13g2_o21ai_1 _15104_ (.B1(_09200_),
    .Y(_00358_),
    .A1(_09053_),
    .A2(_09108_));
 sg13g2_nand2b_1 _15105_ (.Y(_09201_),
    .B(_09106_),
    .A_N(_09082_));
 sg13g2_buf_1 _15106_ (.A(_09201_),
    .X(_09202_));
 sg13g2_buf_1 _15107_ (.A(_09202_),
    .X(_09203_));
 sg13g2_buf_1 _15108_ (.A(net550),
    .X(_09204_));
 sg13g2_buf_1 _15109_ (.A(_09188_),
    .X(_09205_));
 sg13g2_inv_1 _15110_ (.Y(_09206_),
    .A(\top_ihp.oisc.decoder.decoded[15] ));
 sg13g2_nor2_2 _15111_ (.A(_09109_),
    .B(_09206_),
    .Y(_09207_));
 sg13g2_o21ai_1 _15112_ (.B1(_09119_),
    .Y(_09208_),
    .A1(_09063_),
    .A2(_09207_));
 sg13g2_a21oi_1 _15113_ (.A1(_09115_),
    .A2(_09208_),
    .Y(_09209_),
    .B1(_09121_));
 sg13g2_buf_1 _15114_ (.A(_09209_),
    .X(_09210_));
 sg13g2_nor2_1 _15115_ (.A(\top_ihp.wb_dati_rom[23] ),
    .B(net862),
    .Y(_09211_));
 sg13g2_and2_1 _15116_ (.A(_08211_),
    .B(\top_ihp.wb_dati_spi[23] ),
    .X(_09212_));
 sg13g2_inv_1 _15117_ (.Y(_09213_),
    .A(\top_ihp.wb_dati_ram[23] ));
 sg13g2_nor4_1 _15118_ (.A(net981),
    .B(_09213_),
    .C(_08197_),
    .D(net903),
    .Y(_09214_));
 sg13g2_a221oi_1 _15119_ (.B2(_09212_),
    .C1(_09214_),
    .B1(net861),
    .A1(net950),
    .Y(_09215_),
    .A2(_07756_));
 sg13g2_or3_1 _15120_ (.A(net990),
    .B(_09211_),
    .C(_09215_),
    .X(_09216_));
 sg13g2_buf_1 _15121_ (.A(_09216_),
    .X(_09217_));
 sg13g2_nor2_1 _15122_ (.A(\top_ihp.wb_dati_rom[7] ),
    .B(net862),
    .Y(_09218_));
 sg13g2_and2_1 _15123_ (.A(net1012),
    .B(\top_ihp.wb_dati_spi[7] ),
    .X(_09219_));
 sg13g2_inv_1 _15124_ (.Y(_09220_),
    .A(\top_ihp.wb_dati_ram[7] ));
 sg13g2_buf_1 _15125_ (.A(_08197_),
    .X(_09221_));
 sg13g2_nor4_1 _15126_ (.A(net981),
    .B(_09220_),
    .C(net885),
    .D(net903),
    .Y(_09222_));
 sg13g2_a221oi_1 _15127_ (.B2(_09219_),
    .C1(_09222_),
    .B1(net861),
    .A1(net950),
    .Y(_09223_),
    .A2(_07756_));
 sg13g2_or3_1 _15128_ (.A(net980),
    .B(_09218_),
    .C(_09223_),
    .X(_09224_));
 sg13g2_buf_1 _15129_ (.A(_09224_),
    .X(_09225_));
 sg13g2_a21oi_1 _15130_ (.A1(_08215_),
    .A2(\top_ihp.wb_dati_uart[7] ),
    .Y(_09226_),
    .B1(_09136_));
 sg13g2_a22oi_1 _15131_ (.Y(_09227_),
    .B1(_09225_),
    .B2(_09226_),
    .A2(_09217_),
    .A1(_09136_));
 sg13g2_buf_2 _15132_ (.A(_09227_),
    .X(_09228_));
 sg13g2_nor2_1 _15133_ (.A(\top_ihp.wb_dati_rom[31] ),
    .B(_08205_),
    .Y(_09229_));
 sg13g2_and2_1 _15134_ (.A(_08191_),
    .B(\top_ihp.wb_dati_spi[31] ),
    .X(_09230_));
 sg13g2_inv_1 _15135_ (.Y(_09231_),
    .A(\top_ihp.wb_dati_ram[31] ));
 sg13g2_nor4_1 _15136_ (.A(_08194_),
    .B(_09231_),
    .C(_08197_),
    .D(_08199_),
    .Y(_09232_));
 sg13g2_a221oi_1 _15137_ (.B2(_09230_),
    .C1(_09232_),
    .B1(_08190_),
    .A1(_08179_),
    .Y(_09233_),
    .A2(net878));
 sg13g2_or3_1 _15138_ (.A(_09162_),
    .B(_09229_),
    .C(_09233_),
    .X(_09234_));
 sg13g2_buf_1 _15139_ (.A(_09234_),
    .X(_09235_));
 sg13g2_or3_1 _15140_ (.A(net1018),
    .B(_08203_),
    .C(_08209_),
    .X(_09236_));
 sg13g2_o21ai_1 _15141_ (.B1(_09236_),
    .Y(_09237_),
    .A1(_09137_),
    .A2(_09235_));
 sg13g2_buf_1 _15142_ (.A(_09237_),
    .X(_09238_));
 sg13g2_mux2_1 _15143_ (.A0(_09228_),
    .A1(_09238_),
    .S(_09125_),
    .X(_09239_));
 sg13g2_buf_1 _15144_ (.A(_07822_),
    .X(_09240_));
 sg13g2_buf_2 _15145_ (.A(\top_ihp.oisc.decoder.instruction[14] ),
    .X(_09241_));
 sg13g2_nor3_1 _15146_ (.A(_09240_),
    .B(net993),
    .C(_09241_),
    .Y(_09242_));
 sg13g2_a21oi_1 _15147_ (.A1(_09239_),
    .A2(_09242_),
    .Y(_09243_),
    .B1(_09180_));
 sg13g2_buf_2 _15148_ (.A(_09243_),
    .X(_09244_));
 sg13g2_buf_1 _15149_ (.A(_09135_),
    .X(_09245_));
 sg13g2_nor2_1 _15150_ (.A(\top_ihp.wb_dati_rom[10] ),
    .B(net862),
    .Y(_09246_));
 sg13g2_and2_1 _15151_ (.A(net1012),
    .B(\top_ihp.wb_dati_spi[10] ),
    .X(_09247_));
 sg13g2_buf_1 _15152_ (.A(net981),
    .X(_09248_));
 sg13g2_inv_1 _15153_ (.Y(_09249_),
    .A(\top_ihp.wb_dati_ram[10] ));
 sg13g2_buf_1 _15154_ (.A(net903),
    .X(_09250_));
 sg13g2_nor4_1 _15155_ (.A(net914),
    .B(_09249_),
    .C(net885),
    .D(net869),
    .Y(_09251_));
 sg13g2_a221oi_1 _15156_ (.B2(_09247_),
    .C1(_09251_),
    .B1(net839),
    .A1(net950),
    .Y(_09252_),
    .A2(net863));
 sg13g2_nor3_2 _15157_ (.A(net990),
    .B(_09246_),
    .C(_09252_),
    .Y(_09253_));
 sg13g2_nor2_1 _15158_ (.A(\top_ihp.wb_dati_rom[26] ),
    .B(net821),
    .Y(_09254_));
 sg13g2_and3_1 _15159_ (.X(_09255_),
    .A(net918),
    .B(\top_ihp.wb_dati_spi[26] ),
    .C(net839));
 sg13g2_a221oi_1 _15160_ (.B2(\top_ihp.wb_dati_ram[26] ),
    .C1(_09255_),
    .B1(net872),
    .A1(net916),
    .Y(_09256_),
    .A2(net846));
 sg13g2_nor3_2 _15161_ (.A(net951),
    .B(_09254_),
    .C(_09256_),
    .Y(_09257_));
 sg13g2_and2_1 _15162_ (.A(net954),
    .B(_09253_),
    .X(_09258_));
 sg13g2_a21o_1 _15163_ (.A2(_09257_),
    .A1(_09140_),
    .B1(_09258_),
    .X(_09259_));
 sg13g2_a22oi_1 _15164_ (.Y(_09260_),
    .B1(_09259_),
    .B2(net988),
    .A2(_09253_),
    .A1(net949));
 sg13g2_and2_1 _15165_ (.A(_07589_),
    .B(_07594_),
    .X(_09261_));
 sg13g2_o21ai_1 _15166_ (.B1(_09261_),
    .Y(_09262_),
    .A1(_07506_),
    .A2(_07555_));
 sg13g2_buf_1 _15167_ (.A(_09262_),
    .X(_09263_));
 sg13g2_xor2_1 _15168_ (.B(_09263_),
    .A(_07536_),
    .X(_09264_));
 sg13g2_a221oi_1 _15169_ (.B2(net887),
    .C1(net989),
    .B1(_09264_),
    .A1(_09244_),
    .Y(_09265_),
    .A2(_09260_));
 sg13g2_a21oi_1 _15170_ (.A1(\top_ihp.oisc.decoder.instruction[30] ),
    .A2(net870),
    .Y(_09266_),
    .B1(_09265_));
 sg13g2_nand2_1 _15171_ (.Y(_09267_),
    .A(net886),
    .B(_09266_));
 sg13g2_o21ai_1 _15172_ (.B1(_09267_),
    .Y(_09268_),
    .A1(_07534_),
    .A2(net871));
 sg13g2_buf_1 _15173_ (.A(_09268_),
    .X(_09269_));
 sg13g2_buf_2 _15174_ (.A(_09269_),
    .X(_09270_));
 sg13g2_buf_1 _15175_ (.A(_09202_),
    .X(_09271_));
 sg13g2_nand2_1 _15176_ (.Y(_09272_),
    .A(\top_ihp.oisc.regs[0][10] ),
    .B(net549));
 sg13g2_o21ai_1 _15177_ (.B1(_09272_),
    .Y(_00359_),
    .A1(net411),
    .A2(net74));
 sg13g2_nor2_1 _15178_ (.A(\top_ihp.wb_dati_rom[11] ),
    .B(net821),
    .Y(_09273_));
 sg13g2_buf_1 _15179_ (.A(_09169_),
    .X(_09274_));
 sg13g2_and3_1 _15180_ (.X(_09275_),
    .A(net918),
    .B(\top_ihp.wb_dati_spi[11] ),
    .C(net841));
 sg13g2_a221oi_1 _15181_ (.B2(\top_ihp.wb_dati_ram[11] ),
    .C1(_09275_),
    .B1(net872),
    .A1(net884),
    .Y(_09276_),
    .A2(net846));
 sg13g2_nor3_2 _15182_ (.A(_09164_),
    .B(_09273_),
    .C(_09276_),
    .Y(_09277_));
 sg13g2_inv_2 _15183_ (.Y(_09278_),
    .A(net993));
 sg13g2_nand2_1 _15184_ (.Y(_09279_),
    .A(_09278_),
    .B(net1018));
 sg13g2_nor2_1 _15185_ (.A(\top_ihp.wb_dati_rom[27] ),
    .B(net840),
    .Y(_09280_));
 sg13g2_nand2_1 _15186_ (.Y(_09281_),
    .A(\top_ihp.wb_dati_ram[27] ),
    .B(net872));
 sg13g2_nand3_1 _15187_ (.B(\top_ihp.wb_dati_spi[27] ),
    .C(net839),
    .A(net918),
    .Y(_09282_));
 sg13g2_nand3_1 _15188_ (.B(_09281_),
    .C(_09282_),
    .A(net821),
    .Y(_09283_));
 sg13g2_nand3b_1 _15189_ (.B(_09283_),
    .C(_08208_),
    .Y(_09284_),
    .A_N(_09280_));
 sg13g2_buf_1 _15190_ (.A(_09284_),
    .X(_09285_));
 sg13g2_nand2_1 _15191_ (.Y(_09286_),
    .A(net954),
    .B(_09277_));
 sg13g2_o21ai_1 _15192_ (.B1(_09286_),
    .Y(_09287_),
    .A1(_09279_),
    .A2(_09285_));
 sg13g2_a22oi_1 _15193_ (.Y(_09288_),
    .B1(_09287_),
    .B2(net988),
    .A2(_09277_),
    .A1(_09156_));
 sg13g2_and2_1 _15194_ (.A(_09244_),
    .B(_09288_),
    .X(_09289_));
 sg13g2_buf_1 _15195_ (.A(_09191_),
    .X(_09290_));
 sg13g2_a21oi_1 _15196_ (.A1(_07875_),
    .A2(_09263_),
    .Y(_09291_),
    .B1(_07568_));
 sg13g2_xor2_1 _15197_ (.B(_09291_),
    .A(_07533_),
    .X(_09292_));
 sg13g2_o21ai_1 _15198_ (.B1(net955),
    .Y(_09293_),
    .A1(net913),
    .A2(_09292_));
 sg13g2_buf_1 _15199_ (.A(net989),
    .X(_09294_));
 sg13g2_buf_1 _15200_ (.A(\top_ihp.oisc.decoder.instruction[31] ),
    .X(_09295_));
 sg13g2_nor2_1 _15201_ (.A(net995),
    .B(_09116_),
    .Y(_09296_));
 sg13g2_a22oi_1 _15202_ (.Y(_09297_),
    .B1(_09207_),
    .B2(_09296_),
    .A2(_09295_),
    .A1(net995));
 sg13g2_nand4_1 _15203_ (.B(_09114_),
    .C(net995),
    .A(net994),
    .Y(_09298_),
    .D(_09074_));
 sg13g2_o21ai_1 _15204_ (.B1(_09298_),
    .Y(_09299_),
    .A1(net994),
    .A2(_09297_));
 sg13g2_a21oi_1 _15205_ (.A1(net948),
    .A2(_09299_),
    .Y(_09300_),
    .B1(net873));
 sg13g2_o21ai_1 _15206_ (.B1(_09300_),
    .Y(_09301_),
    .A1(_09289_),
    .A2(_09293_));
 sg13g2_o21ai_1 _15207_ (.B1(_09301_),
    .Y(_09302_),
    .A1(_07531_),
    .A2(net871));
 sg13g2_buf_1 _15208_ (.A(_09302_),
    .X(_09303_));
 sg13g2_buf_1 _15209_ (.A(net251),
    .X(_09304_));
 sg13g2_buf_1 _15210_ (.A(_09202_),
    .X(_09305_));
 sg13g2_nand2_1 _15211_ (.Y(_09306_),
    .A(\top_ihp.oisc.regs[0][11] ),
    .B(net548));
 sg13g2_o21ai_1 _15212_ (.B1(_09306_),
    .Y(_00360_),
    .A1(net411),
    .A2(net148));
 sg13g2_buf_1 _15213_ (.A(_09123_),
    .X(_09307_));
 sg13g2_and3_1 _15214_ (.X(_09308_),
    .A(net994),
    .B(net996),
    .C(_09063_));
 sg13g2_buf_1 _15215_ (.A(_09308_),
    .X(_09309_));
 sg13g2_buf_1 _15216_ (.A(_09309_),
    .X(_09310_));
 sg13g2_nor3_2 _15217_ (.A(net994),
    .B(_09063_),
    .C(_09206_),
    .Y(_09311_));
 sg13g2_and2_1 _15218_ (.A(_09114_),
    .B(_09311_),
    .X(_09312_));
 sg13g2_buf_1 _15219_ (.A(_09312_),
    .X(_09313_));
 sg13g2_or2_1 _15220_ (.X(_09314_),
    .B(_09313_),
    .A(net883));
 sg13g2_buf_1 _15221_ (.A(_09314_),
    .X(_09315_));
 sg13g2_nand2_1 _15222_ (.Y(_09316_),
    .A(net994),
    .B(net996));
 sg13g2_nand3_1 _15223_ (.B(_09295_),
    .C(_09316_),
    .A(_09063_),
    .Y(_09317_));
 sg13g2_nand2_1 _15224_ (.Y(_09318_),
    .A(net989),
    .B(_09317_));
 sg13g2_buf_2 _15225_ (.A(_09318_),
    .X(_09319_));
 sg13g2_a21o_1 _15226_ (.A2(_09315_),
    .A1(net988),
    .B1(_09319_),
    .X(_09320_));
 sg13g2_buf_1 _15227_ (.A(net915),
    .X(_09321_));
 sg13g2_nor2_1 _15228_ (.A(_07531_),
    .B(_09291_),
    .Y(_09322_));
 sg13g2_nand2_1 _15229_ (.Y(_09323_),
    .A(_07531_),
    .B(_09291_));
 sg13g2_o21ai_1 _15230_ (.B1(_09323_),
    .Y(_09324_),
    .A1(_07532_),
    .A2(_09322_));
 sg13g2_xnor2_1 _15231_ (.Y(_09325_),
    .A(_07530_),
    .B(_09324_));
 sg13g2_nor2_1 _15232_ (.A(\top_ihp.wb_dati_rom[12] ),
    .B(net862),
    .Y(_09326_));
 sg13g2_and2_1 _15233_ (.A(\top_ihp.wb_dati_spi[12] ),
    .B(net1012),
    .X(_09327_));
 sg13g2_inv_1 _15234_ (.Y(_09328_),
    .A(\top_ihp.wb_dati_ram[12] ));
 sg13g2_nor4_1 _15235_ (.A(net914),
    .B(_09328_),
    .C(net885),
    .D(net903),
    .Y(_09329_));
 sg13g2_a221oi_1 _15236_ (.B2(_09327_),
    .C1(_09329_),
    .B1(net861),
    .A1(net950),
    .Y(_09330_),
    .A2(net863));
 sg13g2_nor3_1 _15237_ (.A(_09163_),
    .B(_09326_),
    .C(_09330_),
    .Y(_09331_));
 sg13g2_buf_1 _15238_ (.A(_09331_),
    .X(_09332_));
 sg13g2_nand2_1 _15239_ (.Y(_09333_),
    .A(net954),
    .B(net804));
 sg13g2_nor2_1 _15240_ (.A(\top_ihp.wb_dati_rom[28] ),
    .B(net840),
    .Y(_09334_));
 sg13g2_and2_1 _15241_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[28] ),
    .X(_09335_));
 sg13g2_inv_1 _15242_ (.Y(_09336_),
    .A(\top_ihp.wb_dati_ram[28] ));
 sg13g2_buf_1 _15243_ (.A(net885),
    .X(_09337_));
 sg13g2_nor4_1 _15244_ (.A(net914),
    .B(_09336_),
    .C(net868),
    .D(net869),
    .Y(_09338_));
 sg13g2_a221oi_1 _15245_ (.B2(_09335_),
    .C1(_09338_),
    .B1(net839),
    .A1(net916),
    .Y(_09339_),
    .A2(net863));
 sg13g2_nor3_2 _15246_ (.A(net990),
    .B(_09334_),
    .C(_09339_),
    .Y(_09340_));
 sg13g2_nand2_1 _15247_ (.Y(_09341_),
    .A(_09140_),
    .B(_09340_));
 sg13g2_nand2_1 _15248_ (.Y(_09342_),
    .A(_09333_),
    .B(_09341_));
 sg13g2_a22oi_1 _15249_ (.Y(_09343_),
    .B1(_09342_),
    .B2(net988),
    .A2(net804),
    .A1(net917));
 sg13g2_nand2_1 _15250_ (.Y(_09344_),
    .A(_09183_),
    .B(_09320_));
 sg13g2_a221oi_1 _15251_ (.B2(_09244_),
    .C1(_09344_),
    .B1(_09343_),
    .A1(_09321_),
    .Y(_09345_),
    .A2(_09325_));
 sg13g2_a221oi_1 _15252_ (.B2(_09320_),
    .C1(_09345_),
    .B1(_09124_),
    .A1(_07528_),
    .Y(_09346_),
    .A2(net860));
 sg13g2_buf_2 _15253_ (.A(_09346_),
    .X(_09347_));
 sg13g2_buf_1 _15254_ (.A(_09347_),
    .X(_09348_));
 sg13g2_nand2_1 _15255_ (.Y(_09349_),
    .A(\top_ihp.oisc.regs[0][12] ),
    .B(net548));
 sg13g2_o21ai_1 _15256_ (.B1(_09349_),
    .Y(_00361_),
    .A1(net411),
    .A2(net250));
 sg13g2_buf_1 _15257_ (.A(_09077_),
    .X(_09350_));
 sg13g2_buf_1 _15258_ (.A(net867),
    .X(_09351_));
 sg13g2_nor2_1 _15259_ (.A(\top_ihp.wb_dati_rom[13] ),
    .B(net862),
    .Y(_09352_));
 sg13g2_and2_1 _15260_ (.A(net1012),
    .B(\top_ihp.wb_dati_spi[13] ),
    .X(_09353_));
 sg13g2_inv_1 _15261_ (.Y(_09354_),
    .A(\top_ihp.wb_dati_ram[13] ));
 sg13g2_nor4_1 _15262_ (.A(net914),
    .B(_09354_),
    .C(net885),
    .D(net903),
    .Y(_09355_));
 sg13g2_a221oi_1 _15263_ (.B2(_09353_),
    .C1(_09355_),
    .B1(net861),
    .A1(net950),
    .Y(_09356_),
    .A2(net863));
 sg13g2_nor3_1 _15264_ (.A(net951),
    .B(_09352_),
    .C(_09356_),
    .Y(_09357_));
 sg13g2_nor2_1 _15265_ (.A(\top_ihp.wb_dati_rom[29] ),
    .B(net821),
    .Y(_09358_));
 sg13g2_and3_1 _15266_ (.X(_09359_),
    .A(net918),
    .B(\top_ihp.wb_dati_spi[29] ),
    .C(net841));
 sg13g2_a221oi_1 _15267_ (.B2(\top_ihp.wb_dati_ram[29] ),
    .C1(_09359_),
    .B1(net872),
    .A1(net884),
    .Y(_09360_),
    .A2(net846));
 sg13g2_nor3_2 _15268_ (.A(net951),
    .B(_09358_),
    .C(_09360_),
    .Y(_09361_));
 sg13g2_or3_1 _15269_ (.A(net990),
    .B(_09352_),
    .C(_09356_),
    .X(_09362_));
 sg13g2_buf_1 _15270_ (.A(_09362_),
    .X(_09363_));
 sg13g2_nor2_1 _15271_ (.A(net1018),
    .B(_09363_),
    .Y(_09364_));
 sg13g2_a21o_1 _15272_ (.A2(_09361_),
    .A1(net991),
    .B1(_09364_),
    .X(_09365_));
 sg13g2_nor2b_1 _15273_ (.A(net993),
    .B_N(net988),
    .Y(_09366_));
 sg13g2_a22oi_1 _15274_ (.Y(_09367_),
    .B1(_09365_),
    .B2(_09366_),
    .A2(_09357_),
    .A1(net949));
 sg13g2_xnor2_1 _15275_ (.Y(_09368_),
    .A(_07527_),
    .B(_07884_));
 sg13g2_a22oi_1 _15276_ (.Y(_09369_),
    .B1(_09368_),
    .B2(_09181_),
    .A2(_09367_),
    .A1(_09244_));
 sg13g2_nor2_1 _15277_ (.A(net948),
    .B(_09369_),
    .Y(_09370_));
 sg13g2_a21oi_1 _15278_ (.A1(net917),
    .A2(_09315_),
    .Y(_09371_),
    .B1(_09319_));
 sg13g2_nor3_1 _15279_ (.A(net860),
    .B(_09370_),
    .C(_09371_),
    .Y(_09372_));
 sg13g2_a21oi_1 _15280_ (.A1(net1034),
    .A2(net859),
    .Y(_09373_),
    .B1(_09372_));
 sg13g2_buf_1 _15281_ (.A(_09373_),
    .X(_09374_));
 sg13g2_buf_8 _15282_ (.A(net147),
    .X(_09375_));
 sg13g2_nand2_1 _15283_ (.Y(_09376_),
    .A(\top_ihp.oisc.regs[0][13] ),
    .B(_09305_));
 sg13g2_o21ai_1 _15284_ (.B1(_09376_),
    .Y(_00362_),
    .A1(net411),
    .A2(net73));
 sg13g2_nor2_1 _15285_ (.A(\top_ihp.wb_dati_rom[14] ),
    .B(net840),
    .Y(_09377_));
 sg13g2_and2_1 _15286_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[14] ),
    .X(_09378_));
 sg13g2_inv_1 _15287_ (.Y(_09379_),
    .A(\top_ihp.wb_dati_ram[14] ));
 sg13g2_nor4_1 _15288_ (.A(net914),
    .B(_09379_),
    .C(net885),
    .D(net869),
    .Y(_09380_));
 sg13g2_a221oi_1 _15289_ (.B2(_09378_),
    .C1(_09380_),
    .B1(net839),
    .A1(net916),
    .Y(_09381_),
    .A2(net863));
 sg13g2_nor3_1 _15290_ (.A(net951),
    .B(_09377_),
    .C(_09381_),
    .Y(_09382_));
 sg13g2_buf_2 _15291_ (.A(_09382_),
    .X(_09383_));
 sg13g2_nor2_1 _15292_ (.A(\top_ihp.wb_dati_rom[30] ),
    .B(net821),
    .Y(_09384_));
 sg13g2_and2_1 _15293_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[30] ),
    .X(_09385_));
 sg13g2_inv_1 _15294_ (.Y(_09386_),
    .A(\top_ihp.wb_dati_ram[30] ));
 sg13g2_nor4_1 _15295_ (.A(net914),
    .B(_09386_),
    .C(net868),
    .D(net869),
    .Y(_09387_));
 sg13g2_a221oi_1 _15296_ (.B2(_09385_),
    .C1(_09387_),
    .B1(net841),
    .A1(net916),
    .Y(_09388_),
    .A2(net846));
 sg13g2_nor3_2 _15297_ (.A(_09164_),
    .B(_09384_),
    .C(_09388_),
    .Y(_09389_));
 sg13g2_or3_1 _15298_ (.A(_09163_),
    .B(_09377_),
    .C(_09381_),
    .X(_09390_));
 sg13g2_buf_2 _15299_ (.A(_09390_),
    .X(_09391_));
 sg13g2_nor2_1 _15300_ (.A(net991),
    .B(_09391_),
    .Y(_09392_));
 sg13g2_a21oi_1 _15301_ (.A1(net991),
    .A2(_09389_),
    .Y(_09393_),
    .B1(_09392_));
 sg13g2_nor2b_1 _15302_ (.A(_09393_),
    .B_N(_09366_),
    .Y(_09394_));
 sg13g2_a21oi_1 _15303_ (.A1(net917),
    .A2(_09383_),
    .Y(_09395_),
    .B1(_09394_));
 sg13g2_a22oi_1 _15304_ (.Y(_09396_),
    .B1(_09263_),
    .B2(_07537_),
    .A2(_07578_),
    .A1(_07575_));
 sg13g2_xnor2_1 _15305_ (.Y(_09397_),
    .A(_07523_),
    .B(_09396_));
 sg13g2_a22oi_1 _15306_ (.Y(_09398_),
    .B1(_09397_),
    .B2(net882),
    .A2(_09395_),
    .A1(_09244_));
 sg13g2_a221oi_1 _15307_ (.B2(_07829_),
    .C1(_09319_),
    .B1(_09313_),
    .A1(_09241_),
    .Y(_09399_),
    .A2(net883));
 sg13g2_nor2_1 _15308_ (.A(_07521_),
    .B(net886),
    .Y(_09400_));
 sg13g2_a21oi_1 _15309_ (.A1(net886),
    .A2(_09399_),
    .Y(_09401_),
    .B1(_09400_));
 sg13g2_o21ai_1 _15310_ (.B1(_09401_),
    .Y(_09402_),
    .A1(_09184_),
    .A2(_09398_));
 sg13g2_buf_1 _15311_ (.A(_09402_),
    .X(_09403_));
 sg13g2_buf_2 _15312_ (.A(_09403_),
    .X(_09404_));
 sg13g2_nand2_1 _15313_ (.Y(_09405_),
    .A(\top_ihp.oisc.regs[0][14] ),
    .B(net548));
 sg13g2_o21ai_1 _15314_ (.B1(_09405_),
    .Y(_00363_),
    .A1(net411),
    .A2(net249));
 sg13g2_nor2_1 _15315_ (.A(_08203_),
    .B(_08209_),
    .Y(_09406_));
 sg13g2_a22oi_1 _15316_ (.Y(_09407_),
    .B1(_09238_),
    .B2(_09366_),
    .A2(_09406_),
    .A1(net917));
 sg13g2_inv_1 _15317_ (.Y(_09408_),
    .A(_07885_));
 sg13g2_o21ai_1 _15318_ (.B1(_07901_),
    .Y(_09409_),
    .A1(_07884_),
    .A2(_09408_));
 sg13g2_buf_1 _15319_ (.A(_09409_),
    .X(_09410_));
 sg13g2_xnor2_1 _15320_ (.Y(_09411_),
    .A(_07511_),
    .B(_09410_));
 sg13g2_xnor2_1 _15321_ (.Y(_09412_),
    .A(net1036),
    .B(_09411_));
 sg13g2_a22oi_1 _15322_ (.Y(_09413_),
    .B1(_09412_),
    .B2(net882),
    .A2(_09407_),
    .A1(_09244_));
 sg13g2_a21oi_1 _15323_ (.A1(\top_ihp.oisc.decoder.instruction[15] ),
    .A2(_09315_),
    .Y(_09414_),
    .B1(_09319_));
 sg13g2_nand2_1 _15324_ (.Y(_09415_),
    .A(net1036),
    .B(net873));
 sg13g2_o21ai_1 _15325_ (.B1(_09415_),
    .Y(_09416_),
    .A1(net867),
    .A2(_09414_));
 sg13g2_o21ai_1 _15326_ (.B1(_09416_),
    .Y(_09417_),
    .A1(_09184_),
    .A2(_09413_));
 sg13g2_buf_2 _15327_ (.A(_09417_),
    .X(_09418_));
 sg13g2_buf_1 _15328_ (.A(_09418_),
    .X(_09419_));
 sg13g2_nand2_1 _15329_ (.Y(_09420_),
    .A(\top_ihp.oisc.regs[0][15] ),
    .B(net548));
 sg13g2_o21ai_1 _15330_ (.B1(_09420_),
    .Y(_00364_),
    .A1(net411),
    .A2(net248));
 sg13g2_inv_1 _15331_ (.Y(_09421_),
    .A(_00103_));
 sg13g2_a221oi_1 _15332_ (.B2(_09421_),
    .C1(_09319_),
    .B1(_09313_),
    .A1(\top_ihp.oisc.decoder.instruction[16] ),
    .Y(_09422_),
    .A2(net883));
 sg13g2_o21ai_1 _15333_ (.B1(_07513_),
    .Y(_09423_),
    .A1(_07904_),
    .A2(_09410_));
 sg13g2_xnor2_1 _15334_ (.Y(_09424_),
    .A(_07509_),
    .B(_09423_));
 sg13g2_nor4_1 _15335_ (.A(_07822_),
    .B(_09125_),
    .C(_09241_),
    .D(_09057_),
    .Y(_09425_));
 sg13g2_nor2_1 _15336_ (.A(_07822_),
    .B(_09125_),
    .Y(_09426_));
 sg13g2_nor3_1 _15337_ (.A(_09241_),
    .B(_09057_),
    .C(_09426_),
    .Y(_09427_));
 sg13g2_nor2_1 _15338_ (.A(_09278_),
    .B(_09057_),
    .Y(_09428_));
 sg13g2_a221oi_1 _15339_ (.B2(_09238_),
    .C1(_09428_),
    .B1(_09427_),
    .A1(_09228_),
    .Y(_09429_),
    .A2(_09425_));
 sg13g2_buf_1 _15340_ (.A(_09429_),
    .X(_09430_));
 sg13g2_nor2_1 _15341_ (.A(_09278_),
    .B(_09134_),
    .Y(_09431_));
 sg13g2_o21ai_1 _15342_ (.B1(net955),
    .Y(_09432_),
    .A1(_09430_),
    .A2(_09431_));
 sg13g2_a21oi_1 _15343_ (.A1(net882),
    .A2(_09424_),
    .Y(_09433_),
    .B1(_09432_));
 sg13g2_nor3_1 _15344_ (.A(_09350_),
    .B(_09422_),
    .C(_09433_),
    .Y(_09434_));
 sg13g2_a21oi_1 _15345_ (.A1(_07507_),
    .A2(net859),
    .Y(_09435_),
    .B1(_09434_));
 sg13g2_buf_2 _15346_ (.A(_09435_),
    .X(_09436_));
 sg13g2_buf_8 _15347_ (.A(net247),
    .X(_09437_));
 sg13g2_nand2_1 _15348_ (.Y(_09438_),
    .A(\top_ihp.oisc.regs[0][16] ),
    .B(net548));
 sg13g2_o21ai_1 _15349_ (.B1(_09438_),
    .Y(_00365_),
    .A1(_09204_),
    .A2(net146));
 sg13g2_nor3_1 _15350_ (.A(net993),
    .B(_09241_),
    .C(_09426_),
    .Y(_09439_));
 sg13g2_nor4_1 _15351_ (.A(_07822_),
    .B(_07823_),
    .C(_09125_),
    .D(_09241_),
    .Y(_09440_));
 sg13g2_a22oi_1 _15352_ (.Y(_09441_),
    .B1(_09440_),
    .B2(_09228_),
    .A2(_09439_),
    .A1(_09238_));
 sg13g2_buf_8 _15353_ (.A(_09441_),
    .X(_09442_));
 sg13g2_inv_4 _15354_ (.A(_09442_),
    .Y(_09443_));
 sg13g2_and2_1 _15355_ (.A(_08191_),
    .B(\top_ihp.wb_dati_spi[17] ),
    .X(_09444_));
 sg13g2_inv_1 _15356_ (.Y(_09445_),
    .A(\top_ihp.wb_dati_ram[17] ));
 sg13g2_nor4_1 _15357_ (.A(net981),
    .B(_09445_),
    .C(_08197_),
    .D(_08199_),
    .Y(_09446_));
 sg13g2_a221oi_1 _15358_ (.B2(_09444_),
    .C1(_09446_),
    .B1(_08190_),
    .A1(_08179_),
    .Y(_09447_),
    .A2(net878));
 sg13g2_buf_1 _15359_ (.A(_09447_),
    .X(_09448_));
 sg13g2_o21ai_1 _15360_ (.B1(_09132_),
    .Y(_09449_),
    .A1(\top_ihp.wb_dati_rom[17] ),
    .A2(_08205_));
 sg13g2_nor3_1 _15361_ (.A(_09278_),
    .B(_09448_),
    .C(_09449_),
    .Y(_09450_));
 sg13g2_nor2_1 _15362_ (.A(_09443_),
    .B(_09450_),
    .Y(_09451_));
 sg13g2_a22oi_1 _15363_ (.Y(_09452_),
    .B1(_09410_),
    .B2(_07515_),
    .A2(_07907_),
    .A1(_07903_));
 sg13g2_xnor2_1 _15364_ (.Y(_09453_),
    .A(_07886_),
    .B(_09452_));
 sg13g2_nor2_1 _15365_ (.A(net913),
    .B(_09453_),
    .Y(_09454_));
 sg13g2_a21oi_1 _15366_ (.A1(net913),
    .A2(_09451_),
    .Y(_09455_),
    .B1(_09454_));
 sg13g2_inv_1 _15367_ (.Y(_09456_),
    .A(_00104_));
 sg13g2_a221oi_1 _15368_ (.B2(_09456_),
    .C1(_09319_),
    .B1(_09313_),
    .A1(\top_ihp.oisc.decoder.instruction[17] ),
    .Y(_09457_),
    .A2(net883));
 sg13g2_nand2_1 _15369_ (.Y(_09458_),
    .A(net1035),
    .B(net873));
 sg13g2_o21ai_1 _15370_ (.B1(_09458_),
    .Y(_09459_),
    .A1(net867),
    .A2(_09457_));
 sg13g2_o21ai_1 _15371_ (.B1(_09459_),
    .Y(_09460_),
    .A1(_09184_),
    .A2(_09455_));
 sg13g2_buf_1 _15372_ (.A(_09460_),
    .X(_09461_));
 sg13g2_buf_1 _15373_ (.A(_09461_),
    .X(_09462_));
 sg13g2_nand2_1 _15374_ (.Y(_09463_),
    .A(\top_ihp.oisc.regs[0][17] ),
    .B(net548));
 sg13g2_o21ai_1 _15375_ (.B1(_09463_),
    .Y(_00366_),
    .A1(net411),
    .A2(net145));
 sg13g2_nand2b_1 _15376_ (.Y(_09464_),
    .B(_07556_),
    .A_N(_07506_));
 sg13g2_nor4_2 _15377_ (.A(_07520_),
    .B(_07565_),
    .C(_07579_),
    .Y(_09465_),
    .D(_07595_));
 sg13g2_nand2_1 _15378_ (.Y(_09466_),
    .A(_09464_),
    .B(_09465_));
 sg13g2_xnor2_1 _15379_ (.Y(_09467_),
    .A(_07608_),
    .B(_09466_));
 sg13g2_and2_1 _15380_ (.A(_08191_),
    .B(\top_ihp.wb_dati_spi[18] ),
    .X(_09468_));
 sg13g2_inv_1 _15381_ (.Y(_09469_),
    .A(\top_ihp.wb_dati_ram[18] ));
 sg13g2_nor4_1 _15382_ (.A(net981),
    .B(_09469_),
    .C(_08197_),
    .D(_08200_),
    .Y(_09470_));
 sg13g2_a221oi_1 _15383_ (.B2(_09468_),
    .C1(_09470_),
    .B1(_09145_),
    .A1(net950),
    .Y(_09471_),
    .A2(net878));
 sg13g2_o21ai_1 _15384_ (.B1(_09132_),
    .Y(_09472_),
    .A1(\top_ihp.wb_dati_rom[18] ),
    .A2(_08205_));
 sg13g2_nor2_1 _15385_ (.A(_09471_),
    .B(_09472_),
    .Y(_09473_));
 sg13g2_nand2_1 _15386_ (.Y(_09474_),
    .A(_09156_),
    .B(_09473_));
 sg13g2_nand3_1 _15387_ (.B(_09442_),
    .C(_09474_),
    .A(_09290_),
    .Y(_09475_));
 sg13g2_o21ai_1 _15388_ (.B1(_09475_),
    .Y(_09476_),
    .A1(net913),
    .A2(_09467_));
 sg13g2_nand2_1 _15389_ (.Y(_09477_),
    .A(net955),
    .B(_09476_));
 sg13g2_a21oi_1 _15390_ (.A1(\top_ihp.oisc.decoder.instruction[18] ),
    .A2(net883),
    .Y(_09478_),
    .B1(_09319_));
 sg13g2_nand2b_1 _15391_ (.Y(_09479_),
    .B(_09313_),
    .A_N(_00105_));
 sg13g2_a21oi_1 _15392_ (.A1(_09478_),
    .A2(_09479_),
    .Y(_09480_),
    .B1(net860));
 sg13g2_a22oi_1 _15393_ (.Y(_09481_),
    .B1(_09477_),
    .B2(_09480_),
    .A2(net859),
    .A1(net1043));
 sg13g2_buf_1 _15394_ (.A(_09481_),
    .X(_09482_));
 sg13g2_buf_1 _15395_ (.A(_09482_),
    .X(_09483_));
 sg13g2_nand2_1 _15396_ (.Y(_09484_),
    .A(\top_ihp.oisc.regs[0][18] ),
    .B(net548));
 sg13g2_o21ai_1 _15397_ (.B1(_09484_),
    .Y(_00367_),
    .A1(net411),
    .A2(net144));
 sg13g2_or3_1 _15398_ (.A(_07897_),
    .B(_09408_),
    .C(_07887_),
    .X(_09485_));
 sg13g2_nor2_1 _15399_ (.A(net1043),
    .B(_07890_),
    .Y(_09486_));
 sg13g2_nand3_1 _15400_ (.B(_07903_),
    .C(_07907_),
    .A(_07516_),
    .Y(_09487_));
 sg13g2_a21oi_1 _15401_ (.A1(_07903_),
    .A2(_07907_),
    .Y(_09488_),
    .B1(_07516_));
 sg13g2_a221oi_1 _15402_ (.B2(_09487_),
    .C1(_09488_),
    .B1(net1035),
    .A1(net1043),
    .Y(_09489_),
    .A2(_07890_));
 sg13g2_nor3_1 _15403_ (.A(_07897_),
    .B(_07887_),
    .C(_07901_),
    .Y(_09490_));
 sg13g2_nor3_1 _15404_ (.A(_09486_),
    .B(_09489_),
    .C(_09490_),
    .Y(_09491_));
 sg13g2_o21ai_1 _15405_ (.B1(_09491_),
    .Y(_09492_),
    .A1(_07884_),
    .A2(_09485_));
 sg13g2_buf_1 _15406_ (.A(_09492_),
    .X(_09493_));
 sg13g2_xnor2_1 _15407_ (.Y(_09494_),
    .A(_07604_),
    .B(_09493_));
 sg13g2_and2_1 _15408_ (.A(net1012),
    .B(\top_ihp.wb_dati_spi[19] ),
    .X(_09495_));
 sg13g2_inv_1 _15409_ (.Y(_09496_),
    .A(\top_ihp.wb_dati_ram[19] ));
 sg13g2_nor4_1 _15410_ (.A(net981),
    .B(_09496_),
    .C(_09221_),
    .D(_08200_),
    .Y(_09497_));
 sg13g2_a221oi_1 _15411_ (.B2(_09495_),
    .C1(_09497_),
    .B1(_09145_),
    .A1(_09168_),
    .Y(_09498_),
    .A2(net878));
 sg13g2_buf_1 _15412_ (.A(_09498_),
    .X(_09499_));
 sg13g2_o21ai_1 _15413_ (.B1(_09132_),
    .Y(_09500_),
    .A1(\top_ihp.wb_dati_rom[19] ),
    .A2(_08206_));
 sg13g2_buf_1 _15414_ (.A(_09500_),
    .X(_09501_));
 sg13g2_nor2_1 _15415_ (.A(_09499_),
    .B(_09501_),
    .Y(_09502_));
 sg13g2_nor2_1 _15416_ (.A(_09278_),
    .B(_09502_),
    .Y(_09503_));
 sg13g2_o21ai_1 _15417_ (.B1(_09078_),
    .Y(_09504_),
    .A1(_09430_),
    .A2(_09503_));
 sg13g2_a21oi_1 _15418_ (.A1(net882),
    .A2(_09494_),
    .Y(_09505_),
    .B1(_09504_));
 sg13g2_inv_1 _15419_ (.Y(_09506_),
    .A(_00106_));
 sg13g2_a221oi_1 _15420_ (.B2(_09506_),
    .C1(_09319_),
    .B1(_09313_),
    .A1(\top_ihp.oisc.decoder.instruction[19] ),
    .Y(_09507_),
    .A2(net883));
 sg13g2_nand2_1 _15421_ (.Y(_09508_),
    .A(net1042),
    .B(net873));
 sg13g2_o21ai_1 _15422_ (.B1(_09508_),
    .Y(_09509_),
    .A1(net867),
    .A2(_09507_));
 sg13g2_nand2b_1 _15423_ (.Y(_09510_),
    .B(_09509_),
    .A_N(_09505_));
 sg13g2_buf_1 _15424_ (.A(_09510_),
    .X(_09511_));
 sg13g2_buf_2 _15425_ (.A(_09511_),
    .X(_09512_));
 sg13g2_nand2_1 _15426_ (.Y(_09513_),
    .A(\top_ihp.oisc.regs[0][19] ),
    .B(_09305_));
 sg13g2_o21ai_1 _15427_ (.B1(_09513_),
    .Y(_00368_),
    .A1(_09204_),
    .A2(net246));
 sg13g2_buf_1 _15428_ (.A(_09203_),
    .X(_09514_));
 sg13g2_nor2_1 _15429_ (.A(\top_ihp.wb_dati_rom[25] ),
    .B(net840),
    .Y(_09515_));
 sg13g2_and2_1 _15430_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[25] ),
    .X(_09516_));
 sg13g2_inv_1 _15431_ (.Y(_09517_),
    .A(\top_ihp.wb_dati_ram[25] ));
 sg13g2_nor4_1 _15432_ (.A(net914),
    .B(_09517_),
    .C(_09337_),
    .D(net869),
    .Y(_09518_));
 sg13g2_a221oi_1 _15433_ (.B2(_09516_),
    .C1(_09518_),
    .B1(net841),
    .A1(net916),
    .Y(_09519_),
    .A2(net863));
 sg13g2_nor3_2 _15434_ (.A(net990),
    .B(_09515_),
    .C(_09519_),
    .Y(_09520_));
 sg13g2_nor3_1 _15435_ (.A(_09127_),
    .B(_09448_),
    .C(_09449_),
    .Y(_09521_));
 sg13g2_a21oi_1 _15436_ (.A1(_09127_),
    .A2(_09520_),
    .Y(_09522_),
    .B1(_09521_));
 sg13g2_and2_1 _15437_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[9] ),
    .X(_09523_));
 sg13g2_mux2_1 _15438_ (.A0(\top_ihp.wb_dati_ram[9] ),
    .A1(_09523_),
    .S(_09174_),
    .X(_09524_));
 sg13g2_mux2_1 _15439_ (.A0(\top_ihp.wb_dati_rom[9] ),
    .A1(_09524_),
    .S(net840),
    .X(_09525_));
 sg13g2_nand2_2 _15440_ (.Y(_09526_),
    .A(_08208_),
    .B(_09525_));
 sg13g2_nand2b_1 _15441_ (.Y(_09527_),
    .B(_09125_),
    .A_N(_07822_));
 sg13g2_buf_1 _15442_ (.A(_09527_),
    .X(_09528_));
 sg13g2_nor2_1 _15443_ (.A(net991),
    .B(_09528_),
    .Y(_09529_));
 sg13g2_a22oi_1 _15444_ (.Y(_09530_),
    .B1(_09526_),
    .B2(_09529_),
    .A2(_09522_),
    .A1(net991));
 sg13g2_nand2_1 _15445_ (.Y(_09531_),
    .A(\top_ihp.wb_dati_ram[1] ),
    .B(_09141_));
 sg13g2_nand3_1 _15446_ (.B(\top_ihp.wb_dati_spi[1] ),
    .C(_09146_),
    .A(_09144_),
    .Y(_09532_));
 sg13g2_a21oi_1 _15447_ (.A1(_09531_),
    .A2(_09532_),
    .Y(_09533_),
    .B1(_08213_));
 sg13g2_a21oi_1 _15448_ (.A1(\top_ihp.wb_dati_rom[1] ),
    .A2(_08213_),
    .Y(_09534_),
    .B1(_09533_));
 sg13g2_nand2_1 _15449_ (.Y(_09535_),
    .A(net954),
    .B(_09528_));
 sg13g2_a22oi_1 _15450_ (.Y(_09536_),
    .B1(_09535_),
    .B2(_09278_),
    .A2(\top_ihp.wb_dati_uart[1] ),
    .A1(net992));
 sg13g2_o21ai_1 _15451_ (.B1(_09536_),
    .Y(_09537_),
    .A1(net980),
    .A2(_09534_));
 sg13g2_o21ai_1 _15452_ (.B1(_09537_),
    .Y(_09538_),
    .A1(net917),
    .A2(_09530_));
 sg13g2_xnor2_1 _15453_ (.Y(_09539_),
    .A(net1041),
    .B(_08174_));
 sg13g2_a21oi_1 _15454_ (.A1(_09321_),
    .A2(_09539_),
    .Y(_09540_),
    .B1(net948));
 sg13g2_o21ai_1 _15455_ (.B1(_09540_),
    .Y(_09541_),
    .A1(net882),
    .A2(_09538_));
 sg13g2_buf_1 _15456_ (.A(\top_ihp.oisc.decoder.instruction[21] ),
    .X(_09542_));
 sg13g2_nand2_1 _15457_ (.Y(_09543_),
    .A(net956),
    .B(_09542_));
 sg13g2_o21ai_1 _15458_ (.B1(_09543_),
    .Y(_09544_),
    .A1(net956),
    .A2(_00099_));
 sg13g2_a21oi_1 _15459_ (.A1(_09311_),
    .A2(_09544_),
    .Y(_09545_),
    .B1(_09122_));
 sg13g2_nor2_1 _15460_ (.A(_09119_),
    .B(net996),
    .Y(_09546_));
 sg13g2_mux2_1 _15461_ (.A0(_09542_),
    .A1(_09055_),
    .S(net956),
    .X(_09547_));
 sg13g2_a22oi_1 _15462_ (.Y(_09548_),
    .B1(_09547_),
    .B2(_09119_),
    .A2(_09546_),
    .A1(_09055_));
 sg13g2_nand2b_1 _15463_ (.Y(_09549_),
    .B(net995),
    .A_N(_09548_));
 sg13g2_a21oi_1 _15464_ (.A1(_09545_),
    .A2(_09549_),
    .Y(_09550_),
    .B1(net860));
 sg13g2_a22oi_1 _15465_ (.Y(_09551_),
    .B1(_09541_),
    .B2(_09550_),
    .A2(net859),
    .A1(net1041));
 sg13g2_buf_1 _15466_ (.A(_09551_),
    .X(_09552_));
 sg13g2_buf_2 _15467_ (.A(_09552_),
    .X(_09553_));
 sg13g2_buf_1 _15468_ (.A(net547),
    .X(_09554_));
 sg13g2_nand2_1 _15469_ (.Y(_09555_),
    .A(\top_ihp.oisc.regs[0][1] ),
    .B(net548));
 sg13g2_o21ai_1 _15470_ (.B1(_09555_),
    .Y(_00369_),
    .A1(net410),
    .A2(net409));
 sg13g2_nor2_1 _15471_ (.A(_07450_),
    .B(_09183_),
    .Y(_09556_));
 sg13g2_inv_1 _15472_ (.Y(_09557_),
    .A(net1042));
 sg13g2_nand2_1 _15473_ (.Y(_09558_),
    .A(_09557_),
    .B(_09493_));
 sg13g2_o21ai_1 _15474_ (.B1(_07453_),
    .Y(_09559_),
    .A1(_09557_),
    .A2(_09493_));
 sg13g2_and3_1 _15475_ (.X(_09560_),
    .A(_07605_),
    .B(_09558_),
    .C(_09559_));
 sg13g2_a21oi_1 _15476_ (.A1(_09558_),
    .A2(_09559_),
    .Y(_09561_),
    .B1(_07605_));
 sg13g2_nor3_1 _15477_ (.A(_09191_),
    .B(_09560_),
    .C(_09561_),
    .Y(_09562_));
 sg13g2_buf_2 _15478_ (.A(_09562_),
    .X(_09563_));
 sg13g2_nor2_1 _15479_ (.A(\top_ihp.wb_dati_rom[20] ),
    .B(net840),
    .Y(_09564_));
 sg13g2_and2_1 _15480_ (.A(_09143_),
    .B(\top_ihp.wb_dati_spi[20] ),
    .X(_09565_));
 sg13g2_inv_1 _15481_ (.Y(_09566_),
    .A(\top_ihp.wb_dati_ram[20] ));
 sg13g2_nor4_1 _15482_ (.A(_09248_),
    .B(_09566_),
    .C(net868),
    .D(_09250_),
    .Y(_09567_));
 sg13g2_a221oi_1 _15483_ (.B2(_09565_),
    .C1(_09567_),
    .B1(net841),
    .A1(net916),
    .Y(_09568_),
    .A2(_07757_));
 sg13g2_nor3_2 _15484_ (.A(net990),
    .B(_09564_),
    .C(_09568_),
    .Y(_09569_));
 sg13g2_a21oi_1 _15485_ (.A1(net949),
    .A2(_09569_),
    .Y(_09570_),
    .B1(_09443_));
 sg13g2_and2_1 _15486_ (.A(_09191_),
    .B(_09570_),
    .X(_09571_));
 sg13g2_nor4_1 _15487_ (.A(net989),
    .B(_09556_),
    .C(_09563_),
    .D(_09571_),
    .Y(_09572_));
 sg13g2_buf_1 _15488_ (.A(_09572_),
    .X(_09573_));
 sg13g2_and2_1 _15489_ (.A(net1019),
    .B(_09309_),
    .X(_09574_));
 sg13g2_buf_1 _15490_ (.A(_09574_),
    .X(_09575_));
 sg13g2_a21o_1 _15491_ (.A2(_09210_),
    .A1(_09295_),
    .B1(_09077_),
    .X(_09576_));
 sg13g2_buf_1 _15492_ (.A(_09576_),
    .X(_09577_));
 sg13g2_a21oi_1 _15493_ (.A1(\top_ihp.oisc.decoder.instruction[20] ),
    .A2(_09575_),
    .Y(_09578_),
    .B1(_09577_));
 sg13g2_nor2_1 _15494_ (.A(_09556_),
    .B(_09578_),
    .Y(_09579_));
 sg13g2_nor2_1 _15495_ (.A(net245),
    .B(_09579_),
    .Y(_09580_));
 sg13g2_buf_8 _15496_ (.A(_09580_),
    .X(_09581_));
 sg13g2_nor2_1 _15497_ (.A(\top_ihp.oisc.regs[0][20] ),
    .B(_09108_),
    .Y(_09582_));
 sg13g2_a21oi_1 _15498_ (.A1(_09108_),
    .A2(_09581_),
    .Y(_00370_),
    .B1(_09582_));
 sg13g2_a21oi_1 _15499_ (.A1(_09542_),
    .A2(_09575_),
    .Y(_09583_),
    .B1(_09577_));
 sg13g2_nor2_2 _15500_ (.A(net1019),
    .B(net915),
    .Y(_09584_));
 sg13g2_nand2b_1 _15501_ (.Y(_09585_),
    .B(_09584_),
    .A_N(_09442_));
 sg13g2_nor2_1 _15502_ (.A(\top_ihp.wb_dati_rom[21] ),
    .B(_09166_),
    .Y(_09586_));
 sg13g2_and3_1 _15503_ (.X(_09587_),
    .A(_09144_),
    .B(\top_ihp.wb_dati_spi[21] ),
    .C(_09146_));
 sg13g2_a221oi_1 _15504_ (.B2(\top_ihp.wb_dati_ram[21] ),
    .C1(_09587_),
    .B1(net872),
    .A1(net884),
    .Y(_09588_),
    .A2(net846));
 sg13g2_nor3_2 _15505_ (.A(net951),
    .B(_09586_),
    .C(_09588_),
    .Y(_09589_));
 sg13g2_nand3_1 _15506_ (.B(_09584_),
    .C(_09589_),
    .A(net949),
    .Y(_09590_));
 sg13g2_nand3_1 _15507_ (.B(_09585_),
    .C(_09590_),
    .A(_09583_),
    .Y(_09591_));
 sg13g2_xnor2_1 _15508_ (.Y(_09592_),
    .A(_07462_),
    .B(_07913_));
 sg13g2_nand2_1 _15509_ (.Y(_09593_),
    .A(_09121_),
    .B(_09181_));
 sg13g2_a21oi_1 _15510_ (.A1(_07461_),
    .A2(_09592_),
    .Y(_09594_),
    .B1(_09593_));
 sg13g2_o21ai_1 _15511_ (.B1(_09188_),
    .Y(_09595_),
    .A1(_09591_),
    .A2(_09592_));
 sg13g2_nand2b_1 _15512_ (.Y(_09596_),
    .B(_09595_),
    .A_N(_07461_));
 sg13g2_o21ai_1 _15513_ (.B1(_09596_),
    .Y(_09597_),
    .A1(_09591_),
    .A2(_09594_));
 sg13g2_buf_2 _15514_ (.A(_09597_),
    .X(_09598_));
 sg13g2_buf_1 _15515_ (.A(_09598_),
    .X(_09599_));
 sg13g2_buf_1 _15516_ (.A(_09202_),
    .X(_09600_));
 sg13g2_nand2_1 _15517_ (.Y(_09601_),
    .A(\top_ihp.oisc.regs[0][21] ),
    .B(net546));
 sg13g2_o21ai_1 _15518_ (.B1(_09601_),
    .Y(_00371_),
    .A1(net410),
    .A2(net72));
 sg13g2_nand2_1 _15519_ (.Y(_09602_),
    .A(\top_ihp.wb_dati_ram[22] ),
    .B(net872));
 sg13g2_nand3_1 _15520_ (.B(\top_ihp.wb_dati_spi[22] ),
    .C(net841),
    .A(net918),
    .Y(_09603_));
 sg13g2_nand3_1 _15521_ (.B(_09602_),
    .C(_09603_),
    .A(net821),
    .Y(_09604_));
 sg13g2_o21ai_1 _15522_ (.B1(_09604_),
    .Y(_09605_),
    .A1(\top_ihp.wb_dati_rom[22] ),
    .A2(_09166_));
 sg13g2_nor2_1 _15523_ (.A(net951),
    .B(_09605_),
    .Y(_09606_));
 sg13g2_nand2_1 _15524_ (.Y(_09607_),
    .A(net949),
    .B(_09606_));
 sg13g2_a21oi_1 _15525_ (.A1(_09442_),
    .A2(_09607_),
    .Y(_09608_),
    .B1(net887));
 sg13g2_a21o_1 _15526_ (.A2(_09465_),
    .A1(_09464_),
    .B1(_08965_),
    .X(_09609_));
 sg13g2_a21oi_1 _15527_ (.A1(_07470_),
    .A2(_09609_),
    .Y(_09610_),
    .B1(_08960_));
 sg13g2_a21oi_1 _15528_ (.A1(_09464_),
    .A2(_09465_),
    .Y(_09611_),
    .B1(_08965_));
 sg13g2_nor3_1 _15529_ (.A(_07599_),
    .B(_07602_),
    .C(_09611_),
    .Y(_09612_));
 sg13g2_nor3_1 _15530_ (.A(_09290_),
    .B(_09610_),
    .C(_09612_),
    .Y(_09613_));
 sg13g2_nor3_1 _15531_ (.A(net948),
    .B(_09608_),
    .C(_09613_),
    .Y(_09614_));
 sg13g2_buf_1 _15532_ (.A(\top_ihp.oisc.decoder.instruction[22] ),
    .X(_09615_));
 sg13g2_nand2_1 _15533_ (.Y(_09616_),
    .A(_09115_),
    .B(_09208_));
 sg13g2_a21o_1 _15534_ (.A2(_09616_),
    .A1(_09295_),
    .B1(_09121_),
    .X(_09617_));
 sg13g2_buf_1 _15535_ (.A(_09617_),
    .X(_09618_));
 sg13g2_a21oi_1 _15536_ (.A1(_09615_),
    .A2(net883),
    .Y(_09619_),
    .B1(_09618_));
 sg13g2_nor3_1 _15537_ (.A(net860),
    .B(_09614_),
    .C(_09619_),
    .Y(_09620_));
 sg13g2_a21oi_1 _15538_ (.A1(_07444_),
    .A2(net859),
    .Y(_09621_),
    .B1(_09620_));
 sg13g2_buf_2 _15539_ (.A(_09621_),
    .X(_09622_));
 sg13g2_buf_2 _15540_ (.A(net244),
    .X(_09623_));
 sg13g2_nand2_1 _15541_ (.Y(_09624_),
    .A(\top_ihp.oisc.regs[0][22] ),
    .B(net546));
 sg13g2_o21ai_1 _15542_ (.B1(_09624_),
    .Y(_00372_),
    .A1(net410),
    .A2(net143));
 sg13g2_buf_1 _15543_ (.A(\top_ihp.oisc.decoder.instruction[23] ),
    .X(_09625_));
 sg13g2_a21oi_1 _15544_ (.A1(_09625_),
    .A2(net883),
    .Y(_09626_),
    .B1(_09618_));
 sg13g2_inv_1 _15545_ (.Y(_09627_),
    .A(_09217_));
 sg13g2_nand2_1 _15546_ (.Y(_09628_),
    .A(_09442_),
    .B(_09584_));
 sg13g2_a21oi_1 _15547_ (.A1(_09157_),
    .A2(_09627_),
    .Y(_09629_),
    .B1(_09628_));
 sg13g2_nand2b_1 _15548_ (.Y(_09630_),
    .B(_07444_),
    .A_N(net1044));
 sg13g2_nor2_1 _15549_ (.A(net1042),
    .B(_07454_),
    .Y(_09631_));
 sg13g2_nand2_1 _15550_ (.Y(_09632_),
    .A(_07452_),
    .B(_09631_));
 sg13g2_o21ai_1 _15551_ (.B1(_07451_),
    .Y(_09633_),
    .A1(_07452_),
    .A2(_09631_));
 sg13g2_nand2_1 _15552_ (.Y(_09634_),
    .A(_09632_),
    .B(_09633_));
 sg13g2_o21ai_1 _15553_ (.B1(_07467_),
    .Y(_09635_),
    .A1(_07464_),
    .A2(_09634_));
 sg13g2_nand2b_1 _15554_ (.Y(_09636_),
    .B(_09635_),
    .A_N(_07446_));
 sg13g2_nor2_1 _15555_ (.A(_07607_),
    .B(_07842_),
    .Y(_09637_));
 sg13g2_a22oi_1 _15556_ (.Y(_09638_),
    .B1(_09637_),
    .B2(_09493_),
    .A2(_09636_),
    .A1(_09630_));
 sg13g2_xor2_1 _15557_ (.B(_09638_),
    .A(_07600_),
    .X(_09639_));
 sg13g2_and2_1 _15558_ (.A(_09192_),
    .B(_09639_),
    .X(_09640_));
 sg13g2_nor4_2 _15559_ (.A(net860),
    .B(_09626_),
    .C(_09629_),
    .Y(_09641_),
    .D(_09640_));
 sg13g2_a21oi_1 _15560_ (.A1(_07442_),
    .A2(_09351_),
    .Y(_09642_),
    .B1(_09641_));
 sg13g2_buf_1 _15561_ (.A(_09642_),
    .X(_09643_));
 sg13g2_nor2_1 _15562_ (.A(\top_ihp.oisc.regs[0][23] ),
    .B(_09108_),
    .Y(_09644_));
 sg13g2_a21oi_1 _15563_ (.A1(_09108_),
    .A2(net243),
    .Y(_00373_),
    .B1(_09644_));
 sg13g2_a21oi_1 _15564_ (.A1(net952),
    .A2(_09172_),
    .Y(_09645_),
    .B1(_09180_));
 sg13g2_nor2_1 _15565_ (.A(_07630_),
    .B(_07632_),
    .Y(_09646_));
 sg13g2_xnor2_1 _15566_ (.Y(_09647_),
    .A(_09646_),
    .B(_07693_));
 sg13g2_a221oi_1 _15567_ (.B2(net887),
    .C1(net989),
    .B1(_09647_),
    .A1(_09442_),
    .Y(_09648_),
    .A2(_09645_));
 sg13g2_buf_1 _15568_ (.A(\top_ihp.oisc.decoder.instruction[24] ),
    .X(_09649_));
 sg13g2_a21oi_1 _15569_ (.A1(_09649_),
    .A2(_09575_),
    .Y(_09650_),
    .B1(_09577_));
 sg13g2_nand2b_1 _15570_ (.Y(_09651_),
    .B(_09650_),
    .A_N(_09648_));
 sg13g2_o21ai_1 _15571_ (.B1(_09651_),
    .Y(_09652_),
    .A1(net1029),
    .A2(_09205_));
 sg13g2_buf_1 _15572_ (.A(_09652_),
    .X(_09653_));
 sg13g2_buf_2 _15573_ (.A(_09653_),
    .X(_09654_));
 sg13g2_nand2_1 _15574_ (.Y(_09655_),
    .A(\top_ihp.oisc.regs[0][24] ),
    .B(_09600_));
 sg13g2_o21ai_1 _15575_ (.B1(_09655_),
    .Y(_00374_),
    .A1(net410),
    .A2(net242));
 sg13g2_nand2_1 _15576_ (.Y(_09656_),
    .A(_07621_),
    .B(net860));
 sg13g2_nor2_1 _15577_ (.A(_07803_),
    .B(_07842_),
    .Y(_09657_));
 sg13g2_a21oi_1 _15578_ (.A1(_07913_),
    .A2(_09657_),
    .Y(_09658_),
    .B1(_07810_));
 sg13g2_nor2_1 _15579_ (.A(_07694_),
    .B(net985),
    .Y(_09659_));
 sg13g2_xor2_1 _15580_ (.B(_09659_),
    .A(_09658_),
    .X(_09660_));
 sg13g2_a21oi_1 _15581_ (.A1(net952),
    .A2(_09520_),
    .Y(_09661_),
    .B1(net887));
 sg13g2_a22oi_1 _15582_ (.Y(_09662_),
    .B1(_09661_),
    .B2(_09442_),
    .A2(_09660_),
    .A1(net882));
 sg13g2_buf_1 _15583_ (.A(\top_ihp.oisc.decoder.instruction[25] ),
    .X(_09663_));
 sg13g2_a21oi_1 _15584_ (.A1(_09663_),
    .A2(_09310_),
    .Y(_09664_),
    .B1(_09618_));
 sg13g2_nor2_1 _15585_ (.A(_09123_),
    .B(_09664_),
    .Y(_09665_));
 sg13g2_o21ai_1 _15586_ (.B1(_09665_),
    .Y(_09666_),
    .A1(net948),
    .A2(_09662_));
 sg13g2_and2_1 _15587_ (.A(_09656_),
    .B(_09666_),
    .X(_09667_));
 sg13g2_buf_1 _15588_ (.A(_09667_),
    .X(_09668_));
 sg13g2_buf_2 _15589_ (.A(_09668_),
    .X(_09669_));
 sg13g2_nand2_1 _15590_ (.Y(_09670_),
    .A(\top_ihp.oisc.regs[0][25] ),
    .B(net546));
 sg13g2_o21ai_1 _15591_ (.B1(_09670_),
    .Y(_00375_),
    .A1(net410),
    .A2(net241));
 sg13g2_or4_1 _15592_ (.A(_07628_),
    .B(_07636_),
    .C(_07638_),
    .D(_07645_),
    .X(_09671_));
 sg13g2_buf_1 _15593_ (.A(\top_ihp.oisc.decoder.instruction[26] ),
    .X(_09672_));
 sg13g2_nand2b_1 _15594_ (.Y(_09673_),
    .B(net952),
    .A_N(_09257_));
 sg13g2_nor2_1 _15595_ (.A(_09189_),
    .B(_09430_),
    .Y(_09674_));
 sg13g2_a221oi_1 _15596_ (.B2(_09674_),
    .C1(_09577_),
    .B1(_09673_),
    .A1(_09672_),
    .Y(_09675_),
    .A2(_09575_));
 sg13g2_o21ai_1 _15597_ (.B1(_09675_),
    .Y(_09676_),
    .A1(_09671_),
    .A2(_09593_));
 sg13g2_o21ai_1 _15598_ (.B1(_09676_),
    .Y(_09677_),
    .A1(net1030),
    .A2(net871));
 sg13g2_buf_2 _15599_ (.A(_09677_),
    .X(_09678_));
 sg13g2_buf_1 _15600_ (.A(_09678_),
    .X(_09679_));
 sg13g2_nand2_1 _15601_ (.Y(_09680_),
    .A(\top_ihp.oisc.regs[0][26] ),
    .B(_09600_));
 sg13g2_o21ai_1 _15602_ (.B1(_09680_),
    .Y(_00376_),
    .A1(_09514_),
    .A2(net142));
 sg13g2_nand3_1 _15603_ (.B(_07613_),
    .C(_07624_),
    .A(net1030),
    .Y(_09681_));
 sg13g2_nand3_1 _15604_ (.B(net1029),
    .C(_07624_),
    .A(net1030),
    .Y(_09682_));
 sg13g2_a22oi_1 _15605_ (.Y(_09683_),
    .B1(_09681_),
    .B2(_09682_),
    .A2(_07611_),
    .A1(_07598_));
 sg13g2_nand2_1 _15606_ (.Y(_09684_),
    .A(net1030),
    .B(net985));
 sg13g2_o21ai_1 _15607_ (.B1(_09684_),
    .Y(_09685_),
    .A1(_07612_),
    .A2(_09682_));
 sg13g2_nor2_1 _15608_ (.A(_09683_),
    .B(_09685_),
    .Y(_09686_));
 sg13g2_a21o_1 _15609_ (.A2(_09309_),
    .A1(\top_ihp.oisc.decoder.instruction[27] ),
    .B1(_09618_),
    .X(_09687_));
 sg13g2_buf_1 _15610_ (.A(_09687_),
    .X(_09688_));
 sg13g2_nand3b_1 _15611_ (.B(net915),
    .C(_09688_),
    .Y(_09689_),
    .A_N(_07697_));
 sg13g2_a21oi_1 _15612_ (.A1(_09245_),
    .A2(_09285_),
    .Y(_09690_),
    .B1(_09430_));
 sg13g2_o21ai_1 _15613_ (.B1(_09688_),
    .Y(_09691_),
    .A1(net989),
    .A2(_09690_));
 sg13g2_o21ai_1 _15614_ (.B1(_09691_),
    .Y(_09692_),
    .A1(_09686_),
    .A2(_09689_));
 sg13g2_a221oi_1 _15615_ (.B2(_09657_),
    .C1(_07810_),
    .B1(_07913_),
    .A1(_07811_),
    .Y(_09693_),
    .A2(_07622_));
 sg13g2_nor3_1 _15616_ (.A(net1030),
    .B(net985),
    .C(_09693_),
    .Y(_09694_));
 sg13g2_or3_1 _15617_ (.A(_07615_),
    .B(_09694_),
    .C(_09689_),
    .X(_09695_));
 sg13g2_nand3_1 _15618_ (.B(net915),
    .C(_09688_),
    .A(_07697_),
    .Y(_09696_));
 sg13g2_nor3_1 _15619_ (.A(_09683_),
    .B(_09685_),
    .C(_09696_),
    .Y(_09697_));
 sg13g2_o21ai_1 _15620_ (.B1(_09697_),
    .Y(_09698_),
    .A1(_07615_),
    .A2(_09694_));
 sg13g2_nand3b_1 _15621_ (.B(_09695_),
    .C(_09698_),
    .Y(_09699_),
    .A_N(_09692_));
 sg13g2_or2_1 _15622_ (.X(_09700_),
    .B(_09205_),
    .A(_07681_));
 sg13g2_o21ai_1 _15623_ (.B1(_09700_),
    .Y(_09701_),
    .A1(_09351_),
    .A2(_09699_));
 sg13g2_buf_8 _15624_ (.A(_09701_),
    .X(_09702_));
 sg13g2_buf_8 _15625_ (.A(net141),
    .X(_09703_));
 sg13g2_nand2_1 _15626_ (.Y(_09704_),
    .A(\top_ihp.oisc.regs[0][27] ),
    .B(net546));
 sg13g2_o21ai_1 _15627_ (.B1(_09704_),
    .Y(_00377_),
    .A1(_09514_),
    .A2(net71));
 sg13g2_buf_1 _15628_ (.A(\top_ihp.oisc.decoder.instruction[28] ),
    .X(_09705_));
 sg13g2_a21o_1 _15629_ (.A2(_09340_),
    .A1(_09245_),
    .B1(_09443_),
    .X(_09706_));
 sg13g2_a221oi_1 _15630_ (.B2(_09706_),
    .C1(_09577_),
    .B1(_09584_),
    .A1(_09705_),
    .Y(_09707_),
    .A2(_09575_));
 sg13g2_a21oi_1 _15631_ (.A1(_07705_),
    .A2(_09707_),
    .Y(_09708_),
    .B1(net867));
 sg13g2_nor3_1 _15632_ (.A(_07701_),
    .B(_07703_),
    .C(_07704_),
    .Y(_09709_));
 sg13g2_a21oi_1 _15633_ (.A1(net1028),
    .A2(_09709_),
    .Y(_09710_),
    .B1(_09593_));
 sg13g2_nand2b_1 _15634_ (.Y(_09711_),
    .B(_09707_),
    .A_N(_09710_));
 sg13g2_o21ai_1 _15635_ (.B1(_09711_),
    .Y(_09712_),
    .A1(net1028),
    .A2(_09708_));
 sg13g2_buf_2 _15636_ (.A(_09712_),
    .X(_09713_));
 sg13g2_buf_8 _15637_ (.A(_09713_),
    .X(_09714_));
 sg13g2_nand2_1 _15638_ (.Y(_09715_),
    .A(\top_ihp.oisc.regs[0][28] ),
    .B(net546));
 sg13g2_o21ai_1 _15639_ (.B1(_09715_),
    .Y(_00378_),
    .A1(net410),
    .A2(net70));
 sg13g2_a21oi_1 _15640_ (.A1(\top_ihp.oisc.decoder.instruction[29] ),
    .A2(_09310_),
    .Y(_09716_),
    .B1(_09618_));
 sg13g2_a21oi_1 _15641_ (.A1(_09157_),
    .A2(_09361_),
    .Y(_09717_),
    .B1(_09628_));
 sg13g2_nor3_1 _15642_ (.A(_09350_),
    .B(_09716_),
    .C(_09717_),
    .Y(_09718_));
 sg13g2_a21oi_1 _15643_ (.A1(_07913_),
    .A2(_07845_),
    .Y(_09719_),
    .B1(_07839_));
 sg13g2_xnor2_1 _15644_ (.Y(_09720_),
    .A(_07916_),
    .B(_09719_));
 sg13g2_nand2_1 _15645_ (.Y(_09721_),
    .A(_09192_),
    .B(_09720_));
 sg13g2_a22oi_1 _15646_ (.Y(_09722_),
    .B1(_09718_),
    .B2(_09721_),
    .A2(net859),
    .A1(_07721_));
 sg13g2_buf_1 _15647_ (.A(_09722_),
    .X(_09723_));
 sg13g2_buf_2 _15648_ (.A(_09723_),
    .X(_09724_));
 sg13g2_nand2_1 _15649_ (.Y(_09725_),
    .A(\top_ihp.oisc.regs[0][29] ),
    .B(net546));
 sg13g2_o21ai_1 _15650_ (.B1(_09725_),
    .Y(_00379_),
    .A1(net410),
    .A2(net140));
 sg13g2_nor2_1 _15651_ (.A(net992),
    .B(_08216_),
    .Y(_09726_));
 sg13g2_and2_1 _15652_ (.A(_09143_),
    .B(\top_ihp.wb_dati_spi[2] ),
    .X(_09727_));
 sg13g2_mux2_1 _15653_ (.A0(\top_ihp.wb_dati_ram[2] ),
    .A1(_09727_),
    .S(net839),
    .X(_09728_));
 sg13g2_mux2_1 _15654_ (.A0(\top_ihp.wb_dati_rom[2] ),
    .A1(_09728_),
    .S(net840),
    .X(_09729_));
 sg13g2_and2_1 _15655_ (.A(net992),
    .B(\top_ihp.wb_dati_uart[2] ),
    .X(_09730_));
 sg13g2_a21o_1 _15656_ (.A2(_09729_),
    .A1(_09726_),
    .B1(_09730_),
    .X(_09731_));
 sg13g2_buf_1 _15657_ (.A(_09731_),
    .X(_09732_));
 sg13g2_a21oi_1 _15658_ (.A1(_09726_),
    .A2(_09729_),
    .Y(_09733_),
    .B1(_09730_));
 sg13g2_buf_2 _15659_ (.A(_09733_),
    .X(_09734_));
 sg13g2_nand2_1 _15660_ (.Y(_09735_),
    .A(_09140_),
    .B(_09473_));
 sg13g2_o21ai_1 _15661_ (.B1(_09735_),
    .Y(_09736_),
    .A1(net991),
    .A2(_09734_));
 sg13g2_a21oi_1 _15662_ (.A1(net991),
    .A2(_09257_),
    .Y(_09737_),
    .B1(_09258_));
 sg13g2_nor2_1 _15663_ (.A(_09160_),
    .B(_09737_),
    .Y(_09738_));
 sg13g2_a221oi_1 _15664_ (.B2(_09528_),
    .C1(_09738_),
    .B1(_09736_),
    .A1(net952),
    .Y(_09739_),
    .A2(_09732_));
 sg13g2_xnor2_1 _15665_ (.Y(_09740_),
    .A(_07472_),
    .B(_07481_));
 sg13g2_xor2_1 _15666_ (.B(_09740_),
    .A(net1040),
    .X(_09741_));
 sg13g2_mux2_1 _15667_ (.A0(_09739_),
    .A1(_09741_),
    .S(net887),
    .X(_09742_));
 sg13g2_nand2_1 _15668_ (.Y(_09743_),
    .A(net955),
    .B(_09742_));
 sg13g2_and2_1 _15669_ (.A(_09109_),
    .B(_09099_),
    .X(_09744_));
 sg13g2_a21oi_1 _15670_ (.A1(_09114_),
    .A2(_09615_),
    .Y(_09745_),
    .B1(_09744_));
 sg13g2_nand2_1 _15671_ (.Y(_09746_),
    .A(_09099_),
    .B(_09546_));
 sg13g2_o21ai_1 _15672_ (.B1(_09746_),
    .Y(_09747_),
    .A1(_09118_),
    .A2(_09745_));
 sg13g2_nand2_1 _15673_ (.Y(_09748_),
    .A(net956),
    .B(_09615_));
 sg13g2_o21ai_1 _15674_ (.B1(_09748_),
    .Y(_09749_),
    .A1(_09110_),
    .A2(_00100_));
 sg13g2_a22oi_1 _15675_ (.Y(_09750_),
    .B1(_09749_),
    .B2(_09311_),
    .A2(_09747_),
    .A1(net995));
 sg13g2_a21oi_1 _15676_ (.A1(net948),
    .A2(_09750_),
    .Y(_09751_),
    .B1(_09307_));
 sg13g2_a22oi_1 _15677_ (.Y(_09752_),
    .B1(_09743_),
    .B2(_09751_),
    .A2(net859),
    .A1(net1040));
 sg13g2_buf_2 _15678_ (.A(_09752_),
    .X(_09753_));
 sg13g2_buf_2 _15679_ (.A(_09753_),
    .X(_09754_));
 sg13g2_nand2_1 _15680_ (.Y(_09755_),
    .A(\top_ihp.oisc.regs[0][2] ),
    .B(net546));
 sg13g2_o21ai_1 _15681_ (.B1(_09755_),
    .Y(_00380_),
    .A1(net410),
    .A2(net240));
 sg13g2_nand2_1 _15682_ (.Y(_09756_),
    .A(_07738_),
    .B(_09192_));
 sg13g2_a21o_1 _15683_ (.A2(_09389_),
    .A1(net952),
    .B1(_09443_),
    .X(_09757_));
 sg13g2_a221oi_1 _15684_ (.B2(_09757_),
    .C1(_09577_),
    .B1(_09584_),
    .A1(\top_ihp.oisc.decoder.instruction[30] ),
    .Y(_09758_),
    .A2(_09575_));
 sg13g2_nand2_1 _15685_ (.Y(_09759_),
    .A(_09756_),
    .B(_09758_));
 sg13g2_o21ai_1 _15686_ (.B1(_09759_),
    .Y(_09760_),
    .A1(net1026),
    .A2(net871));
 sg13g2_buf_2 _15687_ (.A(_09760_),
    .X(_09761_));
 sg13g2_buf_2 _15688_ (.A(_09761_),
    .X(_09762_));
 sg13g2_nand2_1 _15689_ (.Y(_09763_),
    .A(\top_ihp.oisc.regs[0][30] ),
    .B(net546));
 sg13g2_o21ai_1 _15690_ (.B1(_09763_),
    .Y(_00381_),
    .A1(_09271_),
    .A2(net69));
 sg13g2_nor2_1 _15691_ (.A(_09593_),
    .B(net860),
    .Y(_09764_));
 sg13g2_nor2b_1 _15692_ (.A(_07697_),
    .B_N(_08949_),
    .Y(_09765_));
 sg13g2_and2_1 _15693_ (.A(_07615_),
    .B(_09765_),
    .X(_09766_));
 sg13g2_o21ai_1 _15694_ (.B1(_07914_),
    .Y(_09767_),
    .A1(_07815_),
    .A2(_07834_));
 sg13g2_inv_1 _15695_ (.Y(_09768_),
    .A(_07719_));
 sg13g2_o21ai_1 _15696_ (.B1(_09768_),
    .Y(_09769_),
    .A1(net1026),
    .A2(_09767_));
 sg13g2_nand2_1 _15697_ (.Y(_09770_),
    .A(net1026),
    .B(_09767_));
 sg13g2_a21o_1 _15698_ (.A2(_09770_),
    .A1(_09769_),
    .B1(_08948_),
    .X(_09771_));
 sg13g2_a221oi_1 _15699_ (.B2(_09686_),
    .C1(_09771_),
    .B1(_09766_),
    .A1(_09694_),
    .Y(_09772_),
    .A2(_09765_));
 sg13g2_nor2_1 _15700_ (.A(_08982_),
    .B(_09772_),
    .Y(_09773_));
 sg13g2_and2_1 _15701_ (.A(_09189_),
    .B(_09295_),
    .X(_09774_));
 sg13g2_a21o_1 _15702_ (.A2(_09207_),
    .A1(_09119_),
    .B1(net995),
    .X(_09775_));
 sg13g2_nand2_1 _15703_ (.Y(_09776_),
    .A(net917),
    .B(_09235_));
 sg13g2_a22oi_1 _15704_ (.Y(_09777_),
    .B1(_09776_),
    .B2(_09674_),
    .A2(_09775_),
    .A1(_09774_));
 sg13g2_nor2_1 _15705_ (.A(_08946_),
    .B(net886),
    .Y(_09778_));
 sg13g2_a21oi_1 _15706_ (.A1(net871),
    .A2(_09777_),
    .Y(_09779_),
    .B1(_09778_));
 sg13g2_a21oi_1 _15707_ (.A1(_09764_),
    .A2(_09773_),
    .Y(_09780_),
    .B1(_09779_));
 sg13g2_buf_2 _15708_ (.A(_09780_),
    .X(_09781_));
 sg13g2_buf_8 _15709_ (.A(_09781_),
    .X(_09782_));
 sg13g2_nand2_1 _15710_ (.Y(_09783_),
    .A(\top_ihp.oisc.regs[0][31] ),
    .B(_09203_));
 sg13g2_o21ai_1 _15711_ (.B1(_09783_),
    .Y(_00382_),
    .A1(net549),
    .A2(net139));
 sg13g2_or3_1 _15712_ (.A(_09161_),
    .B(_09160_),
    .C(_09277_),
    .X(_09784_));
 sg13g2_or2_1 _15713_ (.X(_09785_),
    .B(_09285_),
    .A(_09160_));
 sg13g2_and2_1 _15714_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[3] ),
    .X(_09786_));
 sg13g2_mux2_1 _15715_ (.A0(\top_ihp.wb_dati_ram[3] ),
    .A1(_09786_),
    .S(net839),
    .X(_09787_));
 sg13g2_mux2_1 _15716_ (.A0(\top_ihp.wb_dati_rom[3] ),
    .A1(_09787_),
    .S(_09165_),
    .X(_09788_));
 sg13g2_a22oi_1 _15717_ (.Y(_09789_),
    .B1(_09726_),
    .B2(_09788_),
    .A2(\top_ihp.wb_dati_uart[3] ),
    .A1(net992));
 sg13g2_buf_1 _15718_ (.A(_09789_),
    .X(_09790_));
 sg13g2_a22oi_1 _15719_ (.Y(_09791_),
    .B1(_09790_),
    .B2(_09160_),
    .A2(_09785_),
    .A1(_09140_));
 sg13g2_nor2_1 _15720_ (.A(_09127_),
    .B(_09279_),
    .Y(_09792_));
 sg13g2_a221oi_1 _15721_ (.B2(_09502_),
    .C1(net882),
    .B1(_09792_),
    .A1(_09784_),
    .Y(_09793_),
    .A2(_09791_));
 sg13g2_xor2_1 _15722_ (.B(_07484_),
    .A(_07485_),
    .X(_09794_));
 sg13g2_xnor2_1 _15723_ (.Y(_09795_),
    .A(net1037),
    .B(_09794_));
 sg13g2_nor2_1 _15724_ (.A(net913),
    .B(_09795_),
    .Y(_09796_));
 sg13g2_o21ai_1 _15725_ (.B1(net955),
    .Y(_09797_),
    .A1(_09793_),
    .A2(_09796_));
 sg13g2_and2_1 _15726_ (.A(net996),
    .B(_09096_),
    .X(_09798_));
 sg13g2_a21oi_1 _15727_ (.A1(_09114_),
    .A2(_09625_),
    .Y(_09799_),
    .B1(_09798_));
 sg13g2_nand2_1 _15728_ (.Y(_09800_),
    .A(_09096_),
    .B(_09546_));
 sg13g2_o21ai_1 _15729_ (.B1(_09800_),
    .Y(_09801_),
    .A1(net994),
    .A2(_09799_));
 sg13g2_nand2_1 _15730_ (.Y(_09802_),
    .A(net956),
    .B(_09625_));
 sg13g2_o21ai_1 _15731_ (.B1(_09802_),
    .Y(_09803_),
    .A1(net956),
    .A2(_00101_));
 sg13g2_a22oi_1 _15732_ (.Y(_09804_),
    .B1(_09803_),
    .B2(_09311_),
    .A2(_09801_),
    .A1(_09111_));
 sg13g2_a21oi_1 _15733_ (.A1(_09294_),
    .A2(_09804_),
    .Y(_09805_),
    .B1(_09307_));
 sg13g2_a22oi_1 _15734_ (.Y(_09806_),
    .B1(_09797_),
    .B2(_09805_),
    .A2(net859),
    .A1(net1037));
 sg13g2_buf_1 _15735_ (.A(_09806_),
    .X(_09807_));
 sg13g2_buf_2 _15736_ (.A(_09807_),
    .X(_09808_));
 sg13g2_nand2_1 _15737_ (.Y(_09809_),
    .A(\top_ihp.oisc.regs[0][3] ),
    .B(net550));
 sg13g2_o21ai_1 _15738_ (.B1(_09809_),
    .Y(_00383_),
    .A1(_09271_),
    .A2(net238));
 sg13g2_and2_1 _15739_ (.A(net996),
    .B(_09087_),
    .X(_09810_));
 sg13g2_a21oi_1 _15740_ (.A1(_09114_),
    .A2(_09649_),
    .Y(_09811_),
    .B1(_09810_));
 sg13g2_nand2_1 _15741_ (.Y(_09812_),
    .A(_09087_),
    .B(_09546_));
 sg13g2_o21ai_1 _15742_ (.B1(_09812_),
    .Y(_09813_),
    .A1(_09118_),
    .A2(_09811_));
 sg13g2_nand2_1 _15743_ (.Y(_09814_),
    .A(net996),
    .B(_09649_));
 sg13g2_o21ai_1 _15744_ (.B1(_09814_),
    .Y(_09815_),
    .A1(_09110_),
    .A2(_00102_));
 sg13g2_a22oi_1 _15745_ (.Y(_09816_),
    .B1(_09815_),
    .B2(_09311_),
    .A2(_09813_),
    .A1(_09111_));
 sg13g2_nand2_1 _15746_ (.Y(_09817_),
    .A(_08215_),
    .B(\top_ihp.wb_dati_uart[4] ));
 sg13g2_nor2_1 _15747_ (.A(\top_ihp.wb_dati_rom[4] ),
    .B(net862),
    .Y(_09818_));
 sg13g2_and2_1 _15748_ (.A(net1012),
    .B(\top_ihp.wb_dati_spi[4] ),
    .X(_09819_));
 sg13g2_inv_1 _15749_ (.Y(_09820_),
    .A(\top_ihp.wb_dati_ram[4] ));
 sg13g2_nor4_1 _15750_ (.A(_09248_),
    .B(_09820_),
    .C(net885),
    .D(net903),
    .Y(_09821_));
 sg13g2_a221oi_1 _15751_ (.B2(_09819_),
    .C1(_09821_),
    .B1(net861),
    .A1(net950),
    .Y(_09822_),
    .A2(net863));
 sg13g2_or3_1 _15752_ (.A(net980),
    .B(_09818_),
    .C(_09822_),
    .X(_09823_));
 sg13g2_nand2_1 _15753_ (.Y(_09824_),
    .A(_09817_),
    .B(_09823_));
 sg13g2_buf_1 _15754_ (.A(_09824_),
    .X(_09825_));
 sg13g2_and2_1 _15755_ (.A(_09817_),
    .B(_09823_),
    .X(_09826_));
 sg13g2_buf_1 _15756_ (.A(_09826_),
    .X(_09827_));
 sg13g2_nand2_1 _15757_ (.Y(_09828_),
    .A(_09140_),
    .B(_09569_));
 sg13g2_o21ai_1 _15758_ (.B1(_09828_),
    .Y(_09829_),
    .A1(net1018),
    .A2(_09827_));
 sg13g2_nand2_1 _15759_ (.Y(_09830_),
    .A(net1018),
    .B(_09340_));
 sg13g2_a21oi_1 _15760_ (.A1(_09333_),
    .A2(_09830_),
    .Y(_09831_),
    .B1(_09160_));
 sg13g2_a221oi_1 _15761_ (.B2(_09528_),
    .C1(_09831_),
    .B1(_09829_),
    .A1(net993),
    .Y(_09832_),
    .A2(_09825_));
 sg13g2_nor2_1 _15762_ (.A(_07852_),
    .B(_07856_),
    .Y(_09833_));
 sg13g2_xnor2_1 _15763_ (.Y(_09834_),
    .A(_07486_),
    .B(_09833_));
 sg13g2_xnor2_1 _15764_ (.Y(_09835_),
    .A(net1039),
    .B(_09834_));
 sg13g2_mux2_1 _15765_ (.A0(_09832_),
    .A1(_09835_),
    .S(net915),
    .X(_09836_));
 sg13g2_mux2_1 _15766_ (.A0(_09816_),
    .A1(_09836_),
    .S(_09121_),
    .X(_09837_));
 sg13g2_nand2_1 _15767_ (.Y(_09838_),
    .A(net886),
    .B(_09837_));
 sg13g2_o21ai_1 _15768_ (.B1(_09838_),
    .Y(_09839_),
    .A1(net1039),
    .A2(net871));
 sg13g2_buf_1 _15769_ (.A(_09839_),
    .X(_09840_));
 sg13g2_buf_2 _15770_ (.A(_09840_),
    .X(_09841_));
 sg13g2_nand2_1 _15771_ (.Y(_09842_),
    .A(\top_ihp.oisc.regs[0][4] ),
    .B(net550));
 sg13g2_o21ai_1 _15772_ (.B1(_09842_),
    .Y(_00384_),
    .A1(net549),
    .A2(net237));
 sg13g2_a21oi_1 _15773_ (.A1(net991),
    .A2(_09361_),
    .Y(_09843_),
    .B1(_09364_));
 sg13g2_nor2_1 _15774_ (.A(\top_ihp.wb_dati_rom[5] ),
    .B(net862),
    .Y(_09844_));
 sg13g2_and2_1 _15775_ (.A(net1012),
    .B(\top_ihp.wb_dati_spi[5] ),
    .X(_09845_));
 sg13g2_inv_1 _15776_ (.Y(_09846_),
    .A(\top_ihp.wb_dati_ram[5] ));
 sg13g2_nor4_1 _15777_ (.A(net981),
    .B(_09846_),
    .C(_09221_),
    .D(net903),
    .Y(_09847_));
 sg13g2_a221oi_1 _15778_ (.B2(_09845_),
    .C1(_09847_),
    .B1(net861),
    .A1(_09168_),
    .Y(_09848_),
    .A2(net878));
 sg13g2_or3_1 _15779_ (.A(net980),
    .B(_09844_),
    .C(_09848_),
    .X(_09849_));
 sg13g2_buf_1 _15780_ (.A(_09849_),
    .X(_09850_));
 sg13g2_nand2_1 _15781_ (.Y(_09851_),
    .A(_08215_),
    .B(\top_ihp.wb_dati_uart[5] ));
 sg13g2_nand2_1 _15782_ (.Y(_09852_),
    .A(_09850_),
    .B(_09851_));
 sg13g2_buf_2 _15783_ (.A(_09852_),
    .X(_09853_));
 sg13g2_and2_1 _15784_ (.A(_09850_),
    .B(_09851_),
    .X(_09854_));
 sg13g2_buf_1 _15785_ (.A(_09854_),
    .X(_09855_));
 sg13g2_nor2_1 _15786_ (.A(net954),
    .B(_09589_),
    .Y(_09856_));
 sg13g2_a21oi_1 _15787_ (.A1(_09138_),
    .A2(net736),
    .Y(_09857_),
    .B1(_09856_));
 sg13g2_nor2_1 _15788_ (.A(net949),
    .B(_09127_),
    .Y(_09858_));
 sg13g2_a22oi_1 _15789_ (.Y(_09859_),
    .B1(_09857_),
    .B2(_09858_),
    .A2(_09853_),
    .A1(net952));
 sg13g2_o21ai_1 _15790_ (.B1(_09859_),
    .Y(_09860_),
    .A1(_09160_),
    .A2(_09843_));
 sg13g2_a21oi_1 _15791_ (.A1(_07488_),
    .A2(_09833_),
    .Y(_09861_),
    .B1(_07501_));
 sg13g2_xnor2_1 _15792_ (.Y(_09862_),
    .A(_07502_),
    .B(_09861_));
 sg13g2_and2_1 _15793_ (.A(net1038),
    .B(net915),
    .X(_09863_));
 sg13g2_a21oi_1 _15794_ (.A1(_09862_),
    .A2(_09863_),
    .Y(_09864_),
    .B1(net948));
 sg13g2_o21ai_1 _15795_ (.B1(_09864_),
    .Y(_09865_),
    .A1(net882),
    .A2(_09860_));
 sg13g2_a21oi_1 _15796_ (.A1(_09663_),
    .A2(net870),
    .Y(_09866_),
    .B1(net867));
 sg13g2_a21oi_1 _15797_ (.A1(_09663_),
    .A2(net870),
    .Y(_09867_),
    .B1(net913));
 sg13g2_nand2b_1 _15798_ (.Y(_09868_),
    .B(_09867_),
    .A_N(_09862_));
 sg13g2_a21oi_1 _15799_ (.A1(net886),
    .A2(_09868_),
    .Y(_09869_),
    .B1(net1038));
 sg13g2_a21o_1 _15800_ (.A2(_09866_),
    .A1(_09865_),
    .B1(_09869_),
    .X(_09870_));
 sg13g2_buf_2 _15801_ (.A(_09870_),
    .X(_09871_));
 sg13g2_buf_2 _15802_ (.A(_09871_),
    .X(_09872_));
 sg13g2_nand2_1 _15803_ (.Y(_09873_),
    .A(\top_ihp.oisc.regs[0][5] ),
    .B(net550));
 sg13g2_o21ai_1 _15804_ (.B1(_09873_),
    .Y(_00385_),
    .A1(net549),
    .A2(net236));
 sg13g2_xnor2_1 _15805_ (.Y(_09874_),
    .A(_07551_),
    .B(_07506_));
 sg13g2_a21oi_1 _15806_ (.A1(_09672_),
    .A2(net870),
    .Y(_09875_),
    .B1(net913));
 sg13g2_a21oi_1 _15807_ (.A1(_09874_),
    .A2(_09875_),
    .Y(_09876_),
    .B1(net867));
 sg13g2_nor2_1 _15808_ (.A(\top_ihp.wb_dati_rom[6] ),
    .B(_09165_),
    .Y(_09877_));
 sg13g2_and2_1 _15809_ (.A(net953),
    .B(\top_ihp.wb_dati_spi[6] ),
    .X(_09878_));
 sg13g2_inv_1 _15810_ (.Y(_09879_),
    .A(\top_ihp.wb_dati_ram[6] ));
 sg13g2_nor4_1 _15811_ (.A(net914),
    .B(_09879_),
    .C(net885),
    .D(_09250_),
    .Y(_09880_));
 sg13g2_a221oi_1 _15812_ (.B2(_09878_),
    .C1(_09880_),
    .B1(_09174_),
    .A1(net916),
    .Y(_09881_),
    .A2(net863));
 sg13g2_or3_1 _15813_ (.A(net980),
    .B(_09877_),
    .C(_09881_),
    .X(_09882_));
 sg13g2_buf_1 _15814_ (.A(_09882_),
    .X(_09883_));
 sg13g2_nand2_1 _15815_ (.Y(_09884_),
    .A(net992),
    .B(\top_ihp.wb_dati_uart[6] ));
 sg13g2_nand2_1 _15816_ (.Y(_09885_),
    .A(_09883_),
    .B(_09884_));
 sg13g2_mux2_1 _15817_ (.A0(_09606_),
    .A1(_09885_),
    .S(net954),
    .X(_09886_));
 sg13g2_o21ai_1 _15818_ (.B1(_09191_),
    .Y(_09887_),
    .A1(_09160_),
    .A2(_09393_));
 sg13g2_a221oi_1 _15819_ (.B2(_09858_),
    .C1(_09887_),
    .B1(_09886_),
    .A1(net952),
    .Y(_09888_),
    .A2(_09885_));
 sg13g2_nand2_1 _15820_ (.Y(_09889_),
    .A(net1031),
    .B(net887));
 sg13g2_o21ai_1 _15821_ (.B1(net955),
    .Y(_09890_),
    .A1(_09874_),
    .A2(_09889_));
 sg13g2_a21oi_1 _15822_ (.A1(_09672_),
    .A2(net870),
    .Y(_09891_),
    .B1(net873));
 sg13g2_o21ai_1 _15823_ (.B1(_09891_),
    .Y(_09892_),
    .A1(_09888_),
    .A2(_09890_));
 sg13g2_o21ai_1 _15824_ (.B1(_09892_),
    .Y(_09893_),
    .A1(net1031),
    .A2(_09876_));
 sg13g2_buf_2 _15825_ (.A(_09893_),
    .X(_09894_));
 sg13g2_buf_2 _15826_ (.A(_09894_),
    .X(_09895_));
 sg13g2_nand2_1 _15827_ (.Y(_09896_),
    .A(\top_ihp.oisc.regs[0][6] ),
    .B(net550));
 sg13g2_o21ai_1 _15828_ (.B1(_09896_),
    .Y(_00386_),
    .A1(net549),
    .A2(net235));
 sg13g2_nor2_1 _15829_ (.A(_07552_),
    .B(_07506_),
    .Y(_09897_));
 sg13g2_a21oi_1 _15830_ (.A1(_07552_),
    .A2(_07506_),
    .Y(_09898_),
    .B1(net1031));
 sg13g2_nor2_1 _15831_ (.A(_09897_),
    .B(_09898_),
    .Y(_09899_));
 sg13g2_xnor2_1 _15832_ (.Y(_09900_),
    .A(_07540_),
    .B(_09899_));
 sg13g2_xor2_1 _15833_ (.B(_09900_),
    .A(net1033),
    .X(_09901_));
 sg13g2_nand2_1 _15834_ (.Y(_09902_),
    .A(net992),
    .B(\top_ihp.wb_dati_uart[7] ));
 sg13g2_a21oi_1 _15835_ (.A1(_09225_),
    .A2(_09902_),
    .Y(_09903_),
    .B1(_09278_));
 sg13g2_nand2_1 _15836_ (.Y(_09904_),
    .A(_09528_),
    .B(_09228_));
 sg13g2_nand2_1 _15837_ (.Y(_09905_),
    .A(_09127_),
    .B(_09238_));
 sg13g2_a21oi_1 _15838_ (.A1(_09904_),
    .A2(_09905_),
    .Y(_09906_),
    .B1(net993));
 sg13g2_o21ai_1 _15839_ (.B1(_09191_),
    .Y(_09907_),
    .A1(_09903_),
    .A2(_09906_));
 sg13g2_o21ai_1 _15840_ (.B1(_09907_),
    .Y(_09908_),
    .A1(_09191_),
    .A2(_09901_));
 sg13g2_a221oi_1 _15841_ (.B2(net955),
    .C1(net873),
    .B1(_09908_),
    .A1(\top_ihp.oisc.decoder.instruction[27] ),
    .Y(_09909_),
    .A2(_09210_));
 sg13g2_buf_2 _15842_ (.A(_09909_),
    .X(_09910_));
 sg13g2_nor2_1 _15843_ (.A(net1033),
    .B(net871),
    .Y(_09911_));
 sg13g2_or2_1 _15844_ (.X(_09912_),
    .B(_09911_),
    .A(net408));
 sg13g2_buf_1 _15845_ (.A(_09912_),
    .X(_09913_));
 sg13g2_buf_2 _15846_ (.A(_09913_),
    .X(_09914_));
 sg13g2_nand2_1 _15847_ (.Y(_09915_),
    .A(\top_ihp.oisc.regs[0][7] ),
    .B(net550));
 sg13g2_o21ai_1 _15848_ (.B1(_09915_),
    .Y(_00387_),
    .A1(net549),
    .A2(net68));
 sg13g2_o21ai_1 _15849_ (.B1(_07871_),
    .Y(_09916_),
    .A1(_07542_),
    .A2(_09899_));
 sg13g2_xnor2_1 _15850_ (.Y(_09917_),
    .A(_07581_),
    .B(_09916_));
 sg13g2_a21oi_1 _15851_ (.A1(_09705_),
    .A2(net870),
    .Y(_09918_),
    .B1(net913));
 sg13g2_a21oi_1 _15852_ (.A1(_09917_),
    .A2(_09918_),
    .Y(_09919_),
    .B1(net867));
 sg13g2_nand2_1 _15853_ (.Y(_09920_),
    .A(net1015),
    .B(net887));
 sg13g2_nand2_1 _15854_ (.Y(_09921_),
    .A(net949),
    .B(_09177_));
 sg13g2_and2_1 _15855_ (.A(_09140_),
    .B(_09172_),
    .X(_09922_));
 sg13g2_o21ai_1 _15856_ (.B1(net988),
    .Y(_09923_),
    .A1(_09178_),
    .A2(_09922_));
 sg13g2_nand3_1 _15857_ (.B(_09921_),
    .C(_09923_),
    .A(_09244_),
    .Y(_09924_));
 sg13g2_o21ai_1 _15858_ (.B1(_09924_),
    .Y(_09925_),
    .A1(_09917_),
    .A2(_09920_));
 sg13g2_a21oi_1 _15859_ (.A1(_09705_),
    .A2(net870),
    .Y(_09926_),
    .B1(net873));
 sg13g2_o21ai_1 _15860_ (.B1(_09926_),
    .Y(_09927_),
    .A1(net948),
    .A2(_09925_));
 sg13g2_o21ai_1 _15861_ (.B1(_09927_),
    .Y(_09928_),
    .A1(net1015),
    .A2(_09919_));
 sg13g2_buf_2 _15862_ (.A(_09928_),
    .X(_09929_));
 sg13g2_buf_2 _15863_ (.A(_09929_),
    .X(_09930_));
 sg13g2_nand2_1 _15864_ (.Y(_09931_),
    .A(\top_ihp.oisc.regs[0][8] ),
    .B(net550));
 sg13g2_o21ai_1 _15865_ (.B1(_09931_),
    .Y(_00388_),
    .A1(net549),
    .A2(net67));
 sg13g2_inv_1 _15866_ (.Y(_09932_),
    .A(_09526_));
 sg13g2_nand2_1 _15867_ (.Y(_09933_),
    .A(_09140_),
    .B(_09520_));
 sg13g2_o21ai_1 _15868_ (.B1(_09933_),
    .Y(_09934_),
    .A1(net1018),
    .A2(_09526_));
 sg13g2_a22oi_1 _15869_ (.Y(_09935_),
    .B1(_09934_),
    .B2(net988),
    .A2(_09932_),
    .A1(net949));
 sg13g2_nand2_1 _15870_ (.Y(_09936_),
    .A(_07865_),
    .B(_07866_));
 sg13g2_a221oi_1 _15871_ (.B2(_09936_),
    .C1(_07872_),
    .B1(_07860_),
    .A1(_07544_),
    .Y(_09937_),
    .A2(_07541_));
 sg13g2_xnor2_1 _15872_ (.Y(_09938_),
    .A(_07549_),
    .B(_09937_));
 sg13g2_a221oi_1 _15873_ (.B2(net915),
    .C1(net989),
    .B1(_09938_),
    .A1(_09244_),
    .Y(_09939_),
    .A2(_09935_));
 sg13g2_a21oi_1 _15874_ (.A1(\top_ihp.oisc.decoder.instruction[29] ),
    .A2(net870),
    .Y(_09940_),
    .B1(_09939_));
 sg13g2_nand2_1 _15875_ (.Y(_09941_),
    .A(net886),
    .B(_09940_));
 sg13g2_o21ai_1 _15876_ (.B1(_09941_),
    .Y(_09942_),
    .A1(net1032),
    .A2(net871));
 sg13g2_buf_1 _15877_ (.A(_09942_),
    .X(_09943_));
 sg13g2_buf_2 _15878_ (.A(_09943_),
    .X(_09944_));
 sg13g2_nand2_1 _15879_ (.Y(_09945_),
    .A(\top_ihp.oisc.regs[0][9] ),
    .B(net550));
 sg13g2_o21ai_1 _15880_ (.B1(_09945_),
    .Y(_00389_),
    .A1(net549),
    .A2(net66));
 sg13g2_buf_2 _15881_ (.A(_09198_),
    .X(_09946_));
 sg13g2_nand2_1 _15882_ (.Y(_09947_),
    .A(net994),
    .B(_09207_));
 sg13g2_nand3_1 _15883_ (.B(net1019),
    .C(_09947_),
    .A(_08992_),
    .Y(_09948_));
 sg13g2_nand3_1 _15884_ (.B(_09102_),
    .C(_09948_),
    .A(_09083_),
    .Y(_09949_));
 sg13g2_buf_1 _15885_ (.A(_09949_),
    .X(_09950_));
 sg13g2_nor2_1 _15886_ (.A(_09054_),
    .B(_09097_),
    .Y(_09951_));
 sg13g2_a21oi_1 _15887_ (.A1(_09054_),
    .A2(_09947_),
    .Y(_09952_),
    .B1(_09951_));
 sg13g2_nor2_1 _15888_ (.A(_08943_),
    .B(_09952_),
    .Y(_09953_));
 sg13g2_nor2_1 _15889_ (.A(_08992_),
    .B(_09947_),
    .Y(_09954_));
 sg13g2_a21oi_1 _15890_ (.A1(_09950_),
    .A2(_09953_),
    .Y(_09955_),
    .B1(_09954_));
 sg13g2_buf_2 _15891_ (.A(_09955_),
    .X(_09956_));
 sg13g2_nand2b_1 _15892_ (.Y(_09957_),
    .B(_09083_),
    .A_N(_09956_));
 sg13g2_buf_2 _15893_ (.A(_09957_),
    .X(_09958_));
 sg13g2_and2_1 _15894_ (.A(_09080_),
    .B(_09073_),
    .X(_09959_));
 sg13g2_buf_1 _15895_ (.A(_09959_),
    .X(_09960_));
 sg13g2_nand2_1 _15896_ (.Y(_09961_),
    .A(_09095_),
    .B(net711));
 sg13g2_buf_2 _15897_ (.A(_09961_),
    .X(_09962_));
 sg13g2_or2_1 _15898_ (.X(_09963_),
    .B(_09962_),
    .A(_09958_));
 sg13g2_buf_1 _15899_ (.A(_09963_),
    .X(_09964_));
 sg13g2_buf_1 _15900_ (.A(_09964_),
    .X(_09965_));
 sg13g2_buf_1 _15901_ (.A(_09964_),
    .X(_09966_));
 sg13g2_nand2_1 _15902_ (.Y(_09967_),
    .A(_00141_),
    .B(net233));
 sg13g2_o21ai_1 _15903_ (.B1(_09967_),
    .Y(_00390_),
    .A1(net407),
    .A2(net234));
 sg13g2_nand2_1 _15904_ (.Y(_09968_),
    .A(\top_ihp.oisc.regs[10][10] ),
    .B(net233));
 sg13g2_o21ai_1 _15905_ (.B1(_09968_),
    .Y(_00391_),
    .A1(net74),
    .A2(net234));
 sg13g2_nand2_1 _15906_ (.Y(_09969_),
    .A(\top_ihp.oisc.regs[10][11] ),
    .B(net233));
 sg13g2_o21ai_1 _15907_ (.B1(_09969_),
    .Y(_00392_),
    .A1(net148),
    .A2(net234));
 sg13g2_nand2_1 _15908_ (.Y(_09970_),
    .A(\top_ihp.oisc.regs[10][12] ),
    .B(net233));
 sg13g2_o21ai_1 _15909_ (.B1(_09970_),
    .Y(_00393_),
    .A1(net250),
    .A2(net234));
 sg13g2_nand2_1 _15910_ (.Y(_09971_),
    .A(\top_ihp.oisc.regs[10][13] ),
    .B(_09966_));
 sg13g2_o21ai_1 _15911_ (.B1(_09971_),
    .Y(_00394_),
    .A1(net73),
    .A2(_09965_));
 sg13g2_nand2_1 _15912_ (.Y(_09972_),
    .A(\top_ihp.oisc.regs[10][14] ),
    .B(net233));
 sg13g2_o21ai_1 _15913_ (.B1(_09972_),
    .Y(_00395_),
    .A1(net249),
    .A2(net234));
 sg13g2_nand2_1 _15914_ (.Y(_09973_),
    .A(\top_ihp.oisc.regs[10][15] ),
    .B(net233));
 sg13g2_o21ai_1 _15915_ (.B1(_09973_),
    .Y(_00396_),
    .A1(net248),
    .A2(net234));
 sg13g2_nand2_1 _15916_ (.Y(_09974_),
    .A(\top_ihp.oisc.regs[10][16] ),
    .B(_09966_));
 sg13g2_o21ai_1 _15917_ (.B1(_09974_),
    .Y(_00397_),
    .A1(net146),
    .A2(_09965_));
 sg13g2_nand2_1 _15918_ (.Y(_09975_),
    .A(\top_ihp.oisc.regs[10][17] ),
    .B(net233));
 sg13g2_o21ai_1 _15919_ (.B1(_09975_),
    .Y(_00398_),
    .A1(net145),
    .A2(net234));
 sg13g2_nand2_1 _15920_ (.Y(_09976_),
    .A(\top_ihp.oisc.regs[10][18] ),
    .B(net233));
 sg13g2_o21ai_1 _15921_ (.B1(_09976_),
    .Y(_00399_),
    .A1(net144),
    .A2(net234));
 sg13g2_buf_1 _15922_ (.A(_09964_),
    .X(_09977_));
 sg13g2_buf_1 _15923_ (.A(_09964_),
    .X(_09978_));
 sg13g2_nand2_1 _15924_ (.Y(_09979_),
    .A(\top_ihp.oisc.regs[10][19] ),
    .B(net231));
 sg13g2_o21ai_1 _15925_ (.B1(_09979_),
    .Y(_00400_),
    .A1(net246),
    .A2(net232));
 sg13g2_nand2_1 _15926_ (.Y(_09980_),
    .A(\top_ihp.oisc.regs[10][1] ),
    .B(net231));
 sg13g2_o21ai_1 _15927_ (.B1(_09980_),
    .Y(_00401_),
    .A1(net409),
    .A2(net232));
 sg13g2_buf_8 _15928_ (.A(_09581_),
    .X(_09981_));
 sg13g2_nor2_1 _15929_ (.A(_09958_),
    .B(_09962_),
    .Y(_09982_));
 sg13g2_nor2_1 _15930_ (.A(\top_ihp.oisc.regs[10][20] ),
    .B(_09982_),
    .Y(_09983_));
 sg13g2_a21oi_1 _15931_ (.A1(net40),
    .A2(_09982_),
    .Y(_00402_),
    .B1(_09983_));
 sg13g2_nand2_1 _15932_ (.Y(_09984_),
    .A(\top_ihp.oisc.regs[10][21] ),
    .B(net231));
 sg13g2_o21ai_1 _15933_ (.B1(_09984_),
    .Y(_00403_),
    .A1(net72),
    .A2(net232));
 sg13g2_nand2_1 _15934_ (.Y(_09985_),
    .A(\top_ihp.oisc.regs[10][22] ),
    .B(net231));
 sg13g2_o21ai_1 _15935_ (.B1(_09985_),
    .Y(_00404_),
    .A1(net143),
    .A2(net232));
 sg13g2_buf_1 _15936_ (.A(net243),
    .X(_09986_));
 sg13g2_nor2_1 _15937_ (.A(\top_ihp.oisc.regs[10][23] ),
    .B(_09982_),
    .Y(_09987_));
 sg13g2_a21oi_1 _15938_ (.A1(net138),
    .A2(_09982_),
    .Y(_00405_),
    .B1(_09987_));
 sg13g2_nand2_1 _15939_ (.Y(_09988_),
    .A(\top_ihp.oisc.regs[10][24] ),
    .B(net231));
 sg13g2_o21ai_1 _15940_ (.B1(_09988_),
    .Y(_00406_),
    .A1(net242),
    .A2(net232));
 sg13g2_nand2_1 _15941_ (.Y(_09989_),
    .A(\top_ihp.oisc.regs[10][25] ),
    .B(net231));
 sg13g2_o21ai_1 _15942_ (.B1(_09989_),
    .Y(_00407_),
    .A1(net241),
    .A2(_09977_));
 sg13g2_nand2_1 _15943_ (.Y(_09990_),
    .A(\top_ihp.oisc.regs[10][26] ),
    .B(_09978_));
 sg13g2_o21ai_1 _15944_ (.B1(_09990_),
    .Y(_00408_),
    .A1(net142),
    .A2(_09977_));
 sg13g2_nand2_1 _15945_ (.Y(_09991_),
    .A(\top_ihp.oisc.regs[10][27] ),
    .B(net231));
 sg13g2_o21ai_1 _15946_ (.B1(_09991_),
    .Y(_00409_),
    .A1(net71),
    .A2(net232));
 sg13g2_nand2_1 _15947_ (.Y(_09992_),
    .A(\top_ihp.oisc.regs[10][28] ),
    .B(net231));
 sg13g2_o21ai_1 _15948_ (.B1(_09992_),
    .Y(_00410_),
    .A1(net70),
    .A2(net232));
 sg13g2_nand2_1 _15949_ (.Y(_09993_),
    .A(\top_ihp.oisc.regs[10][29] ),
    .B(_09978_));
 sg13g2_o21ai_1 _15950_ (.B1(_09993_),
    .Y(_00411_),
    .A1(net140),
    .A2(net232));
 sg13g2_buf_1 _15951_ (.A(_09964_),
    .X(_09994_));
 sg13g2_buf_1 _15952_ (.A(_09964_),
    .X(_09995_));
 sg13g2_nand2_1 _15953_ (.Y(_09996_),
    .A(\top_ihp.oisc.regs[10][2] ),
    .B(net229));
 sg13g2_o21ai_1 _15954_ (.B1(_09996_),
    .Y(_00412_),
    .A1(net240),
    .A2(net230));
 sg13g2_nand2_1 _15955_ (.Y(_09997_),
    .A(\top_ihp.oisc.regs[10][30] ),
    .B(_09995_));
 sg13g2_o21ai_1 _15956_ (.B1(_09997_),
    .Y(_00413_),
    .A1(net69),
    .A2(_09994_));
 sg13g2_nand2_1 _15957_ (.Y(_09998_),
    .A(\top_ihp.oisc.regs[10][31] ),
    .B(_09995_));
 sg13g2_o21ai_1 _15958_ (.B1(_09998_),
    .Y(_00414_),
    .A1(net139),
    .A2(_09994_));
 sg13g2_nand2_1 _15959_ (.Y(_09999_),
    .A(\top_ihp.oisc.regs[10][3] ),
    .B(net229));
 sg13g2_o21ai_1 _15960_ (.B1(_09999_),
    .Y(_00415_),
    .A1(net238),
    .A2(net230));
 sg13g2_nand2_1 _15961_ (.Y(_10000_),
    .A(\top_ihp.oisc.regs[10][4] ),
    .B(net229));
 sg13g2_o21ai_1 _15962_ (.B1(_10000_),
    .Y(_00416_),
    .A1(net237),
    .A2(net230));
 sg13g2_nand2_1 _15963_ (.Y(_10001_),
    .A(\top_ihp.oisc.regs[10][5] ),
    .B(net229));
 sg13g2_o21ai_1 _15964_ (.B1(_10001_),
    .Y(_00417_),
    .A1(net236),
    .A2(net230));
 sg13g2_nand2_1 _15965_ (.Y(_10002_),
    .A(\top_ihp.oisc.regs[10][6] ),
    .B(net229));
 sg13g2_o21ai_1 _15966_ (.B1(_10002_),
    .Y(_00418_),
    .A1(net235),
    .A2(net230));
 sg13g2_nand2_1 _15967_ (.Y(_10003_),
    .A(\top_ihp.oisc.regs[10][7] ),
    .B(net229));
 sg13g2_o21ai_1 _15968_ (.B1(_10003_),
    .Y(_00419_),
    .A1(net68),
    .A2(net230));
 sg13g2_nand2_1 _15969_ (.Y(_10004_),
    .A(\top_ihp.oisc.regs[10][8] ),
    .B(net229));
 sg13g2_o21ai_1 _15970_ (.B1(_10004_),
    .Y(_00420_),
    .A1(net67),
    .A2(net230));
 sg13g2_nand2_1 _15971_ (.Y(_10005_),
    .A(\top_ihp.oisc.regs[10][9] ),
    .B(net229));
 sg13g2_o21ai_1 _15972_ (.B1(_10005_),
    .Y(_00421_),
    .A1(net66),
    .A2(net230));
 sg13g2_nor2b_1 _15973_ (.A(_09956_),
    .B_N(_09083_),
    .Y(_10006_));
 sg13g2_buf_2 _15974_ (.A(_10006_),
    .X(_10007_));
 sg13g2_nor2_1 _15975_ (.A(_09080_),
    .B(_09069_),
    .Y(_10008_));
 sg13g2_buf_2 _15976_ (.A(_10008_),
    .X(_10009_));
 sg13g2_and2_1 _15977_ (.A(_09095_),
    .B(_10009_),
    .X(_10010_));
 sg13g2_buf_1 _15978_ (.A(_10010_),
    .X(_10011_));
 sg13g2_nand2_1 _15979_ (.Y(_10012_),
    .A(_10007_),
    .B(_10011_));
 sg13g2_buf_2 _15980_ (.A(_10012_),
    .X(_10013_));
 sg13g2_buf_1 _15981_ (.A(_10013_),
    .X(_10014_));
 sg13g2_buf_1 _15982_ (.A(_10013_),
    .X(_10015_));
 sg13g2_nand2_1 _15983_ (.Y(_10016_),
    .A(_00142_),
    .B(net227));
 sg13g2_o21ai_1 _15984_ (.B1(_10016_),
    .Y(_00422_),
    .A1(net407),
    .A2(net228));
 sg13g2_nand2_1 _15985_ (.Y(_10017_),
    .A(\top_ihp.oisc.regs[11][10] ),
    .B(net227));
 sg13g2_o21ai_1 _15986_ (.B1(_10017_),
    .Y(_00423_),
    .A1(net74),
    .A2(net228));
 sg13g2_nand2_1 _15987_ (.Y(_10018_),
    .A(\top_ihp.oisc.regs[11][11] ),
    .B(net227));
 sg13g2_o21ai_1 _15988_ (.B1(_10018_),
    .Y(_00424_),
    .A1(net148),
    .A2(net228));
 sg13g2_nand2_1 _15989_ (.Y(_10019_),
    .A(\top_ihp.oisc.regs[11][12] ),
    .B(net227));
 sg13g2_o21ai_1 _15990_ (.B1(_10019_),
    .Y(_00425_),
    .A1(net250),
    .A2(net228));
 sg13g2_buf_1 _15991_ (.A(_10013_),
    .X(_10020_));
 sg13g2_nand2_1 _15992_ (.Y(_10021_),
    .A(\top_ihp.oisc.regs[11][13] ),
    .B(net226));
 sg13g2_o21ai_1 _15993_ (.B1(_10021_),
    .Y(_00426_),
    .A1(net73),
    .A2(_10014_));
 sg13g2_nand2_1 _15994_ (.Y(_10022_),
    .A(\top_ihp.oisc.regs[11][14] ),
    .B(net226));
 sg13g2_o21ai_1 _15995_ (.B1(_10022_),
    .Y(_00427_),
    .A1(net249),
    .A2(net228));
 sg13g2_nand2_1 _15996_ (.Y(_10023_),
    .A(\top_ihp.oisc.regs[11][15] ),
    .B(net226));
 sg13g2_o21ai_1 _15997_ (.B1(_10023_),
    .Y(_00428_),
    .A1(net248),
    .A2(net228));
 sg13g2_nand2_1 _15998_ (.Y(_10024_),
    .A(\top_ihp.oisc.regs[11][16] ),
    .B(net226));
 sg13g2_o21ai_1 _15999_ (.B1(_10024_),
    .Y(_00429_),
    .A1(net146),
    .A2(_10014_));
 sg13g2_nand2_1 _16000_ (.Y(_10025_),
    .A(\top_ihp.oisc.regs[11][17] ),
    .B(net226));
 sg13g2_o21ai_1 _16001_ (.B1(_10025_),
    .Y(_00430_),
    .A1(net145),
    .A2(net228));
 sg13g2_nand2_1 _16002_ (.Y(_10026_),
    .A(\top_ihp.oisc.regs[11][18] ),
    .B(net226));
 sg13g2_o21ai_1 _16003_ (.B1(_10026_),
    .Y(_00431_),
    .A1(net144),
    .A2(net228));
 sg13g2_buf_1 _16004_ (.A(_10013_),
    .X(_10027_));
 sg13g2_nand2_1 _16005_ (.Y(_10028_),
    .A(\top_ihp.oisc.regs[11][19] ),
    .B(net226));
 sg13g2_o21ai_1 _16006_ (.B1(_10028_),
    .Y(_00432_),
    .A1(net246),
    .A2(net225));
 sg13g2_buf_1 _16007_ (.A(_10007_),
    .X(_10029_));
 sg13g2_and2_1 _16008_ (.A(net545),
    .B(_10011_),
    .X(_10030_));
 sg13g2_buf_2 _16009_ (.A(_10030_),
    .X(_10031_));
 sg13g2_mux2_1 _16010_ (.A0(_00143_),
    .A1(net547),
    .S(_10031_),
    .X(_00433_));
 sg13g2_buf_2 _16011_ (.A(net245),
    .X(_10032_));
 sg13g2_mux2_1 _16012_ (.A0(\top_ihp.oisc.regs[11][20] ),
    .A1(net137),
    .S(_10031_),
    .X(_00434_));
 sg13g2_nand2_1 _16013_ (.Y(_10033_),
    .A(\top_ihp.oisc.regs[11][21] ),
    .B(net226));
 sg13g2_o21ai_1 _16014_ (.B1(_10033_),
    .Y(_00435_),
    .A1(net72),
    .A2(net225));
 sg13g2_nand2_1 _16015_ (.Y(_10034_),
    .A(\top_ihp.oisc.regs[11][22] ),
    .B(_10020_));
 sg13g2_o21ai_1 _16016_ (.B1(_10034_),
    .Y(_00436_),
    .A1(net143),
    .A2(net225));
 sg13g2_buf_1 _16017_ (.A(_09641_),
    .X(_10035_));
 sg13g2_buf_1 _16018_ (.A(net406),
    .X(_10036_));
 sg13g2_mux2_1 _16019_ (.A0(\top_ihp.oisc.regs[11][23] ),
    .A1(net224),
    .S(_10031_),
    .X(_00437_));
 sg13g2_nand2_1 _16020_ (.Y(_10037_),
    .A(\top_ihp.oisc.regs[11][24] ),
    .B(_10020_));
 sg13g2_o21ai_1 _16021_ (.B1(_10037_),
    .Y(_00438_),
    .A1(net242),
    .A2(net225));
 sg13g2_buf_1 _16022_ (.A(_10013_),
    .X(_10038_));
 sg13g2_nand2_1 _16023_ (.Y(_10039_),
    .A(\top_ihp.oisc.regs[11][25] ),
    .B(net223));
 sg13g2_o21ai_1 _16024_ (.B1(_10039_),
    .Y(_00439_),
    .A1(net241),
    .A2(net225));
 sg13g2_nand2_1 _16025_ (.Y(_10040_),
    .A(\top_ihp.oisc.regs[11][26] ),
    .B(net223));
 sg13g2_o21ai_1 _16026_ (.B1(_10040_),
    .Y(_00440_),
    .A1(net142),
    .A2(net225));
 sg13g2_nand2_1 _16027_ (.Y(_10041_),
    .A(\top_ihp.oisc.regs[11][27] ),
    .B(net223));
 sg13g2_o21ai_1 _16028_ (.B1(_10041_),
    .Y(_00441_),
    .A1(net71),
    .A2(net225));
 sg13g2_nand2_1 _16029_ (.Y(_10042_),
    .A(\top_ihp.oisc.regs[11][28] ),
    .B(net223));
 sg13g2_o21ai_1 _16030_ (.B1(_10042_),
    .Y(_00442_),
    .A1(net70),
    .A2(_10027_));
 sg13g2_nand2_1 _16031_ (.Y(_10043_),
    .A(\top_ihp.oisc.regs[11][29] ),
    .B(_10038_));
 sg13g2_o21ai_1 _16032_ (.B1(_10043_),
    .Y(_00443_),
    .A1(net140),
    .A2(_10027_));
 sg13g2_buf_1 _16033_ (.A(_09753_),
    .X(_10044_));
 sg13g2_mux2_1 _16034_ (.A0(_00144_),
    .A1(net222),
    .S(_10031_),
    .X(_00444_));
 sg13g2_nand2_1 _16035_ (.Y(_10045_),
    .A(\top_ihp.oisc.regs[11][30] ),
    .B(_10038_));
 sg13g2_o21ai_1 _16036_ (.B1(_10045_),
    .Y(_00445_),
    .A1(net69),
    .A2(net225));
 sg13g2_nand2_1 _16037_ (.Y(_10046_),
    .A(\top_ihp.oisc.regs[11][31] ),
    .B(net223));
 sg13g2_o21ai_1 _16038_ (.B1(_10046_),
    .Y(_00446_),
    .A1(net139),
    .A2(_10015_));
 sg13g2_buf_1 _16039_ (.A(_09807_),
    .X(_10047_));
 sg13g2_mux2_1 _16040_ (.A0(_00145_),
    .A1(net221),
    .S(_10031_),
    .X(_00447_));
 sg13g2_buf_1 _16041_ (.A(_09840_),
    .X(_10048_));
 sg13g2_mux2_1 _16042_ (.A0(_00146_),
    .A1(net220),
    .S(_10031_),
    .X(_00448_));
 sg13g2_nand2_1 _16043_ (.Y(_10049_),
    .A(\top_ihp.oisc.regs[11][5] ),
    .B(net223));
 sg13g2_o21ai_1 _16044_ (.B1(_10049_),
    .Y(_00449_),
    .A1(net236),
    .A2(_10015_));
 sg13g2_nand2_1 _16045_ (.Y(_10050_),
    .A(\top_ihp.oisc.regs[11][6] ),
    .B(net223));
 sg13g2_o21ai_1 _16046_ (.B1(_10050_),
    .Y(_00450_),
    .A1(net235),
    .A2(net227));
 sg13g2_nand2_1 _16047_ (.Y(_10051_),
    .A(\top_ihp.oisc.regs[11][7] ),
    .B(net223));
 sg13g2_o21ai_1 _16048_ (.B1(_10051_),
    .Y(_00451_),
    .A1(net68),
    .A2(net227));
 sg13g2_nand2_1 _16049_ (.Y(_10052_),
    .A(\top_ihp.oisc.regs[11][8] ),
    .B(_10013_));
 sg13g2_o21ai_1 _16050_ (.B1(_10052_),
    .Y(_00452_),
    .A1(net67),
    .A2(net227));
 sg13g2_nand2_1 _16051_ (.Y(_10053_),
    .A(\top_ihp.oisc.regs[11][9] ),
    .B(_10013_));
 sg13g2_o21ai_1 _16052_ (.B1(_10053_),
    .Y(_00453_),
    .A1(net66),
    .A2(net227));
 sg13g2_nor3_1 _16053_ (.A(_08943_),
    .B(_09950_),
    .C(_09952_),
    .Y(_10054_));
 sg13g2_buf_2 _16054_ (.A(_10054_),
    .X(_10055_));
 sg13g2_nor2b_1 _16055_ (.A(_09082_),
    .B_N(_09095_),
    .Y(_10056_));
 sg13g2_buf_2 _16056_ (.A(_10056_),
    .X(_10057_));
 sg13g2_nand2_1 _16057_ (.Y(_10058_),
    .A(_10055_),
    .B(_10057_));
 sg13g2_buf_1 _16058_ (.A(_10058_),
    .X(_10059_));
 sg13g2_buf_1 _16059_ (.A(_10059_),
    .X(_10060_));
 sg13g2_buf_1 _16060_ (.A(net405),
    .X(_10061_));
 sg13g2_nand2_1 _16061_ (.Y(_10062_),
    .A(_00147_),
    .B(net405));
 sg13g2_o21ai_1 _16062_ (.B1(_10062_),
    .Y(_00454_),
    .A1(net407),
    .A2(net219));
 sg13g2_buf_8 _16063_ (.A(_09269_),
    .X(_10063_));
 sg13g2_mux2_1 _16064_ (.A0(net65),
    .A1(_00148_),
    .S(net219),
    .X(_00455_));
 sg13g2_mux2_1 _16065_ (.A0(net251),
    .A1(_00149_),
    .S(net219),
    .X(_00456_));
 sg13g2_buf_8 _16066_ (.A(_09347_),
    .X(_10064_));
 sg13g2_mux2_1 _16067_ (.A0(_10064_),
    .A1(_00150_),
    .S(net219),
    .X(_00457_));
 sg13g2_nand2_1 _16068_ (.Y(_10065_),
    .A(_00151_),
    .B(net405));
 sg13g2_o21ai_1 _16069_ (.B1(_10065_),
    .Y(_00458_),
    .A1(_09372_),
    .A2(net219));
 sg13g2_buf_1 _16070_ (.A(_09403_),
    .X(_10066_));
 sg13g2_buf_2 _16071_ (.A(_10059_),
    .X(_10067_));
 sg13g2_mux2_1 _16072_ (.A0(net217),
    .A1(_00152_),
    .S(net404),
    .X(_00459_));
 sg13g2_buf_1 _16073_ (.A(_09418_),
    .X(_10068_));
 sg13g2_mux2_1 _16074_ (.A0(net216),
    .A1(_00153_),
    .S(net404),
    .X(_00460_));
 sg13g2_nand2_1 _16075_ (.Y(_10069_),
    .A(_00154_),
    .B(net405));
 sg13g2_o21ai_1 _16076_ (.B1(_10069_),
    .Y(_00461_),
    .A1(_09434_),
    .A2(net219));
 sg13g2_buf_1 _16077_ (.A(_09461_),
    .X(_10070_));
 sg13g2_mux2_1 _16078_ (.A0(net136),
    .A1(_00155_),
    .S(net404),
    .X(_00462_));
 sg13g2_buf_1 _16079_ (.A(_09482_),
    .X(_10071_));
 sg13g2_mux2_1 _16080_ (.A0(net135),
    .A1(_00156_),
    .S(net404),
    .X(_00463_));
 sg13g2_buf_1 _16081_ (.A(_09511_),
    .X(_10072_));
 sg13g2_mux2_1 _16082_ (.A0(net215),
    .A1(_00157_),
    .S(net404),
    .X(_00464_));
 sg13g2_mux2_1 _16083_ (.A0(_09553_),
    .A1(_00158_),
    .S(net404),
    .X(_00465_));
 sg13g2_nand2_1 _16084_ (.Y(_10073_),
    .A(_00159_),
    .B(net405));
 sg13g2_o21ai_1 _16085_ (.B1(_10073_),
    .Y(_00466_),
    .A1(net137),
    .A2(net219));
 sg13g2_buf_8 _16086_ (.A(_09598_),
    .X(_10074_));
 sg13g2_mux2_1 _16087_ (.A0(_10074_),
    .A1(_00160_),
    .S(_10067_),
    .X(_00467_));
 sg13g2_nand2_1 _16088_ (.Y(_10075_),
    .A(_00161_),
    .B(_10060_));
 sg13g2_o21ai_1 _16089_ (.B1(_10075_),
    .Y(_00468_),
    .A1(_09620_),
    .A2(_10061_));
 sg13g2_nand2_1 _16090_ (.Y(_10076_),
    .A(_00162_),
    .B(net405));
 sg13g2_o21ai_1 _16091_ (.B1(_10076_),
    .Y(_00469_),
    .A1(net224),
    .A2(net219));
 sg13g2_buf_2 _16092_ (.A(_09653_),
    .X(_10077_));
 sg13g2_mux2_1 _16093_ (.A0(net214),
    .A1(_00163_),
    .S(net404),
    .X(_00470_));
 sg13g2_buf_1 _16094_ (.A(_09668_),
    .X(_10078_));
 sg13g2_mux2_1 _16095_ (.A0(net213),
    .A1(_00164_),
    .S(_10067_),
    .X(_00471_));
 sg13g2_buf_8 _16096_ (.A(_09678_),
    .X(_10079_));
 sg13g2_mux2_1 _16097_ (.A0(net134),
    .A1(_00165_),
    .S(net404),
    .X(_00472_));
 sg13g2_nand2_1 _16098_ (.Y(_10080_),
    .A(_00166_),
    .B(_10060_));
 sg13g2_o21ai_1 _16099_ (.B1(_10080_),
    .Y(_00473_),
    .A1(_09699_),
    .A2(_10061_));
 sg13g2_buf_8 _16100_ (.A(_09713_),
    .X(_10081_));
 sg13g2_buf_2 _16101_ (.A(_10059_),
    .X(_10082_));
 sg13g2_mux2_1 _16102_ (.A0(net63),
    .A1(_00167_),
    .S(net403),
    .X(_00474_));
 sg13g2_buf_1 _16103_ (.A(_09723_),
    .X(_10083_));
 sg13g2_mux2_1 _16104_ (.A0(net133),
    .A1(_00168_),
    .S(_10082_),
    .X(_00475_));
 sg13g2_mux2_1 _16105_ (.A0(net222),
    .A1(_00169_),
    .S(net403),
    .X(_00476_));
 sg13g2_buf_8 _16106_ (.A(_09761_),
    .X(_10084_));
 sg13g2_mux2_1 _16107_ (.A0(net62),
    .A1(_00170_),
    .S(_10082_),
    .X(_00477_));
 sg13g2_mux2_1 _16108_ (.A0(net239),
    .A1(_00171_),
    .S(net403),
    .X(_00478_));
 sg13g2_mux2_1 _16109_ (.A0(net221),
    .A1(_00172_),
    .S(net403),
    .X(_00479_));
 sg13g2_mux2_1 _16110_ (.A0(net220),
    .A1(_00173_),
    .S(net403),
    .X(_00480_));
 sg13g2_buf_2 _16111_ (.A(_09871_),
    .X(_10085_));
 sg13g2_mux2_1 _16112_ (.A0(net212),
    .A1(_00174_),
    .S(net403),
    .X(_00481_));
 sg13g2_buf_2 _16113_ (.A(_09894_),
    .X(_10086_));
 sg13g2_mux2_1 _16114_ (.A0(net211),
    .A1(_00175_),
    .S(net403),
    .X(_00482_));
 sg13g2_mux2_1 _16115_ (.A0(net408),
    .A1(_00176_),
    .S(net403),
    .X(_00483_));
 sg13g2_buf_8 _16116_ (.A(_09929_),
    .X(_10087_));
 sg13g2_mux2_1 _16117_ (.A0(net61),
    .A1(_00177_),
    .S(net405),
    .X(_00484_));
 sg13g2_buf_8 _16118_ (.A(_09943_),
    .X(_10088_));
 sg13g2_mux2_1 _16119_ (.A0(net60),
    .A1(_00178_),
    .S(net405),
    .X(_00485_));
 sg13g2_nand2b_1 _16120_ (.Y(_10089_),
    .B(_09953_),
    .A_N(_09950_));
 sg13g2_buf_2 _16121_ (.A(_10089_),
    .X(_10090_));
 sg13g2_nor2b_1 _16122_ (.A(_09080_),
    .B_N(_09069_),
    .Y(_10091_));
 sg13g2_buf_2 _16123_ (.A(_10091_),
    .X(_10092_));
 sg13g2_nand2_2 _16124_ (.Y(_10093_),
    .A(_09095_),
    .B(net710));
 sg13g2_nor2_1 _16125_ (.A(_10090_),
    .B(_10093_),
    .Y(_10094_));
 sg13g2_buf_1 _16126_ (.A(_10094_),
    .X(_10095_));
 sg13g2_buf_1 _16127_ (.A(_10095_),
    .X(_10096_));
 sg13g2_buf_2 _16128_ (.A(net544),
    .X(_10097_));
 sg13g2_mux2_1 _16129_ (.A0(\top_ihp.oisc.regs[13][0] ),
    .A1(net407),
    .S(net402),
    .X(_00486_));
 sg13g2_nor2_1 _16130_ (.A(_00179_),
    .B(net544),
    .Y(_10098_));
 sg13g2_a21oi_1 _16131_ (.A1(_09267_),
    .A2(net402),
    .Y(_00487_),
    .B1(_10098_));
 sg13g2_nor2_1 _16132_ (.A(_00180_),
    .B(net544),
    .Y(_10099_));
 sg13g2_a21oi_1 _16133_ (.A1(_09301_),
    .A2(net402),
    .Y(_00488_),
    .B1(_10099_));
 sg13g2_mux2_1 _16134_ (.A0(_00181_),
    .A1(net218),
    .S(net402),
    .X(_00489_));
 sg13g2_mux2_1 _16135_ (.A0(_00182_),
    .A1(net147),
    .S(_10097_),
    .X(_00490_));
 sg13g2_buf_2 _16136_ (.A(_10095_),
    .X(_10100_));
 sg13g2_mux2_1 _16137_ (.A0(_00183_),
    .A1(net217),
    .S(net543),
    .X(_00491_));
 sg13g2_mux2_1 _16138_ (.A0(_00184_),
    .A1(net216),
    .S(net543),
    .X(_00492_));
 sg13g2_mux2_1 _16139_ (.A0(_00185_),
    .A1(net247),
    .S(_10100_),
    .X(_00493_));
 sg13g2_mux2_1 _16140_ (.A0(_00186_),
    .A1(net136),
    .S(net543),
    .X(_00494_));
 sg13g2_mux2_1 _16141_ (.A0(_00187_),
    .A1(net135),
    .S(net543),
    .X(_00495_));
 sg13g2_mux2_1 _16142_ (.A0(_00188_),
    .A1(net215),
    .S(net543),
    .X(_00496_));
 sg13g2_nor2_1 _16143_ (.A(\top_ihp.oisc.regs[13][1] ),
    .B(_10096_),
    .Y(_10101_));
 sg13g2_a21oi_1 _16144_ (.A1(net409),
    .A2(net402),
    .Y(_00497_),
    .B1(_10101_));
 sg13g2_mux2_1 _16145_ (.A0(_00189_),
    .A1(_09563_),
    .S(net543),
    .X(_00498_));
 sg13g2_mux2_1 _16146_ (.A0(_00190_),
    .A1(_10074_),
    .S(_10100_),
    .X(_00499_));
 sg13g2_mux2_1 _16147_ (.A0(_00191_),
    .A1(net244),
    .S(net543),
    .X(_00500_));
 sg13g2_mux2_1 _16148_ (.A0(_00192_),
    .A1(net243),
    .S(net543),
    .X(_00501_));
 sg13g2_nor2_1 _16149_ (.A(_00193_),
    .B(_10096_),
    .Y(_10102_));
 sg13g2_a21oi_1 _16150_ (.A1(_09651_),
    .A2(_10097_),
    .Y(_00502_),
    .B1(_10102_));
 sg13g2_buf_2 _16151_ (.A(_10095_),
    .X(_10103_));
 sg13g2_mux2_1 _16152_ (.A0(_00194_),
    .A1(net213),
    .S(net542),
    .X(_00503_));
 sg13g2_mux2_1 _16153_ (.A0(_00195_),
    .A1(net134),
    .S(net542),
    .X(_00504_));
 sg13g2_mux2_1 _16154_ (.A0(_00196_),
    .A1(net141),
    .S(net542),
    .X(_00505_));
 sg13g2_mux2_1 _16155_ (.A0(_00197_),
    .A1(net63),
    .S(net542),
    .X(_00506_));
 sg13g2_mux2_1 _16156_ (.A0(_00198_),
    .A1(net133),
    .S(_10103_),
    .X(_00507_));
 sg13g2_mux2_1 _16157_ (.A0(_00199_),
    .A1(net222),
    .S(net542),
    .X(_00508_));
 sg13g2_mux2_1 _16158_ (.A0(_00200_),
    .A1(net62),
    .S(_10103_),
    .X(_00509_));
 sg13g2_nor2_1 _16159_ (.A(_00201_),
    .B(net544),
    .Y(_10104_));
 sg13g2_a21oi_1 _16160_ (.A1(_09773_),
    .A2(net402),
    .Y(_00510_),
    .B1(_10104_));
 sg13g2_mux2_1 _16161_ (.A0(_00202_),
    .A1(net221),
    .S(net542),
    .X(_00511_));
 sg13g2_nor2_1 _16162_ (.A(_00203_),
    .B(net544),
    .Y(_10105_));
 sg13g2_a21oi_1 _16163_ (.A1(_09838_),
    .A2(net402),
    .Y(_00512_),
    .B1(_10105_));
 sg13g2_mux2_1 _16164_ (.A0(_00204_),
    .A1(net212),
    .S(net542),
    .X(_00513_));
 sg13g2_mux2_1 _16165_ (.A0(_00205_),
    .A1(net211),
    .S(net542),
    .X(_00514_));
 sg13g2_mux2_1 _16166_ (.A0(_00206_),
    .A1(net408),
    .S(net544),
    .X(_00515_));
 sg13g2_mux2_1 _16167_ (.A0(_00207_),
    .A1(net61),
    .S(net544),
    .X(_00516_));
 sg13g2_nor2_1 _16168_ (.A(_00208_),
    .B(net544),
    .Y(_10106_));
 sg13g2_a21oi_1 _16169_ (.A1(_09941_),
    .A2(net402),
    .Y(_00517_),
    .B1(_10106_));
 sg13g2_buf_2 _16170_ (.A(net412),
    .X(_10107_));
 sg13g2_nor2_1 _16171_ (.A(_09962_),
    .B(_10090_),
    .Y(_10108_));
 sg13g2_buf_1 _16172_ (.A(_10108_),
    .X(_10109_));
 sg13g2_mux2_1 _16173_ (.A0(\top_ihp.oisc.regs[14][0] ),
    .A1(net210),
    .S(net541),
    .X(_00518_));
 sg13g2_nand3_1 _16174_ (.B(net711),
    .C(_10055_),
    .A(_09095_),
    .Y(_10110_));
 sg13g2_buf_2 _16175_ (.A(_10110_),
    .X(_10111_));
 sg13g2_buf_1 _16176_ (.A(_10111_),
    .X(_10112_));
 sg13g2_buf_1 _16177_ (.A(_10111_),
    .X(_10113_));
 sg13g2_nand2_1 _16178_ (.Y(_10114_),
    .A(\top_ihp.oisc.regs[14][10] ),
    .B(net539));
 sg13g2_o21ai_1 _16179_ (.B1(_10114_),
    .Y(_00519_),
    .A1(net74),
    .A2(net540));
 sg13g2_nand2_1 _16180_ (.Y(_10115_),
    .A(\top_ihp.oisc.regs[14][11] ),
    .B(_10113_));
 sg13g2_o21ai_1 _16181_ (.B1(_10115_),
    .Y(_00520_),
    .A1(net148),
    .A2(net540));
 sg13g2_nand2_1 _16182_ (.Y(_10116_),
    .A(\top_ihp.oisc.regs[14][12] ),
    .B(net539));
 sg13g2_o21ai_1 _16183_ (.B1(_10116_),
    .Y(_00521_),
    .A1(net250),
    .A2(net540));
 sg13g2_buf_8 _16184_ (.A(net147),
    .X(_10117_));
 sg13g2_nor2_1 _16185_ (.A(\top_ihp.oisc.regs[14][13] ),
    .B(net541),
    .Y(_10118_));
 sg13g2_a21oi_1 _16186_ (.A1(net59),
    .A2(_10109_),
    .Y(_00522_),
    .B1(_10118_));
 sg13g2_nand2_1 _16187_ (.Y(_10119_),
    .A(\top_ihp.oisc.regs[14][14] ),
    .B(_10113_));
 sg13g2_o21ai_1 _16188_ (.B1(_10119_),
    .Y(_00523_),
    .A1(net249),
    .A2(net540));
 sg13g2_buf_1 _16189_ (.A(_10111_),
    .X(_10120_));
 sg13g2_nand2_1 _16190_ (.Y(_10121_),
    .A(\top_ihp.oisc.regs[14][15] ),
    .B(net538));
 sg13g2_o21ai_1 _16191_ (.B1(_10121_),
    .Y(_00524_),
    .A1(net248),
    .A2(net540));
 sg13g2_buf_8 _16192_ (.A(_09436_),
    .X(_10122_));
 sg13g2_nor2_1 _16193_ (.A(\top_ihp.oisc.regs[14][16] ),
    .B(_10109_),
    .Y(_10123_));
 sg13g2_a21oi_1 _16194_ (.A1(_10122_),
    .A2(net541),
    .Y(_00525_),
    .B1(_10123_));
 sg13g2_nand2_1 _16195_ (.Y(_10124_),
    .A(\top_ihp.oisc.regs[14][17] ),
    .B(net538));
 sg13g2_o21ai_1 _16196_ (.B1(_10124_),
    .Y(_00526_),
    .A1(net145),
    .A2(net540));
 sg13g2_nand2_1 _16197_ (.Y(_10125_),
    .A(\top_ihp.oisc.regs[14][18] ),
    .B(net538));
 sg13g2_o21ai_1 _16198_ (.B1(_10125_),
    .Y(_00527_),
    .A1(net144),
    .A2(net540));
 sg13g2_nand2_1 _16199_ (.Y(_10126_),
    .A(\top_ihp.oisc.regs[14][19] ),
    .B(net538));
 sg13g2_o21ai_1 _16200_ (.B1(_10126_),
    .Y(_00528_),
    .A1(net246),
    .A2(net540));
 sg13g2_nand2_1 _16201_ (.Y(_10127_),
    .A(\top_ihp.oisc.regs[14][1] ),
    .B(net538));
 sg13g2_o21ai_1 _16202_ (.B1(_10127_),
    .Y(_00529_),
    .A1(net409),
    .A2(_10112_));
 sg13g2_nor2_1 _16203_ (.A(\top_ihp.oisc.regs[14][20] ),
    .B(net541),
    .Y(_10128_));
 sg13g2_a21oi_1 _16204_ (.A1(net40),
    .A2(net541),
    .Y(_00530_),
    .B1(_10128_));
 sg13g2_nand2_1 _16205_ (.Y(_10129_),
    .A(\top_ihp.oisc.regs[14][21] ),
    .B(net538));
 sg13g2_o21ai_1 _16206_ (.B1(_10129_),
    .Y(_00531_),
    .A1(net72),
    .A2(_10112_));
 sg13g2_buf_1 _16207_ (.A(net244),
    .X(_10130_));
 sg13g2_nor2_1 _16208_ (.A(\top_ihp.oisc.regs[14][22] ),
    .B(net541),
    .Y(_10131_));
 sg13g2_a21oi_1 _16209_ (.A1(net131),
    .A2(net541),
    .Y(_00532_),
    .B1(_10131_));
 sg13g2_nor2_1 _16210_ (.A(\top_ihp.oisc.regs[14][23] ),
    .B(_10108_),
    .Y(_10132_));
 sg13g2_a21oi_1 _16211_ (.A1(_09986_),
    .A2(net541),
    .Y(_00533_),
    .B1(_10132_));
 sg13g2_buf_1 _16212_ (.A(_10111_),
    .X(_10133_));
 sg13g2_nand2_1 _16213_ (.Y(_10134_),
    .A(\top_ihp.oisc.regs[14][24] ),
    .B(net538));
 sg13g2_o21ai_1 _16214_ (.B1(_10134_),
    .Y(_00534_),
    .A1(net242),
    .A2(net537));
 sg13g2_nand2_1 _16215_ (.Y(_10135_),
    .A(\top_ihp.oisc.regs[14][25] ),
    .B(net538));
 sg13g2_o21ai_1 _16216_ (.B1(_10135_),
    .Y(_00535_),
    .A1(net241),
    .A2(net537));
 sg13g2_nand2_1 _16217_ (.Y(_10136_),
    .A(\top_ihp.oisc.regs[14][26] ),
    .B(_10120_));
 sg13g2_o21ai_1 _16218_ (.B1(_10136_),
    .Y(_00536_),
    .A1(net142),
    .A2(net537));
 sg13g2_nand2_1 _16219_ (.Y(_10137_),
    .A(\top_ihp.oisc.regs[14][27] ),
    .B(_10120_));
 sg13g2_o21ai_1 _16220_ (.B1(_10137_),
    .Y(_00537_),
    .A1(net71),
    .A2(net537));
 sg13g2_buf_1 _16221_ (.A(_10111_),
    .X(_10138_));
 sg13g2_nand2_1 _16222_ (.Y(_10139_),
    .A(\top_ihp.oisc.regs[14][28] ),
    .B(net536));
 sg13g2_o21ai_1 _16223_ (.B1(_10139_),
    .Y(_00538_),
    .A1(net70),
    .A2(net537));
 sg13g2_nand2_1 _16224_ (.Y(_10140_),
    .A(\top_ihp.oisc.regs[14][29] ),
    .B(net536));
 sg13g2_o21ai_1 _16225_ (.B1(_10140_),
    .Y(_00539_),
    .A1(net140),
    .A2(net537));
 sg13g2_nand2_1 _16226_ (.Y(_10141_),
    .A(\top_ihp.oisc.regs[14][2] ),
    .B(_10138_));
 sg13g2_o21ai_1 _16227_ (.B1(_10141_),
    .Y(_00540_),
    .A1(net240),
    .A2(net537));
 sg13g2_nand2_1 _16228_ (.Y(_10142_),
    .A(\top_ihp.oisc.regs[14][30] ),
    .B(_10138_));
 sg13g2_o21ai_1 _16229_ (.B1(_10142_),
    .Y(_00541_),
    .A1(net69),
    .A2(_10133_));
 sg13g2_nand2_1 _16230_ (.Y(_10143_),
    .A(\top_ihp.oisc.regs[14][31] ),
    .B(net536));
 sg13g2_o21ai_1 _16231_ (.B1(_10143_),
    .Y(_00542_),
    .A1(net139),
    .A2(_10133_));
 sg13g2_nand2_1 _16232_ (.Y(_10144_),
    .A(\top_ihp.oisc.regs[14][3] ),
    .B(net536));
 sg13g2_o21ai_1 _16233_ (.B1(_10144_),
    .Y(_00543_),
    .A1(net238),
    .A2(net537));
 sg13g2_nand2_1 _16234_ (.Y(_10145_),
    .A(\top_ihp.oisc.regs[14][4] ),
    .B(net536));
 sg13g2_o21ai_1 _16235_ (.B1(_10145_),
    .Y(_00544_),
    .A1(net237),
    .A2(net539));
 sg13g2_nand2_1 _16236_ (.Y(_10146_),
    .A(\top_ihp.oisc.regs[14][5] ),
    .B(net536));
 sg13g2_o21ai_1 _16237_ (.B1(_10146_),
    .Y(_00545_),
    .A1(net236),
    .A2(net539));
 sg13g2_nand2_1 _16238_ (.Y(_10147_),
    .A(\top_ihp.oisc.regs[14][6] ),
    .B(net536));
 sg13g2_o21ai_1 _16239_ (.B1(_10147_),
    .Y(_00546_),
    .A1(net235),
    .A2(net539));
 sg13g2_nand2_1 _16240_ (.Y(_10148_),
    .A(\top_ihp.oisc.regs[14][7] ),
    .B(net536));
 sg13g2_o21ai_1 _16241_ (.B1(_10148_),
    .Y(_00547_),
    .A1(net68),
    .A2(net539));
 sg13g2_nand2_1 _16242_ (.Y(_10149_),
    .A(\top_ihp.oisc.regs[14][8] ),
    .B(_10111_));
 sg13g2_o21ai_1 _16243_ (.B1(_10149_),
    .Y(_00548_),
    .A1(net67),
    .A2(net539));
 sg13g2_nand2_1 _16244_ (.Y(_10150_),
    .A(\top_ihp.oisc.regs[14][9] ),
    .B(_10111_));
 sg13g2_o21ai_1 _16245_ (.B1(_10150_),
    .Y(_00549_),
    .A1(net66),
    .A2(net539));
 sg13g2_buf_1 _16246_ (.A(_10055_),
    .X(_10151_));
 sg13g2_and2_1 _16247_ (.A(_10011_),
    .B(net665),
    .X(_10152_));
 sg13g2_mux2_1 _16248_ (.A0(\top_ihp.oisc.regs[15][0] ),
    .A1(net210),
    .S(_10152_),
    .X(_00550_));
 sg13g2_nand2_1 _16249_ (.Y(_10153_),
    .A(_10011_),
    .B(net665));
 sg13g2_buf_2 _16250_ (.A(_10153_),
    .X(_10154_));
 sg13g2_buf_1 _16251_ (.A(_10154_),
    .X(_10155_));
 sg13g2_buf_1 _16252_ (.A(_10154_),
    .X(_10156_));
 sg13g2_nand2_1 _16253_ (.Y(_10157_),
    .A(\top_ihp.oisc.regs[15][10] ),
    .B(net400));
 sg13g2_o21ai_1 _16254_ (.B1(_10157_),
    .Y(_00551_),
    .A1(net74),
    .A2(net401));
 sg13g2_nand2_1 _16255_ (.Y(_10158_),
    .A(\top_ihp.oisc.regs[15][11] ),
    .B(net400));
 sg13g2_o21ai_1 _16256_ (.B1(_10158_),
    .Y(_00552_),
    .A1(net148),
    .A2(net401));
 sg13g2_nand2_1 _16257_ (.Y(_10159_),
    .A(\top_ihp.oisc.regs[15][12] ),
    .B(net400));
 sg13g2_o21ai_1 _16258_ (.B1(_10159_),
    .Y(_00553_),
    .A1(net250),
    .A2(net401));
 sg13g2_nand2_1 _16259_ (.Y(_10160_),
    .A(\top_ihp.oisc.regs[15][13] ),
    .B(net400));
 sg13g2_o21ai_1 _16260_ (.B1(_10160_),
    .Y(_00554_),
    .A1(net73),
    .A2(net401));
 sg13g2_nand2_1 _16261_ (.Y(_10161_),
    .A(\top_ihp.oisc.regs[15][14] ),
    .B(net400));
 sg13g2_o21ai_1 _16262_ (.B1(_10161_),
    .Y(_00555_),
    .A1(net249),
    .A2(net401));
 sg13g2_nand2_1 _16263_ (.Y(_10162_),
    .A(\top_ihp.oisc.regs[15][15] ),
    .B(net400));
 sg13g2_o21ai_1 _16264_ (.B1(_10162_),
    .Y(_00556_),
    .A1(net248),
    .A2(net401));
 sg13g2_buf_8 _16265_ (.A(net247),
    .X(_10163_));
 sg13g2_nand2_1 _16266_ (.Y(_10164_),
    .A(\top_ihp.oisc.regs[15][16] ),
    .B(_10156_));
 sg13g2_o21ai_1 _16267_ (.B1(_10164_),
    .Y(_00557_),
    .A1(net130),
    .A2(net401));
 sg13g2_nand2_1 _16268_ (.Y(_10165_),
    .A(\top_ihp.oisc.regs[15][17] ),
    .B(net400));
 sg13g2_o21ai_1 _16269_ (.B1(_10165_),
    .Y(_00558_),
    .A1(net145),
    .A2(_10155_));
 sg13g2_nand2_1 _16270_ (.Y(_10166_),
    .A(\top_ihp.oisc.regs[15][18] ),
    .B(net400));
 sg13g2_o21ai_1 _16271_ (.B1(_10166_),
    .Y(_00559_),
    .A1(net144),
    .A2(net401));
 sg13g2_nand2_1 _16272_ (.Y(_10167_),
    .A(\top_ihp.oisc.regs[15][19] ),
    .B(_10156_));
 sg13g2_o21ai_1 _16273_ (.B1(_10167_),
    .Y(_00560_),
    .A1(net246),
    .A2(_10155_));
 sg13g2_buf_1 _16274_ (.A(_10154_),
    .X(_10168_));
 sg13g2_buf_1 _16275_ (.A(_10154_),
    .X(_10169_));
 sg13g2_nand2_1 _16276_ (.Y(_10170_),
    .A(\top_ihp.oisc.regs[15][1] ),
    .B(net398));
 sg13g2_o21ai_1 _16277_ (.B1(_10170_),
    .Y(_00561_),
    .A1(net409),
    .A2(net399));
 sg13g2_nand2_1 _16278_ (.Y(_10171_),
    .A(\top_ihp.oisc.regs[15][20] ),
    .B(_10169_));
 sg13g2_o21ai_1 _16279_ (.B1(_10171_),
    .Y(_00562_),
    .A1(_09563_),
    .A2(_10168_));
 sg13g2_nand2_1 _16280_ (.Y(_10172_),
    .A(\top_ihp.oisc.regs[15][21] ),
    .B(net398));
 sg13g2_o21ai_1 _16281_ (.B1(_10172_),
    .Y(_00563_),
    .A1(net72),
    .A2(net399));
 sg13g2_nand2_1 _16282_ (.Y(_10173_),
    .A(\top_ihp.oisc.regs[15][22] ),
    .B(net398));
 sg13g2_o21ai_1 _16283_ (.B1(_10173_),
    .Y(_00564_),
    .A1(net143),
    .A2(net399));
 sg13g2_mux2_1 _16284_ (.A0(\top_ihp.oisc.regs[15][23] ),
    .A1(net224),
    .S(_10152_),
    .X(_00565_));
 sg13g2_nand2_1 _16285_ (.Y(_10174_),
    .A(\top_ihp.oisc.regs[15][24] ),
    .B(_10169_));
 sg13g2_o21ai_1 _16286_ (.B1(_10174_),
    .Y(_00566_),
    .A1(net242),
    .A2(_10168_));
 sg13g2_nand2_1 _16287_ (.Y(_10175_),
    .A(\top_ihp.oisc.regs[15][25] ),
    .B(net398));
 sg13g2_o21ai_1 _16288_ (.B1(_10175_),
    .Y(_00567_),
    .A1(net241),
    .A2(net399));
 sg13g2_nand2_1 _16289_ (.Y(_10176_),
    .A(\top_ihp.oisc.regs[15][26] ),
    .B(net398));
 sg13g2_o21ai_1 _16290_ (.B1(_10176_),
    .Y(_00568_),
    .A1(net142),
    .A2(net399));
 sg13g2_nand2_1 _16291_ (.Y(_10177_),
    .A(\top_ihp.oisc.regs[15][27] ),
    .B(net398));
 sg13g2_o21ai_1 _16292_ (.B1(_10177_),
    .Y(_00569_),
    .A1(net71),
    .A2(net399));
 sg13g2_nand2_1 _16293_ (.Y(_10178_),
    .A(\top_ihp.oisc.regs[15][28] ),
    .B(net398));
 sg13g2_o21ai_1 _16294_ (.B1(_10178_),
    .Y(_00570_),
    .A1(net70),
    .A2(net399));
 sg13g2_nand2_1 _16295_ (.Y(_10179_),
    .A(\top_ihp.oisc.regs[15][29] ),
    .B(net398));
 sg13g2_o21ai_1 _16296_ (.B1(_10179_),
    .Y(_00571_),
    .A1(net140),
    .A2(net399));
 sg13g2_buf_1 _16297_ (.A(_10154_),
    .X(_10180_));
 sg13g2_buf_1 _16298_ (.A(_10154_),
    .X(_10181_));
 sg13g2_nand2_1 _16299_ (.Y(_10182_),
    .A(\top_ihp.oisc.regs[15][2] ),
    .B(net396));
 sg13g2_o21ai_1 _16300_ (.B1(_10182_),
    .Y(_00572_),
    .A1(net240),
    .A2(net397));
 sg13g2_nand2_1 _16301_ (.Y(_10183_),
    .A(\top_ihp.oisc.regs[15][30] ),
    .B(_10181_));
 sg13g2_o21ai_1 _16302_ (.B1(_10183_),
    .Y(_00573_),
    .A1(net69),
    .A2(_10180_));
 sg13g2_nand2_1 _16303_ (.Y(_10184_),
    .A(\top_ihp.oisc.regs[15][31] ),
    .B(net396));
 sg13g2_o21ai_1 _16304_ (.B1(_10184_),
    .Y(_00574_),
    .A1(net139),
    .A2(_10180_));
 sg13g2_nand2_1 _16305_ (.Y(_10185_),
    .A(\top_ihp.oisc.regs[15][3] ),
    .B(_10181_));
 sg13g2_o21ai_1 _16306_ (.B1(_10185_),
    .Y(_00575_),
    .A1(net238),
    .A2(net397));
 sg13g2_nand2_1 _16307_ (.Y(_10186_),
    .A(\top_ihp.oisc.regs[15][4] ),
    .B(net396));
 sg13g2_o21ai_1 _16308_ (.B1(_10186_),
    .Y(_00576_),
    .A1(net237),
    .A2(net397));
 sg13g2_nand2_1 _16309_ (.Y(_10187_),
    .A(\top_ihp.oisc.regs[15][5] ),
    .B(net396));
 sg13g2_o21ai_1 _16310_ (.B1(_10187_),
    .Y(_00577_),
    .A1(net236),
    .A2(net397));
 sg13g2_nand2_1 _16311_ (.Y(_10188_),
    .A(\top_ihp.oisc.regs[15][6] ),
    .B(net396));
 sg13g2_o21ai_1 _16312_ (.B1(_10188_),
    .Y(_00578_),
    .A1(net235),
    .A2(net397));
 sg13g2_buf_2 _16313_ (.A(net408),
    .X(_10189_));
 sg13g2_nand2_1 _16314_ (.Y(_10190_),
    .A(\top_ihp.oisc.regs[15][7] ),
    .B(net396));
 sg13g2_o21ai_1 _16315_ (.B1(_10190_),
    .Y(_00579_),
    .A1(net209),
    .A2(net397));
 sg13g2_nand2_1 _16316_ (.Y(_10191_),
    .A(\top_ihp.oisc.regs[15][8] ),
    .B(net396));
 sg13g2_o21ai_1 _16317_ (.B1(_10191_),
    .Y(_00580_),
    .A1(net67),
    .A2(net397));
 sg13g2_nand2_1 _16318_ (.Y(_10192_),
    .A(\top_ihp.oisc.regs[15][9] ),
    .B(net396));
 sg13g2_o21ai_1 _16319_ (.B1(_10192_),
    .Y(_00581_),
    .A1(net66),
    .A2(net397));
 sg13g2_buf_1 _16320_ (.A(\top_ihp.oisc.regs[16][0] ),
    .X(_00582_));
 sg13g2_buf_1 _16321_ (.A(\top_ihp.oisc.regs[16][10] ),
    .X(_00583_));
 sg13g2_buf_1 _16322_ (.A(\top_ihp.oisc.regs[16][11] ),
    .X(_00584_));
 sg13g2_buf_1 _16323_ (.A(\top_ihp.oisc.regs[16][12] ),
    .X(_00585_));
 sg13g2_buf_1 _16324_ (.A(\top_ihp.oisc.regs[16][13] ),
    .X(_00586_));
 sg13g2_buf_1 _16325_ (.A(\top_ihp.oisc.regs[16][14] ),
    .X(_00587_));
 sg13g2_buf_1 _16326_ (.A(\top_ihp.oisc.regs[16][15] ),
    .X(_00588_));
 sg13g2_buf_1 _16327_ (.A(\top_ihp.oisc.regs[16][16] ),
    .X(_00589_));
 sg13g2_buf_1 _16328_ (.A(\top_ihp.oisc.regs[16][17] ),
    .X(_00590_));
 sg13g2_buf_1 _16329_ (.A(\top_ihp.oisc.regs[16][18] ),
    .X(_00591_));
 sg13g2_buf_1 _16330_ (.A(\top_ihp.oisc.regs[16][19] ),
    .X(_00592_));
 sg13g2_buf_1 _16331_ (.A(\top_ihp.oisc.regs[16][1] ),
    .X(_00593_));
 sg13g2_buf_1 _16332_ (.A(\top_ihp.oisc.regs[16][20] ),
    .X(_00594_));
 sg13g2_buf_1 _16333_ (.A(\top_ihp.oisc.regs[16][21] ),
    .X(_00595_));
 sg13g2_buf_1 _16334_ (.A(\top_ihp.oisc.regs[16][22] ),
    .X(_00596_));
 sg13g2_buf_1 _16335_ (.A(\top_ihp.oisc.regs[16][23] ),
    .X(_00597_));
 sg13g2_buf_1 _16336_ (.A(\top_ihp.oisc.regs[16][24] ),
    .X(_00598_));
 sg13g2_buf_1 _16337_ (.A(\top_ihp.oisc.regs[16][25] ),
    .X(_00599_));
 sg13g2_buf_1 _16338_ (.A(\top_ihp.oisc.regs[16][26] ),
    .X(_00600_));
 sg13g2_buf_1 _16339_ (.A(\top_ihp.oisc.regs[16][27] ),
    .X(_00601_));
 sg13g2_buf_1 _16340_ (.A(\top_ihp.oisc.regs[16][28] ),
    .X(_00602_));
 sg13g2_buf_1 _16341_ (.A(\top_ihp.oisc.regs[16][29] ),
    .X(_00603_));
 sg13g2_buf_1 _16342_ (.A(\top_ihp.oisc.regs[16][2] ),
    .X(_00604_));
 sg13g2_buf_1 _16343_ (.A(\top_ihp.oisc.regs[16][30] ),
    .X(_00605_));
 sg13g2_buf_1 _16344_ (.A(\top_ihp.oisc.regs[16][31] ),
    .X(_00606_));
 sg13g2_buf_1 _16345_ (.A(\top_ihp.oisc.regs[16][3] ),
    .X(_00607_));
 sg13g2_buf_1 _16346_ (.A(\top_ihp.oisc.regs[16][4] ),
    .X(_00608_));
 sg13g2_buf_1 _16347_ (.A(\top_ihp.oisc.regs[16][5] ),
    .X(_00609_));
 sg13g2_buf_1 _16348_ (.A(\top_ihp.oisc.regs[16][6] ),
    .X(_00610_));
 sg13g2_buf_1 _16349_ (.A(\top_ihp.oisc.regs[16][7] ),
    .X(_00611_));
 sg13g2_buf_1 _16350_ (.A(\top_ihp.oisc.regs[16][8] ),
    .X(_00612_));
 sg13g2_buf_1 _16351_ (.A(\top_ihp.oisc.regs[16][9] ),
    .X(_00613_));
 sg13g2_buf_1 _16352_ (.A(\top_ihp.oisc.regs[17][0] ),
    .X(_00614_));
 sg13g2_buf_1 _16353_ (.A(\top_ihp.oisc.regs[17][10] ),
    .X(_00615_));
 sg13g2_buf_1 _16354_ (.A(\top_ihp.oisc.regs[17][11] ),
    .X(_00616_));
 sg13g2_buf_1 _16355_ (.A(\top_ihp.oisc.regs[17][12] ),
    .X(_00617_));
 sg13g2_buf_1 _16356_ (.A(\top_ihp.oisc.regs[17][13] ),
    .X(_00618_));
 sg13g2_buf_1 _16357_ (.A(\top_ihp.oisc.regs[17][14] ),
    .X(_00619_));
 sg13g2_buf_1 _16358_ (.A(\top_ihp.oisc.regs[17][15] ),
    .X(_00620_));
 sg13g2_buf_1 _16359_ (.A(\top_ihp.oisc.regs[17][16] ),
    .X(_00621_));
 sg13g2_buf_1 _16360_ (.A(\top_ihp.oisc.regs[17][17] ),
    .X(_00622_));
 sg13g2_buf_1 _16361_ (.A(\top_ihp.oisc.regs[17][18] ),
    .X(_00623_));
 sg13g2_buf_1 _16362_ (.A(\top_ihp.oisc.regs[17][19] ),
    .X(_00624_));
 sg13g2_buf_1 _16363_ (.A(\top_ihp.oisc.regs[17][1] ),
    .X(_00625_));
 sg13g2_buf_1 _16364_ (.A(\top_ihp.oisc.regs[17][20] ),
    .X(_00626_));
 sg13g2_buf_1 _16365_ (.A(\top_ihp.oisc.regs[17][21] ),
    .X(_00627_));
 sg13g2_buf_1 _16366_ (.A(\top_ihp.oisc.regs[17][22] ),
    .X(_00628_));
 sg13g2_buf_1 _16367_ (.A(\top_ihp.oisc.regs[17][23] ),
    .X(_00629_));
 sg13g2_buf_1 _16368_ (.A(\top_ihp.oisc.regs[17][24] ),
    .X(_00630_));
 sg13g2_buf_1 _16369_ (.A(\top_ihp.oisc.regs[17][25] ),
    .X(_00631_));
 sg13g2_buf_1 _16370_ (.A(\top_ihp.oisc.regs[17][26] ),
    .X(_00632_));
 sg13g2_buf_1 _16371_ (.A(\top_ihp.oisc.regs[17][27] ),
    .X(_00633_));
 sg13g2_buf_1 _16372_ (.A(\top_ihp.oisc.regs[17][28] ),
    .X(_00634_));
 sg13g2_buf_1 _16373_ (.A(\top_ihp.oisc.regs[17][29] ),
    .X(_00635_));
 sg13g2_buf_1 _16374_ (.A(\top_ihp.oisc.regs[17][2] ),
    .X(_00636_));
 sg13g2_buf_1 _16375_ (.A(\top_ihp.oisc.regs[17][30] ),
    .X(_00637_));
 sg13g2_buf_1 _16376_ (.A(\top_ihp.oisc.regs[17][31] ),
    .X(_00638_));
 sg13g2_buf_1 _16377_ (.A(\top_ihp.oisc.regs[17][3] ),
    .X(_00639_));
 sg13g2_buf_1 _16378_ (.A(\top_ihp.oisc.regs[17][4] ),
    .X(_00640_));
 sg13g2_buf_1 _16379_ (.A(\top_ihp.oisc.regs[17][5] ),
    .X(_00641_));
 sg13g2_buf_1 _16380_ (.A(\top_ihp.oisc.regs[17][6] ),
    .X(_00642_));
 sg13g2_buf_1 _16381_ (.A(\top_ihp.oisc.regs[17][7] ),
    .X(_00643_));
 sg13g2_buf_1 _16382_ (.A(\top_ihp.oisc.regs[17][8] ),
    .X(_00644_));
 sg13g2_buf_1 _16383_ (.A(\top_ihp.oisc.regs[17][9] ),
    .X(_00645_));
 sg13g2_buf_1 _16384_ (.A(\top_ihp.oisc.regs[18][0] ),
    .X(_00646_));
 sg13g2_buf_1 _16385_ (.A(\top_ihp.oisc.regs[18][10] ),
    .X(_00647_));
 sg13g2_buf_1 _16386_ (.A(\top_ihp.oisc.regs[18][11] ),
    .X(_00648_));
 sg13g2_buf_1 _16387_ (.A(\top_ihp.oisc.regs[18][12] ),
    .X(_00649_));
 sg13g2_buf_1 _16388_ (.A(\top_ihp.oisc.regs[18][13] ),
    .X(_00650_));
 sg13g2_buf_1 _16389_ (.A(\top_ihp.oisc.regs[18][14] ),
    .X(_00651_));
 sg13g2_buf_1 _16390_ (.A(\top_ihp.oisc.regs[18][15] ),
    .X(_00652_));
 sg13g2_buf_1 _16391_ (.A(\top_ihp.oisc.regs[18][16] ),
    .X(_00653_));
 sg13g2_buf_1 _16392_ (.A(\top_ihp.oisc.regs[18][17] ),
    .X(_00654_));
 sg13g2_buf_1 _16393_ (.A(\top_ihp.oisc.regs[18][18] ),
    .X(_00655_));
 sg13g2_buf_1 _16394_ (.A(\top_ihp.oisc.regs[18][19] ),
    .X(_00656_));
 sg13g2_buf_1 _16395_ (.A(\top_ihp.oisc.regs[18][1] ),
    .X(_00657_));
 sg13g2_buf_1 _16396_ (.A(\top_ihp.oisc.regs[18][20] ),
    .X(_00658_));
 sg13g2_buf_1 _16397_ (.A(\top_ihp.oisc.regs[18][21] ),
    .X(_00659_));
 sg13g2_buf_1 _16398_ (.A(\top_ihp.oisc.regs[18][22] ),
    .X(_00660_));
 sg13g2_buf_1 _16399_ (.A(\top_ihp.oisc.regs[18][23] ),
    .X(_00661_));
 sg13g2_buf_1 _16400_ (.A(\top_ihp.oisc.regs[18][24] ),
    .X(_00662_));
 sg13g2_buf_1 _16401_ (.A(\top_ihp.oisc.regs[18][25] ),
    .X(_00663_));
 sg13g2_buf_1 _16402_ (.A(\top_ihp.oisc.regs[18][26] ),
    .X(_00664_));
 sg13g2_buf_1 _16403_ (.A(\top_ihp.oisc.regs[18][27] ),
    .X(_00665_));
 sg13g2_buf_1 _16404_ (.A(\top_ihp.oisc.regs[18][28] ),
    .X(_00666_));
 sg13g2_buf_1 _16405_ (.A(\top_ihp.oisc.regs[18][29] ),
    .X(_00667_));
 sg13g2_buf_1 _16406_ (.A(\top_ihp.oisc.regs[18][2] ),
    .X(_00668_));
 sg13g2_buf_1 _16407_ (.A(\top_ihp.oisc.regs[18][30] ),
    .X(_00669_));
 sg13g2_buf_1 _16408_ (.A(\top_ihp.oisc.regs[18][31] ),
    .X(_00670_));
 sg13g2_buf_1 _16409_ (.A(\top_ihp.oisc.regs[18][3] ),
    .X(_00671_));
 sg13g2_buf_1 _16410_ (.A(\top_ihp.oisc.regs[18][4] ),
    .X(_00672_));
 sg13g2_buf_1 _16411_ (.A(\top_ihp.oisc.regs[18][5] ),
    .X(_00673_));
 sg13g2_buf_1 _16412_ (.A(\top_ihp.oisc.regs[18][6] ),
    .X(_00674_));
 sg13g2_buf_1 _16413_ (.A(\top_ihp.oisc.regs[18][7] ),
    .X(_00675_));
 sg13g2_buf_1 _16414_ (.A(\top_ihp.oisc.regs[18][8] ),
    .X(_00676_));
 sg13g2_buf_1 _16415_ (.A(\top_ihp.oisc.regs[18][9] ),
    .X(_00677_));
 sg13g2_buf_1 _16416_ (.A(\top_ihp.oisc.regs[19][0] ),
    .X(_00678_));
 sg13g2_buf_1 _16417_ (.A(\top_ihp.oisc.regs[19][10] ),
    .X(_00679_));
 sg13g2_buf_1 _16418_ (.A(\top_ihp.oisc.regs[19][11] ),
    .X(_00680_));
 sg13g2_buf_1 _16419_ (.A(\top_ihp.oisc.regs[19][12] ),
    .X(_00681_));
 sg13g2_buf_1 _16420_ (.A(\top_ihp.oisc.regs[19][13] ),
    .X(_00682_));
 sg13g2_buf_1 _16421_ (.A(\top_ihp.oisc.regs[19][14] ),
    .X(_00683_));
 sg13g2_buf_1 _16422_ (.A(\top_ihp.oisc.regs[19][15] ),
    .X(_00684_));
 sg13g2_buf_1 _16423_ (.A(\top_ihp.oisc.regs[19][16] ),
    .X(_00685_));
 sg13g2_buf_1 _16424_ (.A(\top_ihp.oisc.regs[19][17] ),
    .X(_00686_));
 sg13g2_buf_1 _16425_ (.A(\top_ihp.oisc.regs[19][18] ),
    .X(_00687_));
 sg13g2_buf_1 _16426_ (.A(\top_ihp.oisc.regs[19][19] ),
    .X(_00688_));
 sg13g2_buf_1 _16427_ (.A(\top_ihp.oisc.regs[19][1] ),
    .X(_00689_));
 sg13g2_buf_1 _16428_ (.A(\top_ihp.oisc.regs[19][20] ),
    .X(_00690_));
 sg13g2_buf_1 _16429_ (.A(\top_ihp.oisc.regs[19][21] ),
    .X(_00691_));
 sg13g2_buf_1 _16430_ (.A(\top_ihp.oisc.regs[19][22] ),
    .X(_00692_));
 sg13g2_buf_1 _16431_ (.A(\top_ihp.oisc.regs[19][23] ),
    .X(_00693_));
 sg13g2_buf_1 _16432_ (.A(\top_ihp.oisc.regs[19][24] ),
    .X(_00694_));
 sg13g2_buf_1 _16433_ (.A(\top_ihp.oisc.regs[19][25] ),
    .X(_00695_));
 sg13g2_buf_1 _16434_ (.A(\top_ihp.oisc.regs[19][26] ),
    .X(_00696_));
 sg13g2_buf_1 _16435_ (.A(\top_ihp.oisc.regs[19][27] ),
    .X(_00697_));
 sg13g2_buf_1 _16436_ (.A(\top_ihp.oisc.regs[19][28] ),
    .X(_00698_));
 sg13g2_buf_1 _16437_ (.A(\top_ihp.oisc.regs[19][29] ),
    .X(_00699_));
 sg13g2_buf_1 _16438_ (.A(\top_ihp.oisc.regs[19][2] ),
    .X(_00700_));
 sg13g2_buf_1 _16439_ (.A(\top_ihp.oisc.regs[19][30] ),
    .X(_00701_));
 sg13g2_buf_1 _16440_ (.A(\top_ihp.oisc.regs[19][31] ),
    .X(_00702_));
 sg13g2_buf_1 _16441_ (.A(\top_ihp.oisc.regs[19][3] ),
    .X(_00703_));
 sg13g2_buf_1 _16442_ (.A(\top_ihp.oisc.regs[19][4] ),
    .X(_00704_));
 sg13g2_buf_1 _16443_ (.A(\top_ihp.oisc.regs[19][5] ),
    .X(_00705_));
 sg13g2_buf_1 _16444_ (.A(\top_ihp.oisc.regs[19][6] ),
    .X(_00706_));
 sg13g2_buf_1 _16445_ (.A(\top_ihp.oisc.regs[19][7] ),
    .X(_00707_));
 sg13g2_buf_1 _16446_ (.A(\top_ihp.oisc.regs[19][8] ),
    .X(_00708_));
 sg13g2_buf_1 _16447_ (.A(\top_ihp.oisc.regs[19][9] ),
    .X(_00709_));
 sg13g2_and2_1 _16448_ (.A(_09106_),
    .B(net710),
    .X(_10193_));
 sg13g2_buf_2 _16449_ (.A(_10193_),
    .X(_10194_));
 sg13g2_mux2_1 _16450_ (.A0(\top_ihp.oisc.regs[1][0] ),
    .A1(net210),
    .S(_10194_),
    .X(_00710_));
 sg13g2_nand2_1 _16451_ (.Y(_10195_),
    .A(_09106_),
    .B(net710));
 sg13g2_buf_1 _16452_ (.A(_10195_),
    .X(_10196_));
 sg13g2_buf_1 _16453_ (.A(net639),
    .X(_10197_));
 sg13g2_buf_1 _16454_ (.A(_10195_),
    .X(_10198_));
 sg13g2_nand2_1 _16455_ (.Y(_10199_),
    .A(\top_ihp.oisc.regs[1][10] ),
    .B(net638));
 sg13g2_o21ai_1 _16456_ (.B1(_10199_),
    .Y(_00711_),
    .A1(net74),
    .A2(net535));
 sg13g2_nand2_1 _16457_ (.Y(_10200_),
    .A(\top_ihp.oisc.regs[1][11] ),
    .B(net638));
 sg13g2_o21ai_1 _16458_ (.B1(_10200_),
    .Y(_00712_),
    .A1(net148),
    .A2(net535));
 sg13g2_buf_1 _16459_ (.A(net639),
    .X(_10201_));
 sg13g2_nand2_1 _16460_ (.Y(_10202_),
    .A(\top_ihp.oisc.regs[1][12] ),
    .B(net534));
 sg13g2_o21ai_1 _16461_ (.B1(_10202_),
    .Y(_00713_),
    .A1(net250),
    .A2(net535));
 sg13g2_buf_8 _16462_ (.A(net147),
    .X(_10203_));
 sg13g2_nand2_1 _16463_ (.Y(_10204_),
    .A(\top_ihp.oisc.regs[1][13] ),
    .B(net534));
 sg13g2_o21ai_1 _16464_ (.B1(_10204_),
    .Y(_00714_),
    .A1(net58),
    .A2(net535));
 sg13g2_nand2_1 _16465_ (.Y(_10205_),
    .A(\top_ihp.oisc.regs[1][14] ),
    .B(net534));
 sg13g2_o21ai_1 _16466_ (.B1(_10205_),
    .Y(_00715_),
    .A1(net249),
    .A2(net535));
 sg13g2_nand2_1 _16467_ (.Y(_10206_),
    .A(\top_ihp.oisc.regs[1][15] ),
    .B(net534));
 sg13g2_o21ai_1 _16468_ (.B1(_10206_),
    .Y(_00716_),
    .A1(net248),
    .A2(net535));
 sg13g2_nand2_1 _16469_ (.Y(_10207_),
    .A(\top_ihp.oisc.regs[1][16] ),
    .B(_10201_));
 sg13g2_o21ai_1 _16470_ (.B1(_10207_),
    .Y(_00717_),
    .A1(net130),
    .A2(net535));
 sg13g2_nand2_1 _16471_ (.Y(_10208_),
    .A(\top_ihp.oisc.regs[1][17] ),
    .B(net534));
 sg13g2_o21ai_1 _16472_ (.B1(_10208_),
    .Y(_00718_),
    .A1(net145),
    .A2(net535));
 sg13g2_nand2_1 _16473_ (.Y(_10209_),
    .A(\top_ihp.oisc.regs[1][18] ),
    .B(net534));
 sg13g2_o21ai_1 _16474_ (.B1(_10209_),
    .Y(_00719_),
    .A1(net144),
    .A2(_10197_));
 sg13g2_nand2_1 _16475_ (.Y(_10210_),
    .A(\top_ihp.oisc.regs[1][19] ),
    .B(_10201_));
 sg13g2_o21ai_1 _16476_ (.B1(_10210_),
    .Y(_00720_),
    .A1(net246),
    .A2(_10197_));
 sg13g2_buf_1 _16477_ (.A(net639),
    .X(_10211_));
 sg13g2_nand2_1 _16478_ (.Y(_10212_),
    .A(\top_ihp.oisc.regs[1][1] ),
    .B(net534));
 sg13g2_o21ai_1 _16479_ (.B1(_10212_),
    .Y(_00721_),
    .A1(net409),
    .A2(net533));
 sg13g2_mux2_1 _16480_ (.A0(\top_ihp.oisc.regs[1][20] ),
    .A1(net137),
    .S(_10194_),
    .X(_00722_));
 sg13g2_nand2_1 _16481_ (.Y(_10213_),
    .A(\top_ihp.oisc.regs[1][21] ),
    .B(net534));
 sg13g2_o21ai_1 _16482_ (.B1(_10213_),
    .Y(_00723_),
    .A1(net72),
    .A2(net533));
 sg13g2_buf_1 _16483_ (.A(net244),
    .X(_10214_));
 sg13g2_buf_1 _16484_ (.A(_10196_),
    .X(_10215_));
 sg13g2_nand2_1 _16485_ (.Y(_10216_),
    .A(\top_ihp.oisc.regs[1][22] ),
    .B(net532));
 sg13g2_o21ai_1 _16486_ (.B1(_10216_),
    .Y(_00724_),
    .A1(net129),
    .A2(net533));
 sg13g2_mux2_1 _16487_ (.A0(\top_ihp.oisc.regs[1][23] ),
    .A1(net224),
    .S(_10194_),
    .X(_00725_));
 sg13g2_nand2_1 _16488_ (.Y(_10217_),
    .A(\top_ihp.oisc.regs[1][24] ),
    .B(net532));
 sg13g2_o21ai_1 _16489_ (.B1(_10217_),
    .Y(_00726_),
    .A1(net242),
    .A2(net533));
 sg13g2_nand2_1 _16490_ (.Y(_10218_),
    .A(\top_ihp.oisc.regs[1][25] ),
    .B(net532));
 sg13g2_o21ai_1 _16491_ (.B1(_10218_),
    .Y(_00727_),
    .A1(net241),
    .A2(net533));
 sg13g2_nand2_1 _16492_ (.Y(_10219_),
    .A(\top_ihp.oisc.regs[1][26] ),
    .B(_10215_));
 sg13g2_o21ai_1 _16493_ (.B1(_10219_),
    .Y(_00728_),
    .A1(net142),
    .A2(_10211_));
 sg13g2_nand2_1 _16494_ (.Y(_10220_),
    .A(\top_ihp.oisc.regs[1][27] ),
    .B(net532));
 sg13g2_o21ai_1 _16495_ (.B1(_10220_),
    .Y(_00729_),
    .A1(net71),
    .A2(net533));
 sg13g2_nand2_1 _16496_ (.Y(_10221_),
    .A(\top_ihp.oisc.regs[1][28] ),
    .B(net532));
 sg13g2_o21ai_1 _16497_ (.B1(_10221_),
    .Y(_00730_),
    .A1(net70),
    .A2(_10211_));
 sg13g2_nand2_1 _16498_ (.Y(_10222_),
    .A(\top_ihp.oisc.regs[1][29] ),
    .B(net532));
 sg13g2_o21ai_1 _16499_ (.B1(_10222_),
    .Y(_00731_),
    .A1(net140),
    .A2(net533));
 sg13g2_nand2_1 _16500_ (.Y(_10223_),
    .A(\top_ihp.oisc.regs[1][2] ),
    .B(net532));
 sg13g2_o21ai_1 _16501_ (.B1(_10223_),
    .Y(_00732_),
    .A1(net240),
    .A2(net533));
 sg13g2_mux2_1 _16502_ (.A0(_00209_),
    .A1(net62),
    .S(_10194_),
    .X(_00733_));
 sg13g2_nand2_1 _16503_ (.Y(_10224_),
    .A(\top_ihp.oisc.regs[1][31] ),
    .B(_10215_));
 sg13g2_o21ai_1 _16504_ (.B1(_10224_),
    .Y(_00734_),
    .A1(net139),
    .A2(net638));
 sg13g2_nand2_1 _16505_ (.Y(_10225_),
    .A(\top_ihp.oisc.regs[1][3] ),
    .B(net532));
 sg13g2_o21ai_1 _16506_ (.B1(_10225_),
    .Y(_00735_),
    .A1(net238),
    .A2(_10198_));
 sg13g2_nand2_1 _16507_ (.Y(_10226_),
    .A(\top_ihp.oisc.regs[1][4] ),
    .B(_10196_));
 sg13g2_o21ai_1 _16508_ (.B1(_10226_),
    .Y(_00736_),
    .A1(net237),
    .A2(_10198_));
 sg13g2_nand2_1 _16509_ (.Y(_10227_),
    .A(\top_ihp.oisc.regs[1][5] ),
    .B(net639));
 sg13g2_o21ai_1 _16510_ (.B1(_10227_),
    .Y(_00737_),
    .A1(net236),
    .A2(net638));
 sg13g2_nand2_1 _16511_ (.Y(_10228_),
    .A(\top_ihp.oisc.regs[1][6] ),
    .B(net639));
 sg13g2_o21ai_1 _16512_ (.B1(_10228_),
    .Y(_00738_),
    .A1(net235),
    .A2(net638));
 sg13g2_nand2_1 _16513_ (.Y(_10229_),
    .A(\top_ihp.oisc.regs[1][7] ),
    .B(net639));
 sg13g2_o21ai_1 _16514_ (.B1(_10229_),
    .Y(_00739_),
    .A1(net209),
    .A2(net638));
 sg13g2_nand2_1 _16515_ (.Y(_10230_),
    .A(\top_ihp.oisc.regs[1][8] ),
    .B(net639));
 sg13g2_o21ai_1 _16516_ (.B1(_10230_),
    .Y(_00740_),
    .A1(net67),
    .A2(net638));
 sg13g2_nand2_1 _16517_ (.Y(_10231_),
    .A(\top_ihp.oisc.regs[1][9] ),
    .B(net639));
 sg13g2_o21ai_1 _16518_ (.B1(_10231_),
    .Y(_00741_),
    .A1(net66),
    .A2(net638));
 sg13g2_buf_1 _16519_ (.A(\top_ihp.oisc.regs[20][0] ),
    .X(_00742_));
 sg13g2_buf_1 _16520_ (.A(\top_ihp.oisc.regs[20][10] ),
    .X(_00743_));
 sg13g2_buf_1 _16521_ (.A(\top_ihp.oisc.regs[20][11] ),
    .X(_00744_));
 sg13g2_buf_1 _16522_ (.A(\top_ihp.oisc.regs[20][12] ),
    .X(_00745_));
 sg13g2_buf_1 _16523_ (.A(\top_ihp.oisc.regs[20][13] ),
    .X(_00746_));
 sg13g2_buf_1 _16524_ (.A(\top_ihp.oisc.regs[20][14] ),
    .X(_00747_));
 sg13g2_buf_1 _16525_ (.A(\top_ihp.oisc.regs[20][15] ),
    .X(_00748_));
 sg13g2_buf_1 _16526_ (.A(\top_ihp.oisc.regs[20][16] ),
    .X(_00749_));
 sg13g2_buf_1 _16527_ (.A(\top_ihp.oisc.regs[20][17] ),
    .X(_00750_));
 sg13g2_buf_1 _16528_ (.A(\top_ihp.oisc.regs[20][18] ),
    .X(_00751_));
 sg13g2_buf_1 _16529_ (.A(\top_ihp.oisc.regs[20][19] ),
    .X(_00752_));
 sg13g2_buf_1 _16530_ (.A(\top_ihp.oisc.regs[20][1] ),
    .X(_00753_));
 sg13g2_buf_1 _16531_ (.A(\top_ihp.oisc.regs[20][20] ),
    .X(_00754_));
 sg13g2_buf_1 _16532_ (.A(\top_ihp.oisc.regs[20][21] ),
    .X(_00755_));
 sg13g2_buf_1 _16533_ (.A(\top_ihp.oisc.regs[20][22] ),
    .X(_00756_));
 sg13g2_buf_1 _16534_ (.A(\top_ihp.oisc.regs[20][23] ),
    .X(_00757_));
 sg13g2_buf_1 _16535_ (.A(\top_ihp.oisc.regs[20][24] ),
    .X(_00758_));
 sg13g2_buf_1 _16536_ (.A(\top_ihp.oisc.regs[20][25] ),
    .X(_00759_));
 sg13g2_buf_1 _16537_ (.A(\top_ihp.oisc.regs[20][26] ),
    .X(_00760_));
 sg13g2_buf_1 _16538_ (.A(\top_ihp.oisc.regs[20][27] ),
    .X(_00761_));
 sg13g2_buf_1 _16539_ (.A(\top_ihp.oisc.regs[20][28] ),
    .X(_00762_));
 sg13g2_buf_1 _16540_ (.A(\top_ihp.oisc.regs[20][29] ),
    .X(_00763_));
 sg13g2_buf_1 _16541_ (.A(\top_ihp.oisc.regs[20][2] ),
    .X(_00764_));
 sg13g2_buf_1 _16542_ (.A(\top_ihp.oisc.regs[20][30] ),
    .X(_00765_));
 sg13g2_buf_1 _16543_ (.A(\top_ihp.oisc.regs[20][31] ),
    .X(_00766_));
 sg13g2_buf_1 _16544_ (.A(\top_ihp.oisc.regs[20][3] ),
    .X(_00767_));
 sg13g2_buf_1 _16545_ (.A(\top_ihp.oisc.regs[20][4] ),
    .X(_00768_));
 sg13g2_buf_1 _16546_ (.A(\top_ihp.oisc.regs[20][5] ),
    .X(_00769_));
 sg13g2_buf_1 _16547_ (.A(\top_ihp.oisc.regs[20][6] ),
    .X(_00770_));
 sg13g2_buf_1 _16548_ (.A(\top_ihp.oisc.regs[20][7] ),
    .X(_00771_));
 sg13g2_buf_1 _16549_ (.A(\top_ihp.oisc.regs[20][8] ),
    .X(_00772_));
 sg13g2_buf_1 _16550_ (.A(\top_ihp.oisc.regs[20][9] ),
    .X(_00773_));
 sg13g2_buf_1 _16551_ (.A(\top_ihp.oisc.regs[21][0] ),
    .X(_00774_));
 sg13g2_buf_1 _16552_ (.A(\top_ihp.oisc.regs[21][10] ),
    .X(_00775_));
 sg13g2_buf_1 _16553_ (.A(\top_ihp.oisc.regs[21][11] ),
    .X(_00776_));
 sg13g2_buf_1 _16554_ (.A(\top_ihp.oisc.regs[21][12] ),
    .X(_00777_));
 sg13g2_buf_1 _16555_ (.A(\top_ihp.oisc.regs[21][13] ),
    .X(_00778_));
 sg13g2_buf_1 _16556_ (.A(\top_ihp.oisc.regs[21][14] ),
    .X(_00779_));
 sg13g2_buf_1 _16557_ (.A(\top_ihp.oisc.regs[21][15] ),
    .X(_00780_));
 sg13g2_buf_1 _16558_ (.A(\top_ihp.oisc.regs[21][16] ),
    .X(_00781_));
 sg13g2_buf_1 _16559_ (.A(\top_ihp.oisc.regs[21][17] ),
    .X(_00782_));
 sg13g2_buf_1 _16560_ (.A(\top_ihp.oisc.regs[21][18] ),
    .X(_00783_));
 sg13g2_buf_1 _16561_ (.A(\top_ihp.oisc.regs[21][19] ),
    .X(_00784_));
 sg13g2_buf_1 _16562_ (.A(\top_ihp.oisc.regs[21][1] ),
    .X(_00785_));
 sg13g2_buf_1 _16563_ (.A(\top_ihp.oisc.regs[21][20] ),
    .X(_00786_));
 sg13g2_buf_1 _16564_ (.A(\top_ihp.oisc.regs[21][21] ),
    .X(_00787_));
 sg13g2_buf_1 _16565_ (.A(\top_ihp.oisc.regs[21][22] ),
    .X(_00788_));
 sg13g2_buf_1 _16566_ (.A(\top_ihp.oisc.regs[21][23] ),
    .X(_00789_));
 sg13g2_buf_1 _16567_ (.A(\top_ihp.oisc.regs[21][24] ),
    .X(_00790_));
 sg13g2_buf_1 _16568_ (.A(\top_ihp.oisc.regs[21][25] ),
    .X(_00791_));
 sg13g2_buf_1 _16569_ (.A(\top_ihp.oisc.regs[21][26] ),
    .X(_00792_));
 sg13g2_buf_1 _16570_ (.A(\top_ihp.oisc.regs[21][27] ),
    .X(_00793_));
 sg13g2_buf_1 _16571_ (.A(\top_ihp.oisc.regs[21][28] ),
    .X(_00794_));
 sg13g2_buf_1 _16572_ (.A(\top_ihp.oisc.regs[21][29] ),
    .X(_00795_));
 sg13g2_buf_1 _16573_ (.A(\top_ihp.oisc.regs[21][2] ),
    .X(_00796_));
 sg13g2_buf_1 _16574_ (.A(\top_ihp.oisc.regs[21][30] ),
    .X(_00797_));
 sg13g2_buf_1 _16575_ (.A(\top_ihp.oisc.regs[21][31] ),
    .X(_00798_));
 sg13g2_buf_1 _16576_ (.A(\top_ihp.oisc.regs[21][3] ),
    .X(_00799_));
 sg13g2_buf_1 _16577_ (.A(\top_ihp.oisc.regs[21][4] ),
    .X(_00800_));
 sg13g2_buf_1 _16578_ (.A(\top_ihp.oisc.regs[21][5] ),
    .X(_00801_));
 sg13g2_buf_1 _16579_ (.A(\top_ihp.oisc.regs[21][6] ),
    .X(_00802_));
 sg13g2_buf_1 _16580_ (.A(\top_ihp.oisc.regs[21][7] ),
    .X(_00803_));
 sg13g2_buf_1 _16581_ (.A(\top_ihp.oisc.regs[21][8] ),
    .X(_00804_));
 sg13g2_buf_1 _16582_ (.A(\top_ihp.oisc.regs[21][9] ),
    .X(_00805_));
 sg13g2_buf_1 _16583_ (.A(\top_ihp.oisc.regs[22][0] ),
    .X(_00806_));
 sg13g2_buf_1 _16584_ (.A(\top_ihp.oisc.regs[22][10] ),
    .X(_00807_));
 sg13g2_buf_1 _16585_ (.A(\top_ihp.oisc.regs[22][11] ),
    .X(_00808_));
 sg13g2_buf_1 _16586_ (.A(\top_ihp.oisc.regs[22][12] ),
    .X(_00809_));
 sg13g2_buf_1 _16587_ (.A(\top_ihp.oisc.regs[22][13] ),
    .X(_00810_));
 sg13g2_buf_1 _16588_ (.A(\top_ihp.oisc.regs[22][14] ),
    .X(_00811_));
 sg13g2_buf_1 _16589_ (.A(\top_ihp.oisc.regs[22][15] ),
    .X(_00812_));
 sg13g2_buf_1 _16590_ (.A(\top_ihp.oisc.regs[22][16] ),
    .X(_00813_));
 sg13g2_buf_1 _16591_ (.A(\top_ihp.oisc.regs[22][17] ),
    .X(_00814_));
 sg13g2_buf_1 _16592_ (.A(\top_ihp.oisc.regs[22][18] ),
    .X(_00815_));
 sg13g2_buf_1 _16593_ (.A(\top_ihp.oisc.regs[22][19] ),
    .X(_00816_));
 sg13g2_buf_1 _16594_ (.A(\top_ihp.oisc.regs[22][1] ),
    .X(_00817_));
 sg13g2_buf_1 _16595_ (.A(\top_ihp.oisc.regs[22][20] ),
    .X(_00818_));
 sg13g2_buf_1 _16596_ (.A(\top_ihp.oisc.regs[22][21] ),
    .X(_00819_));
 sg13g2_buf_1 _16597_ (.A(\top_ihp.oisc.regs[22][22] ),
    .X(_00820_));
 sg13g2_buf_1 _16598_ (.A(\top_ihp.oisc.regs[22][23] ),
    .X(_00821_));
 sg13g2_buf_1 _16599_ (.A(\top_ihp.oisc.regs[22][24] ),
    .X(_00822_));
 sg13g2_buf_1 _16600_ (.A(\top_ihp.oisc.regs[22][25] ),
    .X(_00823_));
 sg13g2_buf_1 _16601_ (.A(\top_ihp.oisc.regs[22][26] ),
    .X(_00824_));
 sg13g2_buf_1 _16602_ (.A(\top_ihp.oisc.regs[22][27] ),
    .X(_00825_));
 sg13g2_buf_1 _16603_ (.A(\top_ihp.oisc.regs[22][28] ),
    .X(_00826_));
 sg13g2_buf_1 _16604_ (.A(\top_ihp.oisc.regs[22][29] ),
    .X(_00827_));
 sg13g2_buf_1 _16605_ (.A(\top_ihp.oisc.regs[22][2] ),
    .X(_00828_));
 sg13g2_buf_1 _16606_ (.A(\top_ihp.oisc.regs[22][30] ),
    .X(_00829_));
 sg13g2_buf_1 _16607_ (.A(\top_ihp.oisc.regs[22][31] ),
    .X(_00830_));
 sg13g2_buf_1 _16608_ (.A(\top_ihp.oisc.regs[22][3] ),
    .X(_00831_));
 sg13g2_buf_1 _16609_ (.A(\top_ihp.oisc.regs[22][4] ),
    .X(_00832_));
 sg13g2_buf_1 _16610_ (.A(\top_ihp.oisc.regs[22][5] ),
    .X(_00833_));
 sg13g2_buf_1 _16611_ (.A(\top_ihp.oisc.regs[22][6] ),
    .X(_00834_));
 sg13g2_buf_1 _16612_ (.A(\top_ihp.oisc.regs[22][7] ),
    .X(_00835_));
 sg13g2_buf_1 _16613_ (.A(\top_ihp.oisc.regs[22][8] ),
    .X(_00836_));
 sg13g2_buf_1 _16614_ (.A(\top_ihp.oisc.regs[22][9] ),
    .X(_00837_));
 sg13g2_buf_1 _16615_ (.A(\top_ihp.oisc.regs[23][0] ),
    .X(_00838_));
 sg13g2_buf_1 _16616_ (.A(\top_ihp.oisc.regs[23][10] ),
    .X(_00839_));
 sg13g2_buf_1 _16617_ (.A(\top_ihp.oisc.regs[23][11] ),
    .X(_00840_));
 sg13g2_buf_1 _16618_ (.A(\top_ihp.oisc.regs[23][12] ),
    .X(_00841_));
 sg13g2_buf_1 _16619_ (.A(\top_ihp.oisc.regs[23][13] ),
    .X(_00842_));
 sg13g2_buf_1 _16620_ (.A(\top_ihp.oisc.regs[23][14] ),
    .X(_00843_));
 sg13g2_buf_1 _16621_ (.A(\top_ihp.oisc.regs[23][15] ),
    .X(_00844_));
 sg13g2_buf_1 _16622_ (.A(\top_ihp.oisc.regs[23][16] ),
    .X(_00845_));
 sg13g2_buf_1 _16623_ (.A(\top_ihp.oisc.regs[23][17] ),
    .X(_00846_));
 sg13g2_buf_1 _16624_ (.A(\top_ihp.oisc.regs[23][18] ),
    .X(_00847_));
 sg13g2_buf_1 _16625_ (.A(\top_ihp.oisc.regs[23][19] ),
    .X(_00848_));
 sg13g2_buf_1 _16626_ (.A(\top_ihp.oisc.regs[23][1] ),
    .X(_00849_));
 sg13g2_buf_1 _16627_ (.A(\top_ihp.oisc.regs[23][20] ),
    .X(_00850_));
 sg13g2_buf_1 _16628_ (.A(\top_ihp.oisc.regs[23][21] ),
    .X(_00851_));
 sg13g2_buf_1 _16629_ (.A(\top_ihp.oisc.regs[23][22] ),
    .X(_00852_));
 sg13g2_buf_1 _16630_ (.A(\top_ihp.oisc.regs[23][23] ),
    .X(_00853_));
 sg13g2_buf_1 _16631_ (.A(\top_ihp.oisc.regs[23][24] ),
    .X(_00854_));
 sg13g2_buf_1 _16632_ (.A(\top_ihp.oisc.regs[23][25] ),
    .X(_00855_));
 sg13g2_buf_1 _16633_ (.A(\top_ihp.oisc.regs[23][26] ),
    .X(_00856_));
 sg13g2_buf_1 _16634_ (.A(\top_ihp.oisc.regs[23][27] ),
    .X(_00857_));
 sg13g2_buf_1 _16635_ (.A(\top_ihp.oisc.regs[23][28] ),
    .X(_00858_));
 sg13g2_buf_1 _16636_ (.A(\top_ihp.oisc.regs[23][29] ),
    .X(_00859_));
 sg13g2_buf_1 _16637_ (.A(\top_ihp.oisc.regs[23][2] ),
    .X(_00860_));
 sg13g2_buf_1 _16638_ (.A(\top_ihp.oisc.regs[23][30] ),
    .X(_00861_));
 sg13g2_buf_1 _16639_ (.A(\top_ihp.oisc.regs[23][31] ),
    .X(_00862_));
 sg13g2_buf_1 _16640_ (.A(\top_ihp.oisc.regs[23][3] ),
    .X(_00863_));
 sg13g2_buf_1 _16641_ (.A(\top_ihp.oisc.regs[23][4] ),
    .X(_00864_));
 sg13g2_buf_1 _16642_ (.A(\top_ihp.oisc.regs[23][5] ),
    .X(_00865_));
 sg13g2_buf_1 _16643_ (.A(\top_ihp.oisc.regs[23][6] ),
    .X(_00866_));
 sg13g2_buf_1 _16644_ (.A(\top_ihp.oisc.regs[23][7] ),
    .X(_00867_));
 sg13g2_buf_1 _16645_ (.A(\top_ihp.oisc.regs[23][8] ),
    .X(_00868_));
 sg13g2_buf_1 _16646_ (.A(\top_ihp.oisc.regs[23][9] ),
    .X(_00869_));
 sg13g2_buf_1 _16647_ (.A(\top_ihp.oisc.regs[24][0] ),
    .X(_00870_));
 sg13g2_buf_1 _16648_ (.A(\top_ihp.oisc.regs[24][10] ),
    .X(_00871_));
 sg13g2_buf_1 _16649_ (.A(\top_ihp.oisc.regs[24][11] ),
    .X(_00872_));
 sg13g2_buf_1 _16650_ (.A(\top_ihp.oisc.regs[24][12] ),
    .X(_00873_));
 sg13g2_buf_1 _16651_ (.A(\top_ihp.oisc.regs[24][13] ),
    .X(_00874_));
 sg13g2_buf_1 _16652_ (.A(\top_ihp.oisc.regs[24][14] ),
    .X(_00875_));
 sg13g2_buf_1 _16653_ (.A(\top_ihp.oisc.regs[24][15] ),
    .X(_00876_));
 sg13g2_buf_1 _16654_ (.A(\top_ihp.oisc.regs[24][16] ),
    .X(_00877_));
 sg13g2_buf_1 _16655_ (.A(\top_ihp.oisc.regs[24][17] ),
    .X(_00878_));
 sg13g2_buf_1 _16656_ (.A(\top_ihp.oisc.regs[24][18] ),
    .X(_00879_));
 sg13g2_buf_1 _16657_ (.A(\top_ihp.oisc.regs[24][19] ),
    .X(_00880_));
 sg13g2_buf_1 _16658_ (.A(\top_ihp.oisc.regs[24][1] ),
    .X(_00881_));
 sg13g2_buf_1 _16659_ (.A(\top_ihp.oisc.regs[24][20] ),
    .X(_00882_));
 sg13g2_buf_1 _16660_ (.A(\top_ihp.oisc.regs[24][21] ),
    .X(_00883_));
 sg13g2_buf_1 _16661_ (.A(\top_ihp.oisc.regs[24][22] ),
    .X(_00884_));
 sg13g2_buf_1 _16662_ (.A(\top_ihp.oisc.regs[24][23] ),
    .X(_00885_));
 sg13g2_buf_1 _16663_ (.A(\top_ihp.oisc.regs[24][24] ),
    .X(_00886_));
 sg13g2_buf_1 _16664_ (.A(\top_ihp.oisc.regs[24][25] ),
    .X(_00887_));
 sg13g2_buf_1 _16665_ (.A(\top_ihp.oisc.regs[24][26] ),
    .X(_00888_));
 sg13g2_buf_1 _16666_ (.A(\top_ihp.oisc.regs[24][27] ),
    .X(_00889_));
 sg13g2_buf_1 _16667_ (.A(\top_ihp.oisc.regs[24][28] ),
    .X(_00890_));
 sg13g2_buf_1 _16668_ (.A(\top_ihp.oisc.regs[24][29] ),
    .X(_00891_));
 sg13g2_buf_1 _16669_ (.A(\top_ihp.oisc.regs[24][2] ),
    .X(_00892_));
 sg13g2_buf_1 _16670_ (.A(\top_ihp.oisc.regs[24][30] ),
    .X(_00893_));
 sg13g2_buf_1 _16671_ (.A(\top_ihp.oisc.regs[24][31] ),
    .X(_00894_));
 sg13g2_buf_1 _16672_ (.A(\top_ihp.oisc.regs[24][3] ),
    .X(_00895_));
 sg13g2_buf_1 _16673_ (.A(\top_ihp.oisc.regs[24][4] ),
    .X(_00896_));
 sg13g2_buf_1 _16674_ (.A(\top_ihp.oisc.regs[24][5] ),
    .X(_00897_));
 sg13g2_buf_1 _16675_ (.A(\top_ihp.oisc.regs[24][6] ),
    .X(_00898_));
 sg13g2_buf_1 _16676_ (.A(\top_ihp.oisc.regs[24][7] ),
    .X(_00899_));
 sg13g2_buf_1 _16677_ (.A(\top_ihp.oisc.regs[24][8] ),
    .X(_00900_));
 sg13g2_buf_1 _16678_ (.A(\top_ihp.oisc.regs[24][9] ),
    .X(_00901_));
 sg13g2_buf_1 _16679_ (.A(\top_ihp.oisc.regs[25][0] ),
    .X(_00902_));
 sg13g2_buf_1 _16680_ (.A(\top_ihp.oisc.regs[25][10] ),
    .X(_00903_));
 sg13g2_buf_1 _16681_ (.A(\top_ihp.oisc.regs[25][11] ),
    .X(_00904_));
 sg13g2_buf_1 _16682_ (.A(\top_ihp.oisc.regs[25][12] ),
    .X(_00905_));
 sg13g2_buf_1 _16683_ (.A(\top_ihp.oisc.regs[25][13] ),
    .X(_00906_));
 sg13g2_buf_1 _16684_ (.A(\top_ihp.oisc.regs[25][14] ),
    .X(_00907_));
 sg13g2_buf_1 _16685_ (.A(\top_ihp.oisc.regs[25][15] ),
    .X(_00908_));
 sg13g2_buf_1 _16686_ (.A(\top_ihp.oisc.regs[25][16] ),
    .X(_00909_));
 sg13g2_buf_1 _16687_ (.A(\top_ihp.oisc.regs[25][17] ),
    .X(_00910_));
 sg13g2_buf_1 _16688_ (.A(\top_ihp.oisc.regs[25][18] ),
    .X(_00911_));
 sg13g2_buf_1 _16689_ (.A(\top_ihp.oisc.regs[25][19] ),
    .X(_00912_));
 sg13g2_buf_1 _16690_ (.A(\top_ihp.oisc.regs[25][1] ),
    .X(_00913_));
 sg13g2_buf_1 _16691_ (.A(\top_ihp.oisc.regs[25][20] ),
    .X(_00914_));
 sg13g2_buf_1 _16692_ (.A(\top_ihp.oisc.regs[25][21] ),
    .X(_00915_));
 sg13g2_buf_1 _16693_ (.A(\top_ihp.oisc.regs[25][22] ),
    .X(_00916_));
 sg13g2_buf_1 _16694_ (.A(\top_ihp.oisc.regs[25][23] ),
    .X(_00917_));
 sg13g2_buf_1 _16695_ (.A(\top_ihp.oisc.regs[25][24] ),
    .X(_00918_));
 sg13g2_buf_1 _16696_ (.A(\top_ihp.oisc.regs[25][25] ),
    .X(_00919_));
 sg13g2_buf_1 _16697_ (.A(\top_ihp.oisc.regs[25][26] ),
    .X(_00920_));
 sg13g2_buf_1 _16698_ (.A(\top_ihp.oisc.regs[25][27] ),
    .X(_00921_));
 sg13g2_buf_1 _16699_ (.A(\top_ihp.oisc.regs[25][28] ),
    .X(_00922_));
 sg13g2_buf_1 _16700_ (.A(\top_ihp.oisc.regs[25][29] ),
    .X(_00923_));
 sg13g2_buf_1 _16701_ (.A(\top_ihp.oisc.regs[25][2] ),
    .X(_00924_));
 sg13g2_buf_1 _16702_ (.A(\top_ihp.oisc.regs[25][30] ),
    .X(_00925_));
 sg13g2_buf_1 _16703_ (.A(\top_ihp.oisc.regs[25][31] ),
    .X(_00926_));
 sg13g2_buf_1 _16704_ (.A(\top_ihp.oisc.regs[25][3] ),
    .X(_00927_));
 sg13g2_buf_1 _16705_ (.A(\top_ihp.oisc.regs[25][4] ),
    .X(_00928_));
 sg13g2_buf_1 _16706_ (.A(\top_ihp.oisc.regs[25][5] ),
    .X(_00929_));
 sg13g2_buf_1 _16707_ (.A(\top_ihp.oisc.regs[25][6] ),
    .X(_00930_));
 sg13g2_buf_1 _16708_ (.A(\top_ihp.oisc.regs[25][7] ),
    .X(_00931_));
 sg13g2_buf_1 _16709_ (.A(\top_ihp.oisc.regs[25][8] ),
    .X(_00932_));
 sg13g2_buf_1 _16710_ (.A(\top_ihp.oisc.regs[25][9] ),
    .X(_00933_));
 sg13g2_buf_1 _16711_ (.A(\top_ihp.oisc.regs[26][0] ),
    .X(_00934_));
 sg13g2_buf_1 _16712_ (.A(\top_ihp.oisc.regs[26][10] ),
    .X(_00935_));
 sg13g2_buf_1 _16713_ (.A(\top_ihp.oisc.regs[26][11] ),
    .X(_00936_));
 sg13g2_buf_1 _16714_ (.A(\top_ihp.oisc.regs[26][12] ),
    .X(_00937_));
 sg13g2_buf_1 _16715_ (.A(\top_ihp.oisc.regs[26][13] ),
    .X(_00938_));
 sg13g2_buf_1 _16716_ (.A(\top_ihp.oisc.regs[26][14] ),
    .X(_00939_));
 sg13g2_buf_1 _16717_ (.A(\top_ihp.oisc.regs[26][15] ),
    .X(_00940_));
 sg13g2_buf_1 _16718_ (.A(\top_ihp.oisc.regs[26][16] ),
    .X(_00941_));
 sg13g2_buf_1 _16719_ (.A(\top_ihp.oisc.regs[26][17] ),
    .X(_00942_));
 sg13g2_buf_1 _16720_ (.A(\top_ihp.oisc.regs[26][18] ),
    .X(_00943_));
 sg13g2_buf_1 _16721_ (.A(\top_ihp.oisc.regs[26][19] ),
    .X(_00944_));
 sg13g2_buf_1 _16722_ (.A(\top_ihp.oisc.regs[26][1] ),
    .X(_00945_));
 sg13g2_buf_1 _16723_ (.A(\top_ihp.oisc.regs[26][20] ),
    .X(_00946_));
 sg13g2_buf_1 _16724_ (.A(\top_ihp.oisc.regs[26][21] ),
    .X(_00947_));
 sg13g2_buf_1 _16725_ (.A(\top_ihp.oisc.regs[26][22] ),
    .X(_00948_));
 sg13g2_buf_1 _16726_ (.A(\top_ihp.oisc.regs[26][23] ),
    .X(_00949_));
 sg13g2_buf_1 _16727_ (.A(\top_ihp.oisc.regs[26][24] ),
    .X(_00950_));
 sg13g2_buf_1 _16728_ (.A(\top_ihp.oisc.regs[26][25] ),
    .X(_00951_));
 sg13g2_buf_1 _16729_ (.A(\top_ihp.oisc.regs[26][26] ),
    .X(_00952_));
 sg13g2_buf_1 _16730_ (.A(\top_ihp.oisc.regs[26][27] ),
    .X(_00953_));
 sg13g2_buf_1 _16731_ (.A(\top_ihp.oisc.regs[26][28] ),
    .X(_00954_));
 sg13g2_buf_1 _16732_ (.A(\top_ihp.oisc.regs[26][29] ),
    .X(_00955_));
 sg13g2_buf_1 _16733_ (.A(\top_ihp.oisc.regs[26][2] ),
    .X(_00956_));
 sg13g2_buf_1 _16734_ (.A(\top_ihp.oisc.regs[26][30] ),
    .X(_00957_));
 sg13g2_buf_1 _16735_ (.A(\top_ihp.oisc.regs[26][31] ),
    .X(_00958_));
 sg13g2_buf_1 _16736_ (.A(\top_ihp.oisc.regs[26][3] ),
    .X(_00959_));
 sg13g2_buf_1 _16737_ (.A(\top_ihp.oisc.regs[26][4] ),
    .X(_00960_));
 sg13g2_buf_1 _16738_ (.A(\top_ihp.oisc.regs[26][5] ),
    .X(_00961_));
 sg13g2_buf_1 _16739_ (.A(\top_ihp.oisc.regs[26][6] ),
    .X(_00962_));
 sg13g2_buf_1 _16740_ (.A(\top_ihp.oisc.regs[26][7] ),
    .X(_00963_));
 sg13g2_buf_1 _16741_ (.A(\top_ihp.oisc.regs[26][8] ),
    .X(_00964_));
 sg13g2_buf_1 _16742_ (.A(\top_ihp.oisc.regs[26][9] ),
    .X(_00965_));
 sg13g2_buf_1 _16743_ (.A(\top_ihp.oisc.regs[27][0] ),
    .X(_00966_));
 sg13g2_buf_1 _16744_ (.A(\top_ihp.oisc.regs[27][10] ),
    .X(_00967_));
 sg13g2_buf_1 _16745_ (.A(\top_ihp.oisc.regs[27][11] ),
    .X(_00968_));
 sg13g2_buf_1 _16746_ (.A(\top_ihp.oisc.regs[27][12] ),
    .X(_00969_));
 sg13g2_buf_1 _16747_ (.A(\top_ihp.oisc.regs[27][13] ),
    .X(_00970_));
 sg13g2_buf_1 _16748_ (.A(\top_ihp.oisc.regs[27][14] ),
    .X(_00971_));
 sg13g2_buf_1 _16749_ (.A(\top_ihp.oisc.regs[27][15] ),
    .X(_00972_));
 sg13g2_buf_1 _16750_ (.A(\top_ihp.oisc.regs[27][16] ),
    .X(_00973_));
 sg13g2_buf_1 _16751_ (.A(\top_ihp.oisc.regs[27][17] ),
    .X(_00974_));
 sg13g2_buf_1 _16752_ (.A(\top_ihp.oisc.regs[27][18] ),
    .X(_00975_));
 sg13g2_buf_1 _16753_ (.A(\top_ihp.oisc.regs[27][19] ),
    .X(_00976_));
 sg13g2_buf_1 _16754_ (.A(\top_ihp.oisc.regs[27][1] ),
    .X(_00977_));
 sg13g2_buf_1 _16755_ (.A(\top_ihp.oisc.regs[27][20] ),
    .X(_00978_));
 sg13g2_buf_1 _16756_ (.A(\top_ihp.oisc.regs[27][21] ),
    .X(_00979_));
 sg13g2_buf_1 _16757_ (.A(\top_ihp.oisc.regs[27][22] ),
    .X(_00980_));
 sg13g2_buf_1 _16758_ (.A(\top_ihp.oisc.regs[27][23] ),
    .X(_00981_));
 sg13g2_buf_1 _16759_ (.A(\top_ihp.oisc.regs[27][24] ),
    .X(_00982_));
 sg13g2_buf_1 _16760_ (.A(\top_ihp.oisc.regs[27][25] ),
    .X(_00983_));
 sg13g2_buf_1 _16761_ (.A(\top_ihp.oisc.regs[27][26] ),
    .X(_00984_));
 sg13g2_buf_1 _16762_ (.A(\top_ihp.oisc.regs[27][27] ),
    .X(_00985_));
 sg13g2_buf_1 _16763_ (.A(\top_ihp.oisc.regs[27][28] ),
    .X(_00986_));
 sg13g2_buf_1 _16764_ (.A(\top_ihp.oisc.regs[27][29] ),
    .X(_00987_));
 sg13g2_buf_1 _16765_ (.A(\top_ihp.oisc.regs[27][2] ),
    .X(_00988_));
 sg13g2_buf_1 _16766_ (.A(\top_ihp.oisc.regs[27][30] ),
    .X(_00989_));
 sg13g2_buf_1 _16767_ (.A(\top_ihp.oisc.regs[27][31] ),
    .X(_00990_));
 sg13g2_buf_1 _16768_ (.A(\top_ihp.oisc.regs[27][3] ),
    .X(_00991_));
 sg13g2_buf_1 _16769_ (.A(\top_ihp.oisc.regs[27][4] ),
    .X(_00992_));
 sg13g2_buf_1 _16770_ (.A(\top_ihp.oisc.regs[27][5] ),
    .X(_00993_));
 sg13g2_buf_1 _16771_ (.A(\top_ihp.oisc.regs[27][6] ),
    .X(_00994_));
 sg13g2_buf_1 _16772_ (.A(\top_ihp.oisc.regs[27][7] ),
    .X(_00995_));
 sg13g2_buf_1 _16773_ (.A(\top_ihp.oisc.regs[27][8] ),
    .X(_00996_));
 sg13g2_buf_1 _16774_ (.A(\top_ihp.oisc.regs[27][9] ),
    .X(_00997_));
 sg13g2_buf_1 _16775_ (.A(\top_ihp.oisc.regs[28][0] ),
    .X(_00998_));
 sg13g2_buf_1 _16776_ (.A(\top_ihp.oisc.regs[28][10] ),
    .X(_00999_));
 sg13g2_buf_1 _16777_ (.A(\top_ihp.oisc.regs[28][11] ),
    .X(_01000_));
 sg13g2_buf_1 _16778_ (.A(\top_ihp.oisc.regs[28][12] ),
    .X(_01001_));
 sg13g2_buf_1 _16779_ (.A(\top_ihp.oisc.regs[28][13] ),
    .X(_01002_));
 sg13g2_buf_1 _16780_ (.A(\top_ihp.oisc.regs[28][14] ),
    .X(_01003_));
 sg13g2_buf_1 _16781_ (.A(\top_ihp.oisc.regs[28][15] ),
    .X(_01004_));
 sg13g2_buf_1 _16782_ (.A(\top_ihp.oisc.regs[28][16] ),
    .X(_01005_));
 sg13g2_buf_1 _16783_ (.A(\top_ihp.oisc.regs[28][17] ),
    .X(_01006_));
 sg13g2_buf_1 _16784_ (.A(\top_ihp.oisc.regs[28][18] ),
    .X(_01007_));
 sg13g2_buf_1 _16785_ (.A(\top_ihp.oisc.regs[28][19] ),
    .X(_01008_));
 sg13g2_buf_1 _16786_ (.A(\top_ihp.oisc.regs[28][1] ),
    .X(_01009_));
 sg13g2_buf_1 _16787_ (.A(\top_ihp.oisc.regs[28][20] ),
    .X(_01010_));
 sg13g2_buf_1 _16788_ (.A(\top_ihp.oisc.regs[28][21] ),
    .X(_01011_));
 sg13g2_buf_1 _16789_ (.A(\top_ihp.oisc.regs[28][22] ),
    .X(_01012_));
 sg13g2_buf_1 _16790_ (.A(\top_ihp.oisc.regs[28][23] ),
    .X(_01013_));
 sg13g2_buf_1 _16791_ (.A(\top_ihp.oisc.regs[28][24] ),
    .X(_01014_));
 sg13g2_buf_1 _16792_ (.A(\top_ihp.oisc.regs[28][25] ),
    .X(_01015_));
 sg13g2_buf_1 _16793_ (.A(\top_ihp.oisc.regs[28][26] ),
    .X(_01016_));
 sg13g2_buf_1 _16794_ (.A(\top_ihp.oisc.regs[28][27] ),
    .X(_01017_));
 sg13g2_buf_1 _16795_ (.A(\top_ihp.oisc.regs[28][28] ),
    .X(_01018_));
 sg13g2_buf_1 _16796_ (.A(\top_ihp.oisc.regs[28][29] ),
    .X(_01019_));
 sg13g2_buf_1 _16797_ (.A(\top_ihp.oisc.regs[28][2] ),
    .X(_01020_));
 sg13g2_buf_1 _16798_ (.A(\top_ihp.oisc.regs[28][30] ),
    .X(_01021_));
 sg13g2_buf_1 _16799_ (.A(\top_ihp.oisc.regs[28][31] ),
    .X(_01022_));
 sg13g2_buf_1 _16800_ (.A(\top_ihp.oisc.regs[28][3] ),
    .X(_01023_));
 sg13g2_buf_1 _16801_ (.A(\top_ihp.oisc.regs[28][4] ),
    .X(_01024_));
 sg13g2_buf_1 _16802_ (.A(\top_ihp.oisc.regs[28][5] ),
    .X(_01025_));
 sg13g2_buf_1 _16803_ (.A(\top_ihp.oisc.regs[28][6] ),
    .X(_01026_));
 sg13g2_buf_1 _16804_ (.A(\top_ihp.oisc.regs[28][7] ),
    .X(_01027_));
 sg13g2_buf_1 _16805_ (.A(\top_ihp.oisc.regs[28][8] ),
    .X(_01028_));
 sg13g2_buf_1 _16806_ (.A(\top_ihp.oisc.regs[28][9] ),
    .X(_01029_));
 sg13g2_buf_1 _16807_ (.A(\top_ihp.oisc.regs[29][0] ),
    .X(_01030_));
 sg13g2_buf_1 _16808_ (.A(\top_ihp.oisc.regs[29][10] ),
    .X(_01031_));
 sg13g2_buf_1 _16809_ (.A(\top_ihp.oisc.regs[29][11] ),
    .X(_01032_));
 sg13g2_buf_1 _16810_ (.A(\top_ihp.oisc.regs[29][12] ),
    .X(_01033_));
 sg13g2_buf_1 _16811_ (.A(\top_ihp.oisc.regs[29][13] ),
    .X(_01034_));
 sg13g2_buf_1 _16812_ (.A(\top_ihp.oisc.regs[29][14] ),
    .X(_01035_));
 sg13g2_buf_1 _16813_ (.A(\top_ihp.oisc.regs[29][15] ),
    .X(_01036_));
 sg13g2_buf_1 _16814_ (.A(\top_ihp.oisc.regs[29][16] ),
    .X(_01037_));
 sg13g2_buf_1 _16815_ (.A(\top_ihp.oisc.regs[29][17] ),
    .X(_01038_));
 sg13g2_buf_1 _16816_ (.A(\top_ihp.oisc.regs[29][18] ),
    .X(_01039_));
 sg13g2_buf_1 _16817_ (.A(\top_ihp.oisc.regs[29][19] ),
    .X(_01040_));
 sg13g2_buf_1 _16818_ (.A(\top_ihp.oisc.regs[29][1] ),
    .X(_01041_));
 sg13g2_buf_1 _16819_ (.A(\top_ihp.oisc.regs[29][20] ),
    .X(_01042_));
 sg13g2_buf_1 _16820_ (.A(\top_ihp.oisc.regs[29][21] ),
    .X(_01043_));
 sg13g2_buf_1 _16821_ (.A(\top_ihp.oisc.regs[29][22] ),
    .X(_01044_));
 sg13g2_buf_1 _16822_ (.A(\top_ihp.oisc.regs[29][23] ),
    .X(_01045_));
 sg13g2_buf_1 _16823_ (.A(\top_ihp.oisc.regs[29][24] ),
    .X(_01046_));
 sg13g2_buf_1 _16824_ (.A(\top_ihp.oisc.regs[29][25] ),
    .X(_01047_));
 sg13g2_buf_1 _16825_ (.A(\top_ihp.oisc.regs[29][26] ),
    .X(_01048_));
 sg13g2_buf_1 _16826_ (.A(\top_ihp.oisc.regs[29][27] ),
    .X(_01049_));
 sg13g2_buf_1 _16827_ (.A(\top_ihp.oisc.regs[29][28] ),
    .X(_01050_));
 sg13g2_buf_1 _16828_ (.A(\top_ihp.oisc.regs[29][29] ),
    .X(_01051_));
 sg13g2_buf_1 _16829_ (.A(\top_ihp.oisc.regs[29][2] ),
    .X(_01052_));
 sg13g2_buf_1 _16830_ (.A(\top_ihp.oisc.regs[29][30] ),
    .X(_01053_));
 sg13g2_buf_1 _16831_ (.A(\top_ihp.oisc.regs[29][31] ),
    .X(_01054_));
 sg13g2_buf_1 _16832_ (.A(\top_ihp.oisc.regs[29][3] ),
    .X(_01055_));
 sg13g2_buf_1 _16833_ (.A(\top_ihp.oisc.regs[29][4] ),
    .X(_01056_));
 sg13g2_buf_1 _16834_ (.A(\top_ihp.oisc.regs[29][5] ),
    .X(_01057_));
 sg13g2_buf_1 _16835_ (.A(\top_ihp.oisc.regs[29][6] ),
    .X(_01058_));
 sg13g2_buf_1 _16836_ (.A(\top_ihp.oisc.regs[29][7] ),
    .X(_01059_));
 sg13g2_buf_1 _16837_ (.A(\top_ihp.oisc.regs[29][8] ),
    .X(_01060_));
 sg13g2_buf_1 _16838_ (.A(\top_ihp.oisc.regs[29][9] ),
    .X(_01061_));
 sg13g2_and2_1 _16839_ (.A(_09106_),
    .B(net711),
    .X(_10232_));
 sg13g2_buf_1 _16840_ (.A(_10232_),
    .X(_10233_));
 sg13g2_mux2_1 _16841_ (.A0(\top_ihp.oisc.regs[2][0] ),
    .A1(net210),
    .S(_10233_),
    .X(_01062_));
 sg13g2_nand2_1 _16842_ (.Y(_10234_),
    .A(_09106_),
    .B(net711));
 sg13g2_buf_1 _16843_ (.A(_10234_),
    .X(_10235_));
 sg13g2_buf_1 _16844_ (.A(_10235_),
    .X(_10236_));
 sg13g2_buf_1 _16845_ (.A(net531),
    .X(_10237_));
 sg13g2_buf_1 _16846_ (.A(_10235_),
    .X(_10238_));
 sg13g2_nand2_1 _16847_ (.Y(_10239_),
    .A(\top_ihp.oisc.regs[2][10] ),
    .B(net530));
 sg13g2_o21ai_1 _16848_ (.B1(_10239_),
    .Y(_01063_),
    .A1(net74),
    .A2(net395));
 sg13g2_buf_1 _16849_ (.A(_10235_),
    .X(_10240_));
 sg13g2_nand2_1 _16850_ (.Y(_10241_),
    .A(\top_ihp.oisc.regs[2][11] ),
    .B(net529));
 sg13g2_o21ai_1 _16851_ (.B1(_10241_),
    .Y(_01064_),
    .A1(net148),
    .A2(net395));
 sg13g2_nand2_1 _16852_ (.Y(_10242_),
    .A(\top_ihp.oisc.regs[2][12] ),
    .B(net529));
 sg13g2_o21ai_1 _16853_ (.B1(_10242_),
    .Y(_01065_),
    .A1(net250),
    .A2(net395));
 sg13g2_nand2_1 _16854_ (.Y(_10243_),
    .A(\top_ihp.oisc.regs[2][13] ),
    .B(_10240_));
 sg13g2_o21ai_1 _16855_ (.B1(_10243_),
    .Y(_01066_),
    .A1(net58),
    .A2(_10237_));
 sg13g2_nand2_1 _16856_ (.Y(_10244_),
    .A(\top_ihp.oisc.regs[2][14] ),
    .B(net529));
 sg13g2_o21ai_1 _16857_ (.B1(_10244_),
    .Y(_01067_),
    .A1(net249),
    .A2(net395));
 sg13g2_nand2_1 _16858_ (.Y(_10245_),
    .A(\top_ihp.oisc.regs[2][15] ),
    .B(net529));
 sg13g2_o21ai_1 _16859_ (.B1(_10245_),
    .Y(_01068_),
    .A1(_09419_),
    .A2(net395));
 sg13g2_nand2_1 _16860_ (.Y(_10246_),
    .A(\top_ihp.oisc.regs[2][16] ),
    .B(_10240_));
 sg13g2_o21ai_1 _16861_ (.B1(_10246_),
    .Y(_01069_),
    .A1(net130),
    .A2(_10237_));
 sg13g2_nand2_1 _16862_ (.Y(_10247_),
    .A(\top_ihp.oisc.regs[2][17] ),
    .B(net529));
 sg13g2_o21ai_1 _16863_ (.B1(_10247_),
    .Y(_01070_),
    .A1(_09462_),
    .A2(net395));
 sg13g2_nand2_1 _16864_ (.Y(_10248_),
    .A(\top_ihp.oisc.regs[2][18] ),
    .B(net529));
 sg13g2_o21ai_1 _16865_ (.B1(_10248_),
    .Y(_01071_),
    .A1(net144),
    .A2(net395));
 sg13g2_nand2_1 _16866_ (.Y(_10249_),
    .A(\top_ihp.oisc.regs[2][19] ),
    .B(net529));
 sg13g2_o21ai_1 _16867_ (.B1(_10249_),
    .Y(_01072_),
    .A1(_09512_),
    .A2(net395));
 sg13g2_buf_1 _16868_ (.A(net531),
    .X(_10250_));
 sg13g2_nand2_1 _16869_ (.Y(_10251_),
    .A(\top_ihp.oisc.regs[2][1] ),
    .B(net529));
 sg13g2_o21ai_1 _16870_ (.B1(_10251_),
    .Y(_01073_),
    .A1(net409),
    .A2(net394));
 sg13g2_nor2_1 _16871_ (.A(\top_ihp.oisc.regs[2][20] ),
    .B(_10233_),
    .Y(_10252_));
 sg13g2_a21oi_1 _16872_ (.A1(net40),
    .A2(_10233_),
    .Y(_01074_),
    .B1(_10252_));
 sg13g2_buf_1 _16873_ (.A(_10235_),
    .X(_10253_));
 sg13g2_nand2_1 _16874_ (.Y(_10254_),
    .A(\top_ihp.oisc.regs[2][21] ),
    .B(net528));
 sg13g2_o21ai_1 _16875_ (.B1(_10254_),
    .Y(_01075_),
    .A1(net72),
    .A2(_10250_));
 sg13g2_nand2_1 _16876_ (.Y(_10255_),
    .A(\top_ihp.oisc.regs[2][22] ),
    .B(net528));
 sg13g2_o21ai_1 _16877_ (.B1(_10255_),
    .Y(_01076_),
    .A1(net129),
    .A2(net394));
 sg13g2_nor2_1 _16878_ (.A(\top_ihp.oisc.regs[2][23] ),
    .B(_10233_),
    .Y(_10256_));
 sg13g2_a21oi_1 _16879_ (.A1(net138),
    .A2(_10233_),
    .Y(_01077_),
    .B1(_10256_));
 sg13g2_nand2_1 _16880_ (.Y(_10257_),
    .A(\top_ihp.oisc.regs[2][24] ),
    .B(_10253_));
 sg13g2_o21ai_1 _16881_ (.B1(_10257_),
    .Y(_01078_),
    .A1(net242),
    .A2(net394));
 sg13g2_nand2_1 _16882_ (.Y(_10258_),
    .A(\top_ihp.oisc.regs[2][25] ),
    .B(_10253_));
 sg13g2_o21ai_1 _16883_ (.B1(_10258_),
    .Y(_01079_),
    .A1(net241),
    .A2(_10250_));
 sg13g2_nand2_1 _16884_ (.Y(_10259_),
    .A(\top_ihp.oisc.regs[2][26] ),
    .B(net528));
 sg13g2_o21ai_1 _16885_ (.B1(_10259_),
    .Y(_01080_),
    .A1(net142),
    .A2(net394));
 sg13g2_nand2_1 _16886_ (.Y(_10260_),
    .A(\top_ihp.oisc.regs[2][27] ),
    .B(net528));
 sg13g2_o21ai_1 _16887_ (.B1(_10260_),
    .Y(_01081_),
    .A1(net71),
    .A2(net394));
 sg13g2_nand2_1 _16888_ (.Y(_10261_),
    .A(\top_ihp.oisc.regs[2][28] ),
    .B(net528));
 sg13g2_o21ai_1 _16889_ (.B1(_10261_),
    .Y(_01082_),
    .A1(net70),
    .A2(net394));
 sg13g2_nand2_1 _16890_ (.Y(_10262_),
    .A(\top_ihp.oisc.regs[2][29] ),
    .B(net528));
 sg13g2_o21ai_1 _16891_ (.B1(_10262_),
    .Y(_01083_),
    .A1(net140),
    .A2(net394));
 sg13g2_nand2_1 _16892_ (.Y(_10263_),
    .A(\top_ihp.oisc.regs[2][2] ),
    .B(net528));
 sg13g2_o21ai_1 _16893_ (.B1(_10263_),
    .Y(_01084_),
    .A1(net240),
    .A2(net394));
 sg13g2_nand2_1 _16894_ (.Y(_10264_),
    .A(\top_ihp.oisc.regs[2][30] ),
    .B(net528));
 sg13g2_o21ai_1 _16895_ (.B1(_10264_),
    .Y(_01085_),
    .A1(net69),
    .A2(net530));
 sg13g2_nand2_1 _16896_ (.Y(_10265_),
    .A(\top_ihp.oisc.regs[2][31] ),
    .B(_10236_));
 sg13g2_o21ai_1 _16897_ (.B1(_10265_),
    .Y(_01086_),
    .A1(net139),
    .A2(_10238_));
 sg13g2_nand2_1 _16898_ (.Y(_10266_),
    .A(\top_ihp.oisc.regs[2][3] ),
    .B(net531));
 sg13g2_o21ai_1 _16899_ (.B1(_10266_),
    .Y(_01087_),
    .A1(net238),
    .A2(net530));
 sg13g2_nand2_1 _16900_ (.Y(_10267_),
    .A(\top_ihp.oisc.regs[2][4] ),
    .B(_10236_));
 sg13g2_o21ai_1 _16901_ (.B1(_10267_),
    .Y(_01088_),
    .A1(net237),
    .A2(_10238_));
 sg13g2_nand2_1 _16902_ (.Y(_10268_),
    .A(\top_ihp.oisc.regs[2][5] ),
    .B(net531));
 sg13g2_o21ai_1 _16903_ (.B1(_10268_),
    .Y(_01089_),
    .A1(net236),
    .A2(net530));
 sg13g2_nand2_1 _16904_ (.Y(_10269_),
    .A(\top_ihp.oisc.regs[2][6] ),
    .B(net531));
 sg13g2_o21ai_1 _16905_ (.B1(_10269_),
    .Y(_01090_),
    .A1(net235),
    .A2(net530));
 sg13g2_nand2_1 _16906_ (.Y(_10270_),
    .A(\top_ihp.oisc.regs[2][7] ),
    .B(net531));
 sg13g2_o21ai_1 _16907_ (.B1(_10270_),
    .Y(_01091_),
    .A1(net68),
    .A2(net530));
 sg13g2_nand2_1 _16908_ (.Y(_10271_),
    .A(\top_ihp.oisc.regs[2][8] ),
    .B(net531));
 sg13g2_o21ai_1 _16909_ (.B1(_10271_),
    .Y(_01092_),
    .A1(net67),
    .A2(net530));
 sg13g2_nand2_1 _16910_ (.Y(_10272_),
    .A(\top_ihp.oisc.regs[2][9] ),
    .B(net531));
 sg13g2_o21ai_1 _16911_ (.B1(_10272_),
    .Y(_01093_),
    .A1(net66),
    .A2(net530));
 sg13g2_buf_1 _16912_ (.A(\top_ihp.oisc.regs[30][0] ),
    .X(_01094_));
 sg13g2_buf_1 _16913_ (.A(\top_ihp.oisc.regs[30][10] ),
    .X(_01095_));
 sg13g2_buf_1 _16914_ (.A(\top_ihp.oisc.regs[30][11] ),
    .X(_01096_));
 sg13g2_buf_1 _16915_ (.A(\top_ihp.oisc.regs[30][12] ),
    .X(_01097_));
 sg13g2_buf_1 _16916_ (.A(\top_ihp.oisc.regs[30][13] ),
    .X(_01098_));
 sg13g2_buf_1 _16917_ (.A(\top_ihp.oisc.regs[30][14] ),
    .X(_01099_));
 sg13g2_buf_1 _16918_ (.A(\top_ihp.oisc.regs[30][15] ),
    .X(_01100_));
 sg13g2_buf_1 _16919_ (.A(\top_ihp.oisc.regs[30][16] ),
    .X(_01101_));
 sg13g2_buf_1 _16920_ (.A(\top_ihp.oisc.regs[30][17] ),
    .X(_01102_));
 sg13g2_buf_1 _16921_ (.A(\top_ihp.oisc.regs[30][18] ),
    .X(_01103_));
 sg13g2_buf_1 _16922_ (.A(\top_ihp.oisc.regs[30][19] ),
    .X(_01104_));
 sg13g2_buf_1 _16923_ (.A(\top_ihp.oisc.regs[30][1] ),
    .X(_01105_));
 sg13g2_buf_1 _16924_ (.A(\top_ihp.oisc.regs[30][20] ),
    .X(_01106_));
 sg13g2_buf_1 _16925_ (.A(\top_ihp.oisc.regs[30][21] ),
    .X(_01107_));
 sg13g2_buf_1 _16926_ (.A(\top_ihp.oisc.regs[30][22] ),
    .X(_01108_));
 sg13g2_buf_1 _16927_ (.A(\top_ihp.oisc.regs[30][23] ),
    .X(_01109_));
 sg13g2_buf_1 _16928_ (.A(\top_ihp.oisc.regs[30][24] ),
    .X(_01110_));
 sg13g2_buf_1 _16929_ (.A(\top_ihp.oisc.regs[30][25] ),
    .X(_01111_));
 sg13g2_buf_1 _16930_ (.A(\top_ihp.oisc.regs[30][26] ),
    .X(_01112_));
 sg13g2_buf_1 _16931_ (.A(\top_ihp.oisc.regs[30][27] ),
    .X(_01113_));
 sg13g2_buf_1 _16932_ (.A(\top_ihp.oisc.regs[30][28] ),
    .X(_01114_));
 sg13g2_buf_1 _16933_ (.A(\top_ihp.oisc.regs[30][29] ),
    .X(_01115_));
 sg13g2_buf_1 _16934_ (.A(\top_ihp.oisc.regs[30][2] ),
    .X(_01116_));
 sg13g2_buf_1 _16935_ (.A(\top_ihp.oisc.regs[30][30] ),
    .X(_01117_));
 sg13g2_buf_1 _16936_ (.A(\top_ihp.oisc.regs[30][31] ),
    .X(_01118_));
 sg13g2_buf_1 _16937_ (.A(\top_ihp.oisc.regs[30][3] ),
    .X(_01119_));
 sg13g2_buf_1 _16938_ (.A(\top_ihp.oisc.regs[30][4] ),
    .X(_01120_));
 sg13g2_buf_1 _16939_ (.A(\top_ihp.oisc.regs[30][5] ),
    .X(_01121_));
 sg13g2_buf_1 _16940_ (.A(\top_ihp.oisc.regs[30][6] ),
    .X(_01122_));
 sg13g2_buf_1 _16941_ (.A(\top_ihp.oisc.regs[30][7] ),
    .X(_01123_));
 sg13g2_buf_1 _16942_ (.A(\top_ihp.oisc.regs[30][8] ),
    .X(_01124_));
 sg13g2_buf_1 _16943_ (.A(\top_ihp.oisc.regs[30][9] ),
    .X(_01125_));
 sg13g2_buf_1 _16944_ (.A(\top_ihp.oisc.regs[31][0] ),
    .X(_01126_));
 sg13g2_buf_1 _16945_ (.A(\top_ihp.oisc.regs[31][10] ),
    .X(_01127_));
 sg13g2_buf_1 _16946_ (.A(\top_ihp.oisc.regs[31][11] ),
    .X(_01128_));
 sg13g2_buf_1 _16947_ (.A(\top_ihp.oisc.regs[31][12] ),
    .X(_01129_));
 sg13g2_buf_1 _16948_ (.A(\top_ihp.oisc.regs[31][13] ),
    .X(_01130_));
 sg13g2_buf_1 _16949_ (.A(\top_ihp.oisc.regs[31][14] ),
    .X(_01131_));
 sg13g2_buf_1 _16950_ (.A(\top_ihp.oisc.regs[31][15] ),
    .X(_01132_));
 sg13g2_buf_1 _16951_ (.A(\top_ihp.oisc.regs[31][16] ),
    .X(_01133_));
 sg13g2_buf_1 _16952_ (.A(\top_ihp.oisc.regs[31][17] ),
    .X(_01134_));
 sg13g2_buf_1 _16953_ (.A(\top_ihp.oisc.regs[31][18] ),
    .X(_01135_));
 sg13g2_buf_1 _16954_ (.A(\top_ihp.oisc.regs[31][19] ),
    .X(_01136_));
 sg13g2_buf_1 _16955_ (.A(\top_ihp.oisc.regs[31][1] ),
    .X(_01137_));
 sg13g2_buf_1 _16956_ (.A(\top_ihp.oisc.regs[31][20] ),
    .X(_01138_));
 sg13g2_buf_1 _16957_ (.A(\top_ihp.oisc.regs[31][21] ),
    .X(_01139_));
 sg13g2_buf_1 _16958_ (.A(\top_ihp.oisc.regs[31][22] ),
    .X(_01140_));
 sg13g2_buf_1 _16959_ (.A(\top_ihp.oisc.regs[31][23] ),
    .X(_01141_));
 sg13g2_buf_1 _16960_ (.A(\top_ihp.oisc.regs[31][24] ),
    .X(_01142_));
 sg13g2_buf_1 _16961_ (.A(\top_ihp.oisc.regs[31][25] ),
    .X(_01143_));
 sg13g2_buf_1 _16962_ (.A(\top_ihp.oisc.regs[31][26] ),
    .X(_01144_));
 sg13g2_buf_1 _16963_ (.A(\top_ihp.oisc.regs[31][27] ),
    .X(_01145_));
 sg13g2_buf_1 _16964_ (.A(\top_ihp.oisc.regs[31][28] ),
    .X(_01146_));
 sg13g2_buf_1 _16965_ (.A(\top_ihp.oisc.regs[31][29] ),
    .X(_01147_));
 sg13g2_buf_1 _16966_ (.A(\top_ihp.oisc.regs[31][2] ),
    .X(_01148_));
 sg13g2_buf_1 _16967_ (.A(\top_ihp.oisc.regs[31][30] ),
    .X(_01149_));
 sg13g2_buf_1 _16968_ (.A(\top_ihp.oisc.regs[31][31] ),
    .X(_01150_));
 sg13g2_buf_1 _16969_ (.A(\top_ihp.oisc.regs[31][3] ),
    .X(_01151_));
 sg13g2_buf_1 _16970_ (.A(\top_ihp.oisc.regs[31][4] ),
    .X(_01152_));
 sg13g2_buf_1 _16971_ (.A(\top_ihp.oisc.regs[31][5] ),
    .X(_01153_));
 sg13g2_buf_1 _16972_ (.A(\top_ihp.oisc.regs[31][6] ),
    .X(_01154_));
 sg13g2_buf_1 _16973_ (.A(\top_ihp.oisc.regs[31][7] ),
    .X(_01155_));
 sg13g2_buf_1 _16974_ (.A(\top_ihp.oisc.regs[31][8] ),
    .X(_01156_));
 sg13g2_buf_1 _16975_ (.A(\top_ihp.oisc.regs[31][9] ),
    .X(_01157_));
 sg13g2_buf_1 _16976_ (.A(\top_ihp.oisc.regs[32][0] ),
    .X(_01158_));
 sg13g2_buf_1 _16977_ (.A(\top_ihp.oisc.regs[32][10] ),
    .X(_01159_));
 sg13g2_buf_1 _16978_ (.A(\top_ihp.oisc.regs[32][11] ),
    .X(_01160_));
 sg13g2_buf_1 _16979_ (.A(\top_ihp.oisc.regs[32][12] ),
    .X(_01161_));
 sg13g2_buf_1 _16980_ (.A(\top_ihp.oisc.regs[32][13] ),
    .X(_01162_));
 sg13g2_buf_1 _16981_ (.A(\top_ihp.oisc.regs[32][14] ),
    .X(_01163_));
 sg13g2_buf_1 _16982_ (.A(\top_ihp.oisc.regs[32][15] ),
    .X(_01164_));
 sg13g2_buf_1 _16983_ (.A(\top_ihp.oisc.regs[32][16] ),
    .X(_01165_));
 sg13g2_buf_1 _16984_ (.A(\top_ihp.oisc.regs[32][17] ),
    .X(_01166_));
 sg13g2_buf_1 _16985_ (.A(\top_ihp.oisc.regs[32][18] ),
    .X(_01167_));
 sg13g2_buf_1 _16986_ (.A(\top_ihp.oisc.regs[32][19] ),
    .X(_01168_));
 sg13g2_buf_1 _16987_ (.A(\top_ihp.oisc.regs[32][1] ),
    .X(_01169_));
 sg13g2_buf_1 _16988_ (.A(\top_ihp.oisc.regs[32][20] ),
    .X(_01170_));
 sg13g2_buf_1 _16989_ (.A(\top_ihp.oisc.regs[32][21] ),
    .X(_01171_));
 sg13g2_buf_1 _16990_ (.A(\top_ihp.oisc.regs[32][22] ),
    .X(_01172_));
 sg13g2_buf_1 _16991_ (.A(\top_ihp.oisc.regs[32][23] ),
    .X(_01173_));
 sg13g2_buf_1 _16992_ (.A(\top_ihp.oisc.regs[32][24] ),
    .X(_01174_));
 sg13g2_buf_1 _16993_ (.A(\top_ihp.oisc.regs[32][25] ),
    .X(_01175_));
 sg13g2_buf_1 _16994_ (.A(\top_ihp.oisc.regs[32][26] ),
    .X(_01176_));
 sg13g2_buf_1 _16995_ (.A(\top_ihp.oisc.regs[32][27] ),
    .X(_01177_));
 sg13g2_buf_1 _16996_ (.A(\top_ihp.oisc.regs[32][28] ),
    .X(_01178_));
 sg13g2_buf_1 _16997_ (.A(\top_ihp.oisc.regs[32][29] ),
    .X(_01179_));
 sg13g2_buf_1 _16998_ (.A(\top_ihp.oisc.regs[32][2] ),
    .X(_01180_));
 sg13g2_buf_1 _16999_ (.A(\top_ihp.oisc.regs[32][30] ),
    .X(_01181_));
 sg13g2_buf_1 _17000_ (.A(\top_ihp.oisc.regs[32][31] ),
    .X(_01182_));
 sg13g2_buf_1 _17001_ (.A(\top_ihp.oisc.regs[32][3] ),
    .X(_01183_));
 sg13g2_buf_1 _17002_ (.A(\top_ihp.oisc.regs[32][4] ),
    .X(_01184_));
 sg13g2_buf_1 _17003_ (.A(\top_ihp.oisc.regs[32][5] ),
    .X(_01185_));
 sg13g2_buf_1 _17004_ (.A(\top_ihp.oisc.regs[32][6] ),
    .X(_01186_));
 sg13g2_buf_1 _17005_ (.A(\top_ihp.oisc.regs[32][7] ),
    .X(_01187_));
 sg13g2_buf_1 _17006_ (.A(\top_ihp.oisc.regs[32][8] ),
    .X(_01188_));
 sg13g2_buf_1 _17007_ (.A(\top_ihp.oisc.regs[32][9] ),
    .X(_01189_));
 sg13g2_nor3_1 _17008_ (.A(_09067_),
    .B(_09085_),
    .C(_09093_),
    .Y(_10273_));
 sg13g2_buf_2 _17009_ (.A(_10273_),
    .X(_10274_));
 sg13g2_nand2_1 _17010_ (.Y(_10275_),
    .A(net710),
    .B(_10274_));
 sg13g2_buf_2 _17011_ (.A(_10275_),
    .X(_10276_));
 sg13g2_nor2b_1 _17012_ (.A(_10276_),
    .B_N(net737),
    .Y(_10277_));
 sg13g2_buf_1 _17013_ (.A(_10277_),
    .X(_10278_));
 sg13g2_mux2_1 _17014_ (.A0(\top_ihp.oisc.regs[33][0] ),
    .A1(net210),
    .S(net527),
    .X(_01190_));
 sg13g2_nand3_1 _17015_ (.B(net710),
    .C(_10274_),
    .A(net737),
    .Y(_10279_));
 sg13g2_buf_2 _17016_ (.A(_10279_),
    .X(_10280_));
 sg13g2_buf_1 _17017_ (.A(_10280_),
    .X(_10281_));
 sg13g2_buf_1 _17018_ (.A(_10280_),
    .X(_10282_));
 sg13g2_nand2_1 _17019_ (.Y(_10283_),
    .A(\top_ihp.oisc.regs[33][10] ),
    .B(net636));
 sg13g2_o21ai_1 _17020_ (.B1(_10283_),
    .Y(_01191_),
    .A1(_09270_),
    .A2(net637));
 sg13g2_nand2_1 _17021_ (.Y(_10284_),
    .A(\top_ihp.oisc.regs[33][11] ),
    .B(net636));
 sg13g2_o21ai_1 _17022_ (.B1(_10284_),
    .Y(_01192_),
    .A1(net148),
    .A2(net637));
 sg13g2_nand2_1 _17023_ (.Y(_10285_),
    .A(\top_ihp.oisc.regs[33][12] ),
    .B(net636));
 sg13g2_o21ai_1 _17024_ (.B1(_10285_),
    .Y(_01193_),
    .A1(_09348_),
    .A2(net637));
 sg13g2_nor2_1 _17025_ (.A(\top_ihp.oisc.regs[33][13] ),
    .B(net527),
    .Y(_10286_));
 sg13g2_a21oi_1 _17026_ (.A1(net59),
    .A2(net527),
    .Y(_01194_),
    .B1(_10286_));
 sg13g2_nand2_1 _17027_ (.Y(_10287_),
    .A(\top_ihp.oisc.regs[33][14] ),
    .B(net636));
 sg13g2_o21ai_1 _17028_ (.B1(_10287_),
    .Y(_01195_),
    .A1(_09404_),
    .A2(net637));
 sg13g2_buf_1 _17029_ (.A(_10280_),
    .X(_10288_));
 sg13g2_nand2_1 _17030_ (.Y(_10289_),
    .A(\top_ihp.oisc.regs[33][15] ),
    .B(net635));
 sg13g2_o21ai_1 _17031_ (.B1(_10289_),
    .Y(_01196_),
    .A1(_09419_),
    .A2(net637));
 sg13g2_nor2_1 _17032_ (.A(\top_ihp.oisc.regs[33][16] ),
    .B(net527),
    .Y(_10290_));
 sg13g2_a21oi_1 _17033_ (.A1(_10122_),
    .A2(net527),
    .Y(_01197_),
    .B1(_10290_));
 sg13g2_nand2_1 _17034_ (.Y(_10291_),
    .A(\top_ihp.oisc.regs[33][17] ),
    .B(net635));
 sg13g2_o21ai_1 _17035_ (.B1(_10291_),
    .Y(_01198_),
    .A1(_09462_),
    .A2(net637));
 sg13g2_nand2_1 _17036_ (.Y(_10292_),
    .A(\top_ihp.oisc.regs[33][18] ),
    .B(net635));
 sg13g2_o21ai_1 _17037_ (.B1(_10292_),
    .Y(_01199_),
    .A1(_09483_),
    .A2(net637));
 sg13g2_nand2_1 _17038_ (.Y(_10293_),
    .A(\top_ihp.oisc.regs[33][19] ),
    .B(net635));
 sg13g2_o21ai_1 _17039_ (.B1(_10293_),
    .Y(_01200_),
    .A1(_09512_),
    .A2(net637));
 sg13g2_nand2_1 _17040_ (.Y(_10294_),
    .A(\top_ihp.oisc.regs[33][1] ),
    .B(_10288_));
 sg13g2_o21ai_1 _17041_ (.B1(_10294_),
    .Y(_01201_),
    .A1(_09554_),
    .A2(_10281_));
 sg13g2_nor2_1 _17042_ (.A(\top_ihp.oisc.regs[33][20] ),
    .B(net527),
    .Y(_10295_));
 sg13g2_a21oi_1 _17043_ (.A1(net40),
    .A2(net527),
    .Y(_01202_),
    .B1(_10295_));
 sg13g2_nand2_1 _17044_ (.Y(_10296_),
    .A(\top_ihp.oisc.regs[33][21] ),
    .B(net635));
 sg13g2_o21ai_1 _17045_ (.B1(_10296_),
    .Y(_01203_),
    .A1(_09599_),
    .A2(_10281_));
 sg13g2_nor2_1 _17046_ (.A(\top_ihp.oisc.regs[33][22] ),
    .B(_10278_),
    .Y(_10297_));
 sg13g2_a21oi_1 _17047_ (.A1(net131),
    .A2(_10278_),
    .Y(_01204_),
    .B1(_10297_));
 sg13g2_nor2_1 _17048_ (.A(\top_ihp.oisc.regs[33][23] ),
    .B(_10277_),
    .Y(_10298_));
 sg13g2_a21oi_1 _17049_ (.A1(_09986_),
    .A2(net527),
    .Y(_01205_),
    .B1(_10298_));
 sg13g2_buf_1 _17050_ (.A(_10280_),
    .X(_10299_));
 sg13g2_nand2_1 _17051_ (.Y(_10300_),
    .A(\top_ihp.oisc.regs[33][24] ),
    .B(net635));
 sg13g2_o21ai_1 _17052_ (.B1(_10300_),
    .Y(_01206_),
    .A1(_09654_),
    .A2(net634));
 sg13g2_nand2_1 _17053_ (.Y(_10301_),
    .A(\top_ihp.oisc.regs[33][25] ),
    .B(_10288_));
 sg13g2_o21ai_1 _17054_ (.B1(_10301_),
    .Y(_01207_),
    .A1(_09669_),
    .A2(_10299_));
 sg13g2_nand2_1 _17055_ (.Y(_10302_),
    .A(\top_ihp.oisc.regs[33][26] ),
    .B(net635));
 sg13g2_o21ai_1 _17056_ (.B1(_10302_),
    .Y(_01208_),
    .A1(net142),
    .A2(net634));
 sg13g2_nand2_1 _17057_ (.Y(_10303_),
    .A(\top_ihp.oisc.regs[33][27] ),
    .B(net635));
 sg13g2_o21ai_1 _17058_ (.B1(_10303_),
    .Y(_01209_),
    .A1(net71),
    .A2(_10299_));
 sg13g2_buf_1 _17059_ (.A(_10280_),
    .X(_10304_));
 sg13g2_nand2_1 _17060_ (.Y(_10305_),
    .A(\top_ihp.oisc.regs[33][28] ),
    .B(net633));
 sg13g2_o21ai_1 _17061_ (.B1(_10305_),
    .Y(_01210_),
    .A1(net70),
    .A2(net634));
 sg13g2_nand2_1 _17062_ (.Y(_10306_),
    .A(\top_ihp.oisc.regs[33][29] ),
    .B(net633));
 sg13g2_o21ai_1 _17063_ (.B1(_10306_),
    .Y(_01211_),
    .A1(net140),
    .A2(net634));
 sg13g2_nand2_1 _17064_ (.Y(_10307_),
    .A(\top_ihp.oisc.regs[33][2] ),
    .B(net633));
 sg13g2_o21ai_1 _17065_ (.B1(_10307_),
    .Y(_01212_),
    .A1(_09754_),
    .A2(net634));
 sg13g2_nand2_1 _17066_ (.Y(_10308_),
    .A(\top_ihp.oisc.regs[33][30] ),
    .B(net633));
 sg13g2_o21ai_1 _17067_ (.B1(_10308_),
    .Y(_01213_),
    .A1(net69),
    .A2(net634));
 sg13g2_nand2_1 _17068_ (.Y(_10309_),
    .A(\top_ihp.oisc.regs[33][31] ),
    .B(_10304_));
 sg13g2_o21ai_1 _17069_ (.B1(_10309_),
    .Y(_01214_),
    .A1(net139),
    .A2(net634));
 sg13g2_nand2_1 _17070_ (.Y(_10310_),
    .A(\top_ihp.oisc.regs[33][3] ),
    .B(_10304_));
 sg13g2_o21ai_1 _17071_ (.B1(_10310_),
    .Y(_01215_),
    .A1(net238),
    .A2(net634));
 sg13g2_nand2_1 _17072_ (.Y(_10311_),
    .A(\top_ihp.oisc.regs[33][4] ),
    .B(net633));
 sg13g2_o21ai_1 _17073_ (.B1(_10311_),
    .Y(_01216_),
    .A1(net237),
    .A2(net636));
 sg13g2_nand2_1 _17074_ (.Y(_10312_),
    .A(\top_ihp.oisc.regs[33][5] ),
    .B(net633));
 sg13g2_o21ai_1 _17075_ (.B1(_10312_),
    .Y(_01217_),
    .A1(_09872_),
    .A2(_10282_));
 sg13g2_nand2_1 _17076_ (.Y(_10313_),
    .A(\top_ihp.oisc.regs[33][6] ),
    .B(net633));
 sg13g2_o21ai_1 _17077_ (.B1(_10313_),
    .Y(_01218_),
    .A1(_09895_),
    .A2(_10282_));
 sg13g2_nand2_1 _17078_ (.Y(_10314_),
    .A(\top_ihp.oisc.regs[33][7] ),
    .B(net633));
 sg13g2_o21ai_1 _17079_ (.B1(_10314_),
    .Y(_01219_),
    .A1(net209),
    .A2(net636));
 sg13g2_nand2_1 _17080_ (.Y(_10315_),
    .A(\top_ihp.oisc.regs[33][8] ),
    .B(_10280_));
 sg13g2_o21ai_1 _17081_ (.B1(_10315_),
    .Y(_01220_),
    .A1(net67),
    .A2(net636));
 sg13g2_nand2_1 _17082_ (.Y(_10316_),
    .A(\top_ihp.oisc.regs[33][9] ),
    .B(_10280_));
 sg13g2_o21ai_1 _17083_ (.B1(_10316_),
    .Y(_01221_),
    .A1(net66),
    .A2(net636));
 sg13g2_and2_1 _17084_ (.A(_09960_),
    .B(_10274_),
    .X(_10317_));
 sg13g2_buf_1 _17085_ (.A(_10317_),
    .X(_10318_));
 sg13g2_and2_1 _17086_ (.A(net737),
    .B(_10318_),
    .X(_10319_));
 sg13g2_buf_2 _17087_ (.A(_10319_),
    .X(_10320_));
 sg13g2_mux2_1 _17088_ (.A0(\top_ihp.oisc.regs[34][0] ),
    .A1(net210),
    .S(_10320_),
    .X(_01222_));
 sg13g2_nand2_1 _17089_ (.Y(_10321_),
    .A(net737),
    .B(net664));
 sg13g2_buf_1 _17090_ (.A(_10321_),
    .X(_10322_));
 sg13g2_buf_1 _17091_ (.A(net526),
    .X(_10323_));
 sg13g2_buf_1 _17092_ (.A(net526),
    .X(_10324_));
 sg13g2_nand2_1 _17093_ (.Y(_10325_),
    .A(\top_ihp.oisc.regs[34][10] ),
    .B(net392));
 sg13g2_o21ai_1 _17094_ (.B1(_10325_),
    .Y(_01223_),
    .A1(net74),
    .A2(net393));
 sg13g2_nand2_1 _17095_ (.Y(_10326_),
    .A(\top_ihp.oisc.regs[34][11] ),
    .B(net392));
 sg13g2_o21ai_1 _17096_ (.B1(_10326_),
    .Y(_01224_),
    .A1(_09304_),
    .A2(net393));
 sg13g2_nand2_1 _17097_ (.Y(_10327_),
    .A(\top_ihp.oisc.regs[34][12] ),
    .B(net392));
 sg13g2_o21ai_1 _17098_ (.B1(_10327_),
    .Y(_01225_),
    .A1(net250),
    .A2(_10323_));
 sg13g2_buf_1 _17099_ (.A(net526),
    .X(_10328_));
 sg13g2_nand2_1 _17100_ (.Y(_10329_),
    .A(\top_ihp.oisc.regs[34][13] ),
    .B(net391));
 sg13g2_o21ai_1 _17101_ (.B1(_10329_),
    .Y(_01226_),
    .A1(net58),
    .A2(net393));
 sg13g2_nand2_1 _17102_ (.Y(_10330_),
    .A(\top_ihp.oisc.regs[34][14] ),
    .B(net391));
 sg13g2_o21ai_1 _17103_ (.B1(_10330_),
    .Y(_01227_),
    .A1(_09404_),
    .A2(net393));
 sg13g2_mux2_1 _17104_ (.A0(_00210_),
    .A1(net216),
    .S(_10320_),
    .X(_01228_));
 sg13g2_nand2_1 _17105_ (.Y(_10331_),
    .A(\top_ihp.oisc.regs[34][16] ),
    .B(net391));
 sg13g2_o21ai_1 _17106_ (.B1(_10331_),
    .Y(_01229_),
    .A1(net130),
    .A2(net393));
 sg13g2_nand2_1 _17107_ (.Y(_10332_),
    .A(\top_ihp.oisc.regs[34][17] ),
    .B(net391));
 sg13g2_o21ai_1 _17108_ (.B1(_10332_),
    .Y(_01230_),
    .A1(net145),
    .A2(net393));
 sg13g2_nand2_1 _17109_ (.Y(_10333_),
    .A(\top_ihp.oisc.regs[34][18] ),
    .B(_10328_));
 sg13g2_o21ai_1 _17110_ (.B1(_10333_),
    .Y(_01231_),
    .A1(net144),
    .A2(net393));
 sg13g2_nand2_1 _17111_ (.Y(_10334_),
    .A(\top_ihp.oisc.regs[34][19] ),
    .B(net391));
 sg13g2_o21ai_1 _17112_ (.B1(_10334_),
    .Y(_01232_),
    .A1(net246),
    .A2(net393));
 sg13g2_nand2_1 _17113_ (.Y(_10335_),
    .A(\top_ihp.oisc.regs[34][1] ),
    .B(net391));
 sg13g2_o21ai_1 _17114_ (.B1(_10335_),
    .Y(_01233_),
    .A1(_09554_),
    .A2(_10323_));
 sg13g2_nor2_1 _17115_ (.A(\top_ihp.oisc.regs[34][20] ),
    .B(_10320_),
    .Y(_10336_));
 sg13g2_a21oi_1 _17116_ (.A1(net40),
    .A2(_10320_),
    .Y(_01234_),
    .B1(_10336_));
 sg13g2_buf_1 _17117_ (.A(net526),
    .X(_10337_));
 sg13g2_nand2_1 _17118_ (.Y(_10338_),
    .A(\top_ihp.oisc.regs[34][21] ),
    .B(_10328_));
 sg13g2_o21ai_1 _17119_ (.B1(_10338_),
    .Y(_01235_),
    .A1(net72),
    .A2(net390));
 sg13g2_nand2_1 _17120_ (.Y(_10339_),
    .A(\top_ihp.oisc.regs[34][22] ),
    .B(net391));
 sg13g2_o21ai_1 _17121_ (.B1(_10339_),
    .Y(_01236_),
    .A1(_10214_),
    .A2(net390));
 sg13g2_nor2_1 _17122_ (.A(\top_ihp.oisc.regs[34][23] ),
    .B(_10320_),
    .Y(_10340_));
 sg13g2_a21oi_1 _17123_ (.A1(net138),
    .A2(_10320_),
    .Y(_01237_),
    .B1(_10340_));
 sg13g2_nand2_1 _17124_ (.Y(_10341_),
    .A(\top_ihp.oisc.regs[34][24] ),
    .B(net391));
 sg13g2_o21ai_1 _17125_ (.B1(_10341_),
    .Y(_01238_),
    .A1(net242),
    .A2(net390));
 sg13g2_buf_1 _17126_ (.A(net526),
    .X(_10342_));
 sg13g2_nand2_1 _17127_ (.Y(_10343_),
    .A(\top_ihp.oisc.regs[34][25] ),
    .B(net389));
 sg13g2_o21ai_1 _17128_ (.B1(_10343_),
    .Y(_01239_),
    .A1(net241),
    .A2(net390));
 sg13g2_nand2_1 _17129_ (.Y(_10344_),
    .A(\top_ihp.oisc.regs[34][26] ),
    .B(net389));
 sg13g2_o21ai_1 _17130_ (.B1(_10344_),
    .Y(_01240_),
    .A1(_09679_),
    .A2(net390));
 sg13g2_nand2_1 _17131_ (.Y(_10345_),
    .A(\top_ihp.oisc.regs[34][27] ),
    .B(net389));
 sg13g2_o21ai_1 _17132_ (.B1(_10345_),
    .Y(_01241_),
    .A1(_09703_),
    .A2(_10337_));
 sg13g2_nand2_1 _17133_ (.Y(_10346_),
    .A(\top_ihp.oisc.regs[34][28] ),
    .B(_10342_));
 sg13g2_o21ai_1 _17134_ (.B1(_10346_),
    .Y(_01242_),
    .A1(_09714_),
    .A2(_10337_));
 sg13g2_nand2_1 _17135_ (.Y(_10347_),
    .A(\top_ihp.oisc.regs[34][29] ),
    .B(_10342_));
 sg13g2_o21ai_1 _17136_ (.B1(_10347_),
    .Y(_01243_),
    .A1(_09724_),
    .A2(net390));
 sg13g2_nand2_1 _17137_ (.Y(_10348_),
    .A(\top_ihp.oisc.regs[34][2] ),
    .B(net389));
 sg13g2_o21ai_1 _17138_ (.B1(_10348_),
    .Y(_01244_),
    .A1(net240),
    .A2(net390));
 sg13g2_nand2_1 _17139_ (.Y(_10349_),
    .A(\top_ihp.oisc.regs[34][30] ),
    .B(net389));
 sg13g2_o21ai_1 _17140_ (.B1(_10349_),
    .Y(_01245_),
    .A1(net69),
    .A2(net390));
 sg13g2_mux2_1 _17141_ (.A0(_00211_),
    .A1(net239),
    .S(_10320_),
    .X(_01246_));
 sg13g2_nand2_1 _17142_ (.Y(_10350_),
    .A(\top_ihp.oisc.regs[34][3] ),
    .B(net389));
 sg13g2_o21ai_1 _17143_ (.B1(_10350_),
    .Y(_01247_),
    .A1(net238),
    .A2(net392));
 sg13g2_nand2_1 _17144_ (.Y(_10351_),
    .A(\top_ihp.oisc.regs[34][4] ),
    .B(net389));
 sg13g2_o21ai_1 _17145_ (.B1(_10351_),
    .Y(_01248_),
    .A1(net237),
    .A2(net392));
 sg13g2_nand2_1 _17146_ (.Y(_10352_),
    .A(\top_ihp.oisc.regs[34][5] ),
    .B(net389));
 sg13g2_o21ai_1 _17147_ (.B1(_10352_),
    .Y(_01249_),
    .A1(net236),
    .A2(net392));
 sg13g2_nand2_1 _17148_ (.Y(_10353_),
    .A(\top_ihp.oisc.regs[34][6] ),
    .B(net526));
 sg13g2_o21ai_1 _17149_ (.B1(_10353_),
    .Y(_01250_),
    .A1(net235),
    .A2(net392));
 sg13g2_nand2_1 _17150_ (.Y(_10354_),
    .A(\top_ihp.oisc.regs[34][7] ),
    .B(net526));
 sg13g2_o21ai_1 _17151_ (.B1(_10354_),
    .Y(_01251_),
    .A1(net68),
    .A2(_10324_));
 sg13g2_nand2_1 _17152_ (.Y(_10355_),
    .A(\top_ihp.oisc.regs[34][8] ),
    .B(_10322_));
 sg13g2_o21ai_1 _17153_ (.B1(_10355_),
    .Y(_01252_),
    .A1(_09930_),
    .A2(_10324_));
 sg13g2_nand2_1 _17154_ (.Y(_10356_),
    .A(\top_ihp.oisc.regs[34][9] ),
    .B(net526));
 sg13g2_o21ai_1 _17155_ (.B1(_10356_),
    .Y(_01253_),
    .A1(_09944_),
    .A2(net392));
 sg13g2_and2_1 _17156_ (.A(_10009_),
    .B(_10274_),
    .X(_10357_));
 sg13g2_buf_2 _17157_ (.A(_10357_),
    .X(_10358_));
 sg13g2_and2_1 _17158_ (.A(net737),
    .B(_10358_),
    .X(_10359_));
 sg13g2_buf_2 _17159_ (.A(_10359_),
    .X(_10360_));
 sg13g2_mux2_1 _17160_ (.A0(\top_ihp.oisc.regs[35][0] ),
    .A1(net210),
    .S(_10360_),
    .X(_01254_));
 sg13g2_nand2_1 _17161_ (.Y(_10361_),
    .A(net737),
    .B(_10358_));
 sg13g2_buf_1 _17162_ (.A(_10361_),
    .X(_10362_));
 sg13g2_buf_1 _17163_ (.A(net525),
    .X(_10363_));
 sg13g2_buf_1 _17164_ (.A(net525),
    .X(_10364_));
 sg13g2_nand2_1 _17165_ (.Y(_10365_),
    .A(\top_ihp.oisc.regs[35][10] ),
    .B(net387));
 sg13g2_o21ai_1 _17166_ (.B1(_10365_),
    .Y(_01255_),
    .A1(_09270_),
    .A2(_10363_));
 sg13g2_nor2_1 _17167_ (.A(_00212_),
    .B(_10360_),
    .Y(_10366_));
 sg13g2_a21oi_1 _17168_ (.A1(_09301_),
    .A2(_10360_),
    .Y(_01256_),
    .B1(_10366_));
 sg13g2_nand2_1 _17169_ (.Y(_10367_),
    .A(\top_ihp.oisc.regs[35][12] ),
    .B(net387));
 sg13g2_o21ai_1 _17170_ (.B1(_10367_),
    .Y(_01257_),
    .A1(_09348_),
    .A2(net388));
 sg13g2_nand2_1 _17171_ (.Y(_10368_),
    .A(\top_ihp.oisc.regs[35][13] ),
    .B(net387));
 sg13g2_o21ai_1 _17172_ (.B1(_10368_),
    .Y(_01258_),
    .A1(net58),
    .A2(net388));
 sg13g2_buf_1 _17173_ (.A(net525),
    .X(_10369_));
 sg13g2_nand2_1 _17174_ (.Y(_10370_),
    .A(\top_ihp.oisc.regs[35][14] ),
    .B(net386));
 sg13g2_o21ai_1 _17175_ (.B1(_10370_),
    .Y(_01259_),
    .A1(net249),
    .A2(net388));
 sg13g2_nand2_1 _17176_ (.Y(_10371_),
    .A(\top_ihp.oisc.regs[35][15] ),
    .B(net386));
 sg13g2_o21ai_1 _17177_ (.B1(_10371_),
    .Y(_01260_),
    .A1(net248),
    .A2(net388));
 sg13g2_nand2_1 _17178_ (.Y(_10372_),
    .A(\top_ihp.oisc.regs[35][16] ),
    .B(net386));
 sg13g2_o21ai_1 _17179_ (.B1(_10372_),
    .Y(_01261_),
    .A1(net130),
    .A2(net388));
 sg13g2_nand2_1 _17180_ (.Y(_10373_),
    .A(\top_ihp.oisc.regs[35][17] ),
    .B(net386));
 sg13g2_o21ai_1 _17181_ (.B1(_10373_),
    .Y(_01262_),
    .A1(net145),
    .A2(net388));
 sg13g2_nand2_1 _17182_ (.Y(_10374_),
    .A(\top_ihp.oisc.regs[35][18] ),
    .B(net386));
 sg13g2_o21ai_1 _17183_ (.B1(_10374_),
    .Y(_01263_),
    .A1(_09483_),
    .A2(net388));
 sg13g2_nand2_1 _17184_ (.Y(_10375_),
    .A(\top_ihp.oisc.regs[35][19] ),
    .B(net386));
 sg13g2_o21ai_1 _17185_ (.B1(_10375_),
    .Y(_01264_),
    .A1(net246),
    .A2(net388));
 sg13g2_nand2_1 _17186_ (.Y(_10376_),
    .A(\top_ihp.oisc.regs[35][1] ),
    .B(net386));
 sg13g2_o21ai_1 _17187_ (.B1(_10376_),
    .Y(_01265_),
    .A1(net409),
    .A2(_10363_));
 sg13g2_mux2_1 _17188_ (.A0(\top_ihp.oisc.regs[35][20] ),
    .A1(net137),
    .S(_10360_),
    .X(_01266_));
 sg13g2_buf_1 _17189_ (.A(net525),
    .X(_10377_));
 sg13g2_nand2_1 _17190_ (.Y(_10378_),
    .A(\top_ihp.oisc.regs[35][21] ),
    .B(_10369_));
 sg13g2_o21ai_1 _17191_ (.B1(_10378_),
    .Y(_01267_),
    .A1(_09599_),
    .A2(net385));
 sg13g2_nand2_1 _17192_ (.Y(_10379_),
    .A(\top_ihp.oisc.regs[35][22] ),
    .B(_10369_));
 sg13g2_o21ai_1 _17193_ (.B1(_10379_),
    .Y(_01268_),
    .A1(_10214_),
    .A2(net385));
 sg13g2_mux2_1 _17194_ (.A0(\top_ihp.oisc.regs[35][23] ),
    .A1(net224),
    .S(_10360_),
    .X(_01269_));
 sg13g2_nand2_1 _17195_ (.Y(_10380_),
    .A(\top_ihp.oisc.regs[35][24] ),
    .B(net386));
 sg13g2_o21ai_1 _17196_ (.B1(_10380_),
    .Y(_01270_),
    .A1(_09654_),
    .A2(net385));
 sg13g2_buf_1 _17197_ (.A(net525),
    .X(_10381_));
 sg13g2_nand2_1 _17198_ (.Y(_10382_),
    .A(\top_ihp.oisc.regs[35][25] ),
    .B(net384));
 sg13g2_o21ai_1 _17199_ (.B1(_10382_),
    .Y(_01271_),
    .A1(_09669_),
    .A2(net385));
 sg13g2_nand2_1 _17200_ (.Y(_10383_),
    .A(\top_ihp.oisc.regs[35][26] ),
    .B(net384));
 sg13g2_o21ai_1 _17201_ (.B1(_10383_),
    .Y(_01272_),
    .A1(_09679_),
    .A2(net385));
 sg13g2_nand2_1 _17202_ (.Y(_10384_),
    .A(\top_ihp.oisc.regs[35][27] ),
    .B(_10381_));
 sg13g2_o21ai_1 _17203_ (.B1(_10384_),
    .Y(_01273_),
    .A1(_09703_),
    .A2(_10377_));
 sg13g2_nand2_1 _17204_ (.Y(_10385_),
    .A(\top_ihp.oisc.regs[35][28] ),
    .B(_10381_));
 sg13g2_o21ai_1 _17205_ (.B1(_10385_),
    .Y(_01274_),
    .A1(_09714_),
    .A2(net385));
 sg13g2_nand2_1 _17206_ (.Y(_10386_),
    .A(\top_ihp.oisc.regs[35][29] ),
    .B(net384));
 sg13g2_o21ai_1 _17207_ (.B1(_10386_),
    .Y(_01275_),
    .A1(_09724_),
    .A2(net385));
 sg13g2_nand2_1 _17208_ (.Y(_10387_),
    .A(\top_ihp.oisc.regs[35][2] ),
    .B(net384));
 sg13g2_o21ai_1 _17209_ (.B1(_10387_),
    .Y(_01276_),
    .A1(_09754_),
    .A2(net385));
 sg13g2_nand2_1 _17210_ (.Y(_10388_),
    .A(\top_ihp.oisc.regs[35][30] ),
    .B(net384));
 sg13g2_o21ai_1 _17211_ (.B1(_10388_),
    .Y(_01277_),
    .A1(_09762_),
    .A2(_10377_));
 sg13g2_mux2_1 _17212_ (.A0(_00213_),
    .A1(net239),
    .S(_10360_),
    .X(_01278_));
 sg13g2_nand2_1 _17213_ (.Y(_10389_),
    .A(\top_ihp.oisc.regs[35][3] ),
    .B(net384));
 sg13g2_o21ai_1 _17214_ (.B1(_10389_),
    .Y(_01279_),
    .A1(_09808_),
    .A2(net387));
 sg13g2_nand2_1 _17215_ (.Y(_10390_),
    .A(\top_ihp.oisc.regs[35][4] ),
    .B(net384));
 sg13g2_o21ai_1 _17216_ (.B1(_10390_),
    .Y(_01280_),
    .A1(_09841_),
    .A2(net387));
 sg13g2_nand2_1 _17217_ (.Y(_10391_),
    .A(\top_ihp.oisc.regs[35][5] ),
    .B(net384));
 sg13g2_o21ai_1 _17218_ (.B1(_10391_),
    .Y(_01281_),
    .A1(_09872_),
    .A2(net387));
 sg13g2_nand2_1 _17219_ (.Y(_10392_),
    .A(\top_ihp.oisc.regs[35][6] ),
    .B(net525));
 sg13g2_o21ai_1 _17220_ (.B1(_10392_),
    .Y(_01282_),
    .A1(_09895_),
    .A2(_10364_));
 sg13g2_nand2_1 _17221_ (.Y(_10393_),
    .A(\top_ihp.oisc.regs[35][7] ),
    .B(net525));
 sg13g2_o21ai_1 _17222_ (.B1(_10393_),
    .Y(_01283_),
    .A1(net209),
    .A2(net387));
 sg13g2_nand2_1 _17223_ (.Y(_10394_),
    .A(\top_ihp.oisc.regs[35][8] ),
    .B(_10362_));
 sg13g2_o21ai_1 _17224_ (.B1(_10394_),
    .Y(_01284_),
    .A1(_09930_),
    .A2(_10364_));
 sg13g2_nand2_1 _17225_ (.Y(_10395_),
    .A(\top_ihp.oisc.regs[35][9] ),
    .B(net525));
 sg13g2_o21ai_1 _17226_ (.B1(_10395_),
    .Y(_01285_),
    .A1(_09944_),
    .A2(net387));
 sg13g2_nor3_1 _17227_ (.A(_09954_),
    .B(_09950_),
    .C(_09953_),
    .Y(_10396_));
 sg13g2_buf_2 _17228_ (.A(_10396_),
    .X(_10397_));
 sg13g2_buf_1 _17229_ (.A(_10397_),
    .X(_10398_));
 sg13g2_nand2b_1 _17230_ (.Y(_10399_),
    .B(_10274_),
    .A_N(net737));
 sg13g2_nor2_1 _17231_ (.A(_09082_),
    .B(_10399_),
    .Y(_10400_));
 sg13g2_buf_2 _17232_ (.A(_10400_),
    .X(_10401_));
 sg13g2_and2_1 _17233_ (.A(net663),
    .B(_10401_),
    .X(_10402_));
 sg13g2_buf_1 _17234_ (.A(_10402_),
    .X(_10403_));
 sg13g2_mux2_1 _17235_ (.A0(\top_ihp.oisc.regs[36][0] ),
    .A1(net210),
    .S(_10403_),
    .X(_01286_));
 sg13g2_buf_8 _17236_ (.A(net65),
    .X(_10404_));
 sg13g2_nand2_1 _17237_ (.Y(_10405_),
    .A(_10397_),
    .B(_10401_));
 sg13g2_buf_1 _17238_ (.A(_10405_),
    .X(_10406_));
 sg13g2_buf_1 _17239_ (.A(_10406_),
    .X(_10407_));
 sg13g2_buf_2 _17240_ (.A(net383),
    .X(_10408_));
 sg13g2_buf_1 _17241_ (.A(_10406_),
    .X(_10409_));
 sg13g2_nand2_1 _17242_ (.Y(_10410_),
    .A(\top_ihp.oisc.regs[36][10] ),
    .B(net382));
 sg13g2_o21ai_1 _17243_ (.B1(_10410_),
    .Y(_01287_),
    .A1(net39),
    .A2(_10408_));
 sg13g2_buf_1 _17244_ (.A(_10406_),
    .X(_10411_));
 sg13g2_nand2_1 _17245_ (.Y(_10412_),
    .A(\top_ihp.oisc.regs[36][11] ),
    .B(net381));
 sg13g2_o21ai_1 _17246_ (.B1(_10412_),
    .Y(_01288_),
    .A1(_09304_),
    .A2(net208));
 sg13g2_buf_1 _17247_ (.A(net218),
    .X(_10413_));
 sg13g2_nand2_1 _17248_ (.Y(_10414_),
    .A(\top_ihp.oisc.regs[36][12] ),
    .B(_10411_));
 sg13g2_o21ai_1 _17249_ (.B1(_10414_),
    .Y(_01289_),
    .A1(net128),
    .A2(net208));
 sg13g2_nand2_1 _17250_ (.Y(_10415_),
    .A(\top_ihp.oisc.regs[36][13] ),
    .B(net381));
 sg13g2_o21ai_1 _17251_ (.B1(_10415_),
    .Y(_01290_),
    .A1(net58),
    .A2(net208));
 sg13g2_buf_1 _17252_ (.A(net217),
    .X(_10416_));
 sg13g2_nand2_1 _17253_ (.Y(_10417_),
    .A(\top_ihp.oisc.regs[36][14] ),
    .B(_10411_));
 sg13g2_o21ai_1 _17254_ (.B1(_10417_),
    .Y(_01291_),
    .A1(_10416_),
    .A2(_10408_));
 sg13g2_nand2_1 _17255_ (.Y(_10418_),
    .A(\top_ihp.oisc.regs[36][15] ),
    .B(net381));
 sg13g2_o21ai_1 _17256_ (.B1(_10418_),
    .Y(_01292_),
    .A1(net248),
    .A2(net208));
 sg13g2_nand2_1 _17257_ (.Y(_10419_),
    .A(\top_ihp.oisc.regs[36][16] ),
    .B(net381));
 sg13g2_o21ai_1 _17258_ (.B1(_10419_),
    .Y(_01293_),
    .A1(net130),
    .A2(net208));
 sg13g2_buf_1 _17259_ (.A(net136),
    .X(_10420_));
 sg13g2_nand2_1 _17260_ (.Y(_10421_),
    .A(\top_ihp.oisc.regs[36][17] ),
    .B(net381));
 sg13g2_o21ai_1 _17261_ (.B1(_10421_),
    .Y(_01294_),
    .A1(net57),
    .A2(net208));
 sg13g2_buf_1 _17262_ (.A(net135),
    .X(_10422_));
 sg13g2_nand2_1 _17263_ (.Y(_10423_),
    .A(\top_ihp.oisc.regs[36][18] ),
    .B(net381));
 sg13g2_o21ai_1 _17264_ (.B1(_10423_),
    .Y(_01295_),
    .A1(_10422_),
    .A2(net208));
 sg13g2_buf_1 _17265_ (.A(net215),
    .X(_10424_));
 sg13g2_nand2_1 _17266_ (.Y(_10425_),
    .A(\top_ihp.oisc.regs[36][19] ),
    .B(net381));
 sg13g2_o21ai_1 _17267_ (.B1(_10425_),
    .Y(_01296_),
    .A1(net126),
    .A2(net208));
 sg13g2_buf_1 _17268_ (.A(net547),
    .X(_10426_));
 sg13g2_buf_2 _17269_ (.A(net383),
    .X(_10427_));
 sg13g2_nand2_1 _17270_ (.Y(_10428_),
    .A(\top_ihp.oisc.regs[36][1] ),
    .B(net381));
 sg13g2_o21ai_1 _17271_ (.B1(_10428_),
    .Y(_01297_),
    .A1(net380),
    .A2(net207));
 sg13g2_mux2_1 _17272_ (.A0(\top_ihp.oisc.regs[36][20] ),
    .A1(net137),
    .S(_10403_),
    .X(_01298_));
 sg13g2_buf_8 _17273_ (.A(net64),
    .X(_10429_));
 sg13g2_buf_2 _17274_ (.A(_10406_),
    .X(_10430_));
 sg13g2_nand2_1 _17275_ (.Y(_10431_),
    .A(\top_ihp.oisc.regs[36][21] ),
    .B(net379));
 sg13g2_o21ai_1 _17276_ (.B1(_10431_),
    .Y(_01299_),
    .A1(net38),
    .A2(net207));
 sg13g2_nand2_1 _17277_ (.Y(_10432_),
    .A(\top_ihp.oisc.regs[36][22] ),
    .B(_10430_));
 sg13g2_o21ai_1 _17278_ (.B1(_10432_),
    .Y(_01300_),
    .A1(net129),
    .A2(_10427_));
 sg13g2_mux2_1 _17279_ (.A0(\top_ihp.oisc.regs[36][23] ),
    .A1(net224),
    .S(_10403_),
    .X(_01301_));
 sg13g2_buf_1 _17280_ (.A(net214),
    .X(_10433_));
 sg13g2_nand2_1 _17281_ (.Y(_10434_),
    .A(\top_ihp.oisc.regs[36][24] ),
    .B(net379));
 sg13g2_o21ai_1 _17282_ (.B1(_10434_),
    .Y(_01302_),
    .A1(net125),
    .A2(net207));
 sg13g2_buf_2 _17283_ (.A(net213),
    .X(_10435_));
 sg13g2_nand2_1 _17284_ (.Y(_10436_),
    .A(\top_ihp.oisc.regs[36][25] ),
    .B(net379));
 sg13g2_o21ai_1 _17285_ (.B1(_10436_),
    .Y(_01303_),
    .A1(net124),
    .A2(net207));
 sg13g2_buf_8 _17286_ (.A(net134),
    .X(_10437_));
 sg13g2_nand2_1 _17287_ (.Y(_10438_),
    .A(\top_ihp.oisc.regs[36][26] ),
    .B(net379));
 sg13g2_o21ai_1 _17288_ (.B1(_10438_),
    .Y(_01304_),
    .A1(net55),
    .A2(net207));
 sg13g2_buf_8 _17289_ (.A(net141),
    .X(_10439_));
 sg13g2_nand2_1 _17290_ (.Y(_10440_),
    .A(\top_ihp.oisc.regs[36][27] ),
    .B(net379));
 sg13g2_o21ai_1 _17291_ (.B1(_10440_),
    .Y(_01305_),
    .A1(net54),
    .A2(_10427_));
 sg13g2_buf_8 _17292_ (.A(_10081_),
    .X(_10441_));
 sg13g2_nand2_1 _17293_ (.Y(_10442_),
    .A(\top_ihp.oisc.regs[36][28] ),
    .B(_10430_));
 sg13g2_o21ai_1 _17294_ (.B1(_10442_),
    .Y(_01306_),
    .A1(_10441_),
    .A2(net207));
 sg13g2_buf_2 _17295_ (.A(net133),
    .X(_10443_));
 sg13g2_nand2_1 _17296_ (.Y(_10444_),
    .A(\top_ihp.oisc.regs[36][29] ),
    .B(net379));
 sg13g2_o21ai_1 _17297_ (.B1(_10444_),
    .Y(_01307_),
    .A1(net53),
    .A2(net207));
 sg13g2_nand2_1 _17298_ (.Y(_10445_),
    .A(\top_ihp.oisc.regs[36][2] ),
    .B(net379));
 sg13g2_o21ai_1 _17299_ (.B1(_10445_),
    .Y(_01308_),
    .A1(net240),
    .A2(net207));
 sg13g2_nand2_1 _17300_ (.Y(_10446_),
    .A(\top_ihp.oisc.regs[36][30] ),
    .B(net379));
 sg13g2_o21ai_1 _17301_ (.B1(_10446_),
    .Y(_01309_),
    .A1(_09762_),
    .A2(_10409_));
 sg13g2_nand2_1 _17302_ (.Y(_10447_),
    .A(\top_ihp.oisc.regs[36][31] ),
    .B(_10407_));
 sg13g2_o21ai_1 _17303_ (.B1(_10447_),
    .Y(_01310_),
    .A1(_09782_),
    .A2(net382));
 sg13g2_nand2_1 _17304_ (.Y(_10448_),
    .A(\top_ihp.oisc.regs[36][3] ),
    .B(_10407_));
 sg13g2_o21ai_1 _17305_ (.B1(_10448_),
    .Y(_01311_),
    .A1(_09808_),
    .A2(_10409_));
 sg13g2_nand2_1 _17306_ (.Y(_10449_),
    .A(\top_ihp.oisc.regs[36][4] ),
    .B(net383));
 sg13g2_o21ai_1 _17307_ (.B1(_10449_),
    .Y(_01312_),
    .A1(_09841_),
    .A2(net382));
 sg13g2_buf_2 _17308_ (.A(net212),
    .X(_10450_));
 sg13g2_nand2_1 _17309_ (.Y(_10451_),
    .A(\top_ihp.oisc.regs[36][5] ),
    .B(net383));
 sg13g2_o21ai_1 _17310_ (.B1(_10451_),
    .Y(_01313_),
    .A1(net123),
    .A2(net382));
 sg13g2_buf_1 _17311_ (.A(net211),
    .X(_10452_));
 sg13g2_nand2_1 _17312_ (.Y(_10453_),
    .A(\top_ihp.oisc.regs[36][6] ),
    .B(net383));
 sg13g2_o21ai_1 _17313_ (.B1(_10453_),
    .Y(_01314_),
    .A1(net122),
    .A2(net382));
 sg13g2_nand2_1 _17314_ (.Y(_10454_),
    .A(\top_ihp.oisc.regs[36][7] ),
    .B(net383));
 sg13g2_o21ai_1 _17315_ (.B1(_10454_),
    .Y(_01315_),
    .A1(net209),
    .A2(net382));
 sg13g2_buf_1 _17316_ (.A(net61),
    .X(_10455_));
 sg13g2_nand2_1 _17317_ (.Y(_10456_),
    .A(\top_ihp.oisc.regs[36][8] ),
    .B(net383));
 sg13g2_o21ai_1 _17318_ (.B1(_10456_),
    .Y(_01316_),
    .A1(net36),
    .A2(net382));
 sg13g2_buf_8 _17319_ (.A(net60),
    .X(_10457_));
 sg13g2_nand2_1 _17320_ (.Y(_10458_),
    .A(\top_ihp.oisc.regs[36][9] ),
    .B(net383));
 sg13g2_o21ai_1 _17321_ (.B1(_10458_),
    .Y(_01317_),
    .A1(net35),
    .A2(net382));
 sg13g2_or3_1 _17322_ (.A(_09954_),
    .B(_09950_),
    .C(_09953_),
    .X(_10459_));
 sg13g2_buf_2 _17323_ (.A(_10459_),
    .X(_10460_));
 sg13g2_nor2_1 _17324_ (.A(_10276_),
    .B(net682),
    .Y(_10461_));
 sg13g2_buf_1 _17325_ (.A(_10461_),
    .X(_10462_));
 sg13g2_mux2_1 _17326_ (.A0(\top_ihp.oisc.regs[37][0] ),
    .A1(_10107_),
    .S(_10462_),
    .X(_01318_));
 sg13g2_nand2b_1 _17327_ (.Y(_10463_),
    .B(net663),
    .A_N(_10276_));
 sg13g2_buf_2 _17328_ (.A(_10463_),
    .X(_10464_));
 sg13g2_buf_1 _17329_ (.A(_10464_),
    .X(_10465_));
 sg13g2_buf_1 _17330_ (.A(_10464_),
    .X(_10466_));
 sg13g2_nand2_1 _17331_ (.Y(_10467_),
    .A(\top_ihp.oisc.regs[37][10] ),
    .B(net377));
 sg13g2_o21ai_1 _17332_ (.B1(_10467_),
    .Y(_01319_),
    .A1(_10404_),
    .A2(net378));
 sg13g2_buf_1 _17333_ (.A(net251),
    .X(_10468_));
 sg13g2_nand2_1 _17334_ (.Y(_10469_),
    .A(\top_ihp.oisc.regs[37][11] ),
    .B(net377));
 sg13g2_o21ai_1 _17335_ (.B1(_10469_),
    .Y(_01320_),
    .A1(net121),
    .A2(net378));
 sg13g2_nand2_1 _17336_ (.Y(_10470_),
    .A(\top_ihp.oisc.regs[37][12] ),
    .B(net377));
 sg13g2_o21ai_1 _17337_ (.B1(_10470_),
    .Y(_01321_),
    .A1(net128),
    .A2(net378));
 sg13g2_nor2_1 _17338_ (.A(\top_ihp.oisc.regs[37][13] ),
    .B(net524),
    .Y(_10471_));
 sg13g2_a21oi_1 _17339_ (.A1(net59),
    .A2(net524),
    .Y(_01322_),
    .B1(_10471_));
 sg13g2_nand2_1 _17340_ (.Y(_10472_),
    .A(\top_ihp.oisc.regs[37][14] ),
    .B(net377));
 sg13g2_o21ai_1 _17341_ (.B1(_10472_),
    .Y(_01323_),
    .A1(net127),
    .A2(net378));
 sg13g2_buf_1 _17342_ (.A(net216),
    .X(_10473_));
 sg13g2_buf_2 _17343_ (.A(_10464_),
    .X(_10474_));
 sg13g2_nand2_1 _17344_ (.Y(_10475_),
    .A(\top_ihp.oisc.regs[37][15] ),
    .B(net376));
 sg13g2_o21ai_1 _17345_ (.B1(_10475_),
    .Y(_01324_),
    .A1(net120),
    .A2(net378));
 sg13g2_nor2_1 _17346_ (.A(\top_ihp.oisc.regs[37][16] ),
    .B(net524),
    .Y(_10476_));
 sg13g2_a21oi_1 _17347_ (.A1(net132),
    .A2(net524),
    .Y(_01325_),
    .B1(_10476_));
 sg13g2_nand2_1 _17348_ (.Y(_10477_),
    .A(\top_ihp.oisc.regs[37][17] ),
    .B(net376));
 sg13g2_o21ai_1 _17349_ (.B1(_10477_),
    .Y(_01326_),
    .A1(net57),
    .A2(net378));
 sg13g2_nand2_1 _17350_ (.Y(_10478_),
    .A(\top_ihp.oisc.regs[37][18] ),
    .B(net376));
 sg13g2_o21ai_1 _17351_ (.B1(_10478_),
    .Y(_01327_),
    .A1(net56),
    .A2(_10465_));
 sg13g2_nand2_1 _17352_ (.Y(_10479_),
    .A(\top_ihp.oisc.regs[37][19] ),
    .B(net376));
 sg13g2_o21ai_1 _17353_ (.B1(_10479_),
    .Y(_01328_),
    .A1(net126),
    .A2(net378));
 sg13g2_nand2_1 _17354_ (.Y(_10480_),
    .A(\top_ihp.oisc.regs[37][1] ),
    .B(net376));
 sg13g2_o21ai_1 _17355_ (.B1(_10480_),
    .Y(_01329_),
    .A1(_10426_),
    .A2(_10465_));
 sg13g2_nor2_1 _17356_ (.A(\top_ihp.oisc.regs[37][20] ),
    .B(net524),
    .Y(_10481_));
 sg13g2_a21oi_1 _17357_ (.A1(net40),
    .A2(net524),
    .Y(_01330_),
    .B1(_10481_));
 sg13g2_nand2_1 _17358_ (.Y(_10482_),
    .A(\top_ihp.oisc.regs[37][21] ),
    .B(net376));
 sg13g2_o21ai_1 _17359_ (.B1(_10482_),
    .Y(_01331_),
    .A1(_10429_),
    .A2(net378));
 sg13g2_nor2_1 _17360_ (.A(\top_ihp.oisc.regs[37][22] ),
    .B(net524),
    .Y(_10483_));
 sg13g2_a21oi_1 _17361_ (.A1(net131),
    .A2(_10462_),
    .Y(_01332_),
    .B1(_10483_));
 sg13g2_nor2_1 _17362_ (.A(\top_ihp.oisc.regs[37][23] ),
    .B(_10461_),
    .Y(_10484_));
 sg13g2_a21oi_1 _17363_ (.A1(net138),
    .A2(net524),
    .Y(_01333_),
    .B1(_10484_));
 sg13g2_buf_1 _17364_ (.A(_10464_),
    .X(_10485_));
 sg13g2_nand2_1 _17365_ (.Y(_10486_),
    .A(\top_ihp.oisc.regs[37][24] ),
    .B(net376));
 sg13g2_o21ai_1 _17366_ (.B1(_10486_),
    .Y(_01334_),
    .A1(net125),
    .A2(net375));
 sg13g2_nand2_1 _17367_ (.Y(_10487_),
    .A(\top_ihp.oisc.regs[37][25] ),
    .B(net376));
 sg13g2_o21ai_1 _17368_ (.B1(_10487_),
    .Y(_01335_),
    .A1(net124),
    .A2(net375));
 sg13g2_nand2_1 _17369_ (.Y(_10488_),
    .A(\top_ihp.oisc.regs[37][26] ),
    .B(_10474_));
 sg13g2_o21ai_1 _17370_ (.B1(_10488_),
    .Y(_01336_),
    .A1(net55),
    .A2(net375));
 sg13g2_nand2_1 _17371_ (.Y(_10489_),
    .A(\top_ihp.oisc.regs[37][27] ),
    .B(_10474_));
 sg13g2_o21ai_1 _17372_ (.B1(_10489_),
    .Y(_01337_),
    .A1(net54),
    .A2(_10485_));
 sg13g2_buf_1 _17373_ (.A(_10464_),
    .X(_10490_));
 sg13g2_nand2_1 _17374_ (.Y(_10491_),
    .A(\top_ihp.oisc.regs[37][28] ),
    .B(net374));
 sg13g2_o21ai_1 _17375_ (.B1(_10491_),
    .Y(_01338_),
    .A1(net37),
    .A2(_10485_));
 sg13g2_nand2_1 _17376_ (.Y(_10492_),
    .A(\top_ihp.oisc.regs[37][29] ),
    .B(net374));
 sg13g2_o21ai_1 _17377_ (.B1(_10492_),
    .Y(_01339_),
    .A1(net53),
    .A2(net375));
 sg13g2_buf_2 _17378_ (.A(net222),
    .X(_10493_));
 sg13g2_nand2_1 _17379_ (.Y(_10494_),
    .A(\top_ihp.oisc.regs[37][2] ),
    .B(_10490_));
 sg13g2_o21ai_1 _17380_ (.B1(_10494_),
    .Y(_01340_),
    .A1(net119),
    .A2(net375));
 sg13g2_buf_1 _17381_ (.A(net62),
    .X(_10495_));
 sg13g2_nand2_1 _17382_ (.Y(_10496_),
    .A(\top_ihp.oisc.regs[37][30] ),
    .B(_10490_));
 sg13g2_o21ai_1 _17383_ (.B1(_10496_),
    .Y(_01341_),
    .A1(net34),
    .A2(net375));
 sg13g2_nand2_1 _17384_ (.Y(_10497_),
    .A(\top_ihp.oisc.regs[37][31] ),
    .B(net374));
 sg13g2_o21ai_1 _17385_ (.B1(_10497_),
    .Y(_01342_),
    .A1(_09782_),
    .A2(net375));
 sg13g2_buf_1 _17386_ (.A(net221),
    .X(_10498_));
 sg13g2_nand2_1 _17387_ (.Y(_10499_),
    .A(\top_ihp.oisc.regs[37][3] ),
    .B(net374));
 sg13g2_o21ai_1 _17388_ (.B1(_10499_),
    .Y(_01343_),
    .A1(net118),
    .A2(net375));
 sg13g2_buf_2 _17389_ (.A(net220),
    .X(_10500_));
 sg13g2_nand2_1 _17390_ (.Y(_10501_),
    .A(\top_ihp.oisc.regs[37][4] ),
    .B(net374));
 sg13g2_o21ai_1 _17391_ (.B1(_10501_),
    .Y(_01344_),
    .A1(net117),
    .A2(net377));
 sg13g2_nand2_1 _17392_ (.Y(_10502_),
    .A(\top_ihp.oisc.regs[37][5] ),
    .B(net374));
 sg13g2_o21ai_1 _17393_ (.B1(_10502_),
    .Y(_01345_),
    .A1(net123),
    .A2(net377));
 sg13g2_nand2_1 _17394_ (.Y(_10503_),
    .A(\top_ihp.oisc.regs[37][6] ),
    .B(net374));
 sg13g2_o21ai_1 _17395_ (.B1(_10503_),
    .Y(_01346_),
    .A1(net122),
    .A2(_10466_));
 sg13g2_nand2_1 _17396_ (.Y(_10504_),
    .A(\top_ihp.oisc.regs[37][7] ),
    .B(net374));
 sg13g2_o21ai_1 _17397_ (.B1(_10504_),
    .Y(_01347_),
    .A1(net209),
    .A2(net377));
 sg13g2_nand2_1 _17398_ (.Y(_10505_),
    .A(\top_ihp.oisc.regs[37][8] ),
    .B(_10464_));
 sg13g2_o21ai_1 _17399_ (.B1(_10505_),
    .Y(_01348_),
    .A1(net36),
    .A2(net377));
 sg13g2_nand2_1 _17400_ (.Y(_10506_),
    .A(\top_ihp.oisc.regs[37][9] ),
    .B(_10464_));
 sg13g2_o21ai_1 _17401_ (.B1(_10506_),
    .Y(_01349_),
    .A1(net35),
    .A2(_10466_));
 sg13g2_and2_1 _17402_ (.A(net664),
    .B(net663),
    .X(_10507_));
 sg13g2_buf_1 _17403_ (.A(_10507_),
    .X(_10508_));
 sg13g2_mux2_1 _17404_ (.A0(\top_ihp.oisc.regs[38][0] ),
    .A1(_10107_),
    .S(_10508_),
    .X(_01350_));
 sg13g2_nand2_1 _17405_ (.Y(_10509_),
    .A(net664),
    .B(net663));
 sg13g2_buf_1 _17406_ (.A(_10509_),
    .X(_10510_));
 sg13g2_buf_1 _17407_ (.A(_10510_),
    .X(_10511_));
 sg13g2_buf_1 _17408_ (.A(net373),
    .X(_10512_));
 sg13g2_buf_1 _17409_ (.A(_10510_),
    .X(_10513_));
 sg13g2_nand2_1 _17410_ (.Y(_10514_),
    .A(\top_ihp.oisc.regs[38][10] ),
    .B(net372));
 sg13g2_o21ai_1 _17411_ (.B1(_10514_),
    .Y(_01351_),
    .A1(net39),
    .A2(net206));
 sg13g2_buf_1 _17412_ (.A(_10510_),
    .X(_10515_));
 sg13g2_nand2_1 _17413_ (.Y(_10516_),
    .A(\top_ihp.oisc.regs[38][11] ),
    .B(net371));
 sg13g2_o21ai_1 _17414_ (.B1(_10516_),
    .Y(_01352_),
    .A1(net121),
    .A2(_10512_));
 sg13g2_nand2_1 _17415_ (.Y(_10517_),
    .A(\top_ihp.oisc.regs[38][12] ),
    .B(net371));
 sg13g2_o21ai_1 _17416_ (.B1(_10517_),
    .Y(_01353_),
    .A1(net128),
    .A2(_10512_));
 sg13g2_nand2_1 _17417_ (.Y(_10518_),
    .A(\top_ihp.oisc.regs[38][13] ),
    .B(_10515_));
 sg13g2_o21ai_1 _17418_ (.B1(_10518_),
    .Y(_01354_),
    .A1(net58),
    .A2(net206));
 sg13g2_nand2_1 _17419_ (.Y(_10519_),
    .A(\top_ihp.oisc.regs[38][14] ),
    .B(net371));
 sg13g2_o21ai_1 _17420_ (.B1(_10519_),
    .Y(_01355_),
    .A1(net127),
    .A2(net206));
 sg13g2_nand2_1 _17421_ (.Y(_10520_),
    .A(\top_ihp.oisc.regs[38][15] ),
    .B(net371));
 sg13g2_o21ai_1 _17422_ (.B1(_10520_),
    .Y(_01356_),
    .A1(net120),
    .A2(net206));
 sg13g2_nand2_1 _17423_ (.Y(_10521_),
    .A(\top_ihp.oisc.regs[38][16] ),
    .B(_10515_));
 sg13g2_o21ai_1 _17424_ (.B1(_10521_),
    .Y(_01357_),
    .A1(net130),
    .A2(net206));
 sg13g2_nand2_1 _17425_ (.Y(_10522_),
    .A(\top_ihp.oisc.regs[38][17] ),
    .B(net371));
 sg13g2_o21ai_1 _17426_ (.B1(_10522_),
    .Y(_01358_),
    .A1(_10420_),
    .A2(net206));
 sg13g2_nand2_1 _17427_ (.Y(_10523_),
    .A(\top_ihp.oisc.regs[38][18] ),
    .B(net371));
 sg13g2_o21ai_1 _17428_ (.B1(_10523_),
    .Y(_01359_),
    .A1(net56),
    .A2(net206));
 sg13g2_nand2_1 _17429_ (.Y(_10524_),
    .A(\top_ihp.oisc.regs[38][19] ),
    .B(net371));
 sg13g2_o21ai_1 _17430_ (.B1(_10524_),
    .Y(_01360_),
    .A1(net126),
    .A2(net206));
 sg13g2_buf_1 _17431_ (.A(_10511_),
    .X(_10525_));
 sg13g2_nand2_1 _17432_ (.Y(_10526_),
    .A(\top_ihp.oisc.regs[38][1] ),
    .B(net371));
 sg13g2_o21ai_1 _17433_ (.B1(_10526_),
    .Y(_01361_),
    .A1(net380),
    .A2(net205));
 sg13g2_nor2_1 _17434_ (.A(\top_ihp.oisc.regs[38][20] ),
    .B(_10508_),
    .Y(_10527_));
 sg13g2_a21oi_1 _17435_ (.A1(net40),
    .A2(_10508_),
    .Y(_01362_),
    .B1(_10527_));
 sg13g2_buf_1 _17436_ (.A(_10510_),
    .X(_10528_));
 sg13g2_nand2_1 _17437_ (.Y(_10529_),
    .A(\top_ihp.oisc.regs[38][21] ),
    .B(net370));
 sg13g2_o21ai_1 _17438_ (.B1(_10529_),
    .Y(_01363_),
    .A1(net38),
    .A2(net205));
 sg13g2_nand2_1 _17439_ (.Y(_10530_),
    .A(\top_ihp.oisc.regs[38][22] ),
    .B(net370));
 sg13g2_o21ai_1 _17440_ (.B1(_10530_),
    .Y(_01364_),
    .A1(net129),
    .A2(net205));
 sg13g2_nor2_1 _17441_ (.A(\top_ihp.oisc.regs[38][23] ),
    .B(_10508_),
    .Y(_10531_));
 sg13g2_a21oi_1 _17442_ (.A1(net138),
    .A2(_10508_),
    .Y(_01365_),
    .B1(_10531_));
 sg13g2_nand2_1 _17443_ (.Y(_10532_),
    .A(\top_ihp.oisc.regs[38][24] ),
    .B(_10528_));
 sg13g2_o21ai_1 _17444_ (.B1(_10532_),
    .Y(_01366_),
    .A1(_10433_),
    .A2(_10525_));
 sg13g2_nand2_1 _17445_ (.Y(_10533_),
    .A(\top_ihp.oisc.regs[38][25] ),
    .B(net370));
 sg13g2_o21ai_1 _17446_ (.B1(_10533_),
    .Y(_01367_),
    .A1(net124),
    .A2(net205));
 sg13g2_nand2_1 _17447_ (.Y(_10534_),
    .A(\top_ihp.oisc.regs[38][26] ),
    .B(net370));
 sg13g2_o21ai_1 _17448_ (.B1(_10534_),
    .Y(_01368_),
    .A1(net55),
    .A2(net205));
 sg13g2_nand2_1 _17449_ (.Y(_10535_),
    .A(\top_ihp.oisc.regs[38][27] ),
    .B(net370));
 sg13g2_o21ai_1 _17450_ (.B1(_10535_),
    .Y(_01369_),
    .A1(net54),
    .A2(net205));
 sg13g2_nand2_1 _17451_ (.Y(_10536_),
    .A(\top_ihp.oisc.regs[38][28] ),
    .B(net370));
 sg13g2_o21ai_1 _17452_ (.B1(_10536_),
    .Y(_01370_),
    .A1(net37),
    .A2(_10525_));
 sg13g2_nand2_1 _17453_ (.Y(_10537_),
    .A(\top_ihp.oisc.regs[38][29] ),
    .B(net370));
 sg13g2_o21ai_1 _17454_ (.B1(_10537_),
    .Y(_01371_),
    .A1(net53),
    .A2(net205));
 sg13g2_nand2_1 _17455_ (.Y(_10538_),
    .A(\top_ihp.oisc.regs[38][2] ),
    .B(net370));
 sg13g2_o21ai_1 _17456_ (.B1(_10538_),
    .Y(_01372_),
    .A1(net119),
    .A2(net205));
 sg13g2_nand2_1 _17457_ (.Y(_10539_),
    .A(\top_ihp.oisc.regs[38][30] ),
    .B(_10528_));
 sg13g2_o21ai_1 _17458_ (.B1(_10539_),
    .Y(_01373_),
    .A1(net34),
    .A2(net372));
 sg13g2_buf_8 _17459_ (.A(net239),
    .X(_10540_));
 sg13g2_nand2_1 _17460_ (.Y(_10541_),
    .A(\top_ihp.oisc.regs[38][31] ),
    .B(net373));
 sg13g2_o21ai_1 _17461_ (.B1(_10541_),
    .Y(_01374_),
    .A1(net116),
    .A2(_10513_));
 sg13g2_nand2_1 _17462_ (.Y(_10542_),
    .A(\top_ihp.oisc.regs[38][3] ),
    .B(net373));
 sg13g2_o21ai_1 _17463_ (.B1(_10542_),
    .Y(_01375_),
    .A1(net118),
    .A2(net372));
 sg13g2_nand2_1 _17464_ (.Y(_10543_),
    .A(\top_ihp.oisc.regs[38][4] ),
    .B(_10511_));
 sg13g2_o21ai_1 _17465_ (.B1(_10543_),
    .Y(_01376_),
    .A1(_10500_),
    .A2(_10513_));
 sg13g2_nand2_1 _17466_ (.Y(_10544_),
    .A(\top_ihp.oisc.regs[38][5] ),
    .B(net373));
 sg13g2_o21ai_1 _17467_ (.B1(_10544_),
    .Y(_01377_),
    .A1(net123),
    .A2(net372));
 sg13g2_nand2_1 _17468_ (.Y(_10545_),
    .A(\top_ihp.oisc.regs[38][6] ),
    .B(net373));
 sg13g2_o21ai_1 _17469_ (.B1(_10545_),
    .Y(_01378_),
    .A1(net122),
    .A2(net372));
 sg13g2_nand2_1 _17470_ (.Y(_10546_),
    .A(\top_ihp.oisc.regs[38][7] ),
    .B(net373));
 sg13g2_o21ai_1 _17471_ (.B1(_10546_),
    .Y(_01379_),
    .A1(net68),
    .A2(net372));
 sg13g2_nand2_1 _17472_ (.Y(_10547_),
    .A(\top_ihp.oisc.regs[38][8] ),
    .B(net373));
 sg13g2_o21ai_1 _17473_ (.B1(_10547_),
    .Y(_01380_),
    .A1(net36),
    .A2(net372));
 sg13g2_nand2_1 _17474_ (.Y(_10548_),
    .A(\top_ihp.oisc.regs[38][9] ),
    .B(net373));
 sg13g2_o21ai_1 _17475_ (.B1(_10548_),
    .Y(_01381_),
    .A1(net35),
    .A2(net372));
 sg13g2_buf_2 _17476_ (.A(net412),
    .X(_10549_));
 sg13g2_and2_1 _17477_ (.A(_10358_),
    .B(_10398_),
    .X(_10550_));
 sg13g2_buf_1 _17478_ (.A(_10550_),
    .X(_10551_));
 sg13g2_mux2_1 _17479_ (.A0(\top_ihp.oisc.regs[39][0] ),
    .A1(net204),
    .S(_10551_),
    .X(_01382_));
 sg13g2_nand2_1 _17480_ (.Y(_10552_),
    .A(_10358_),
    .B(_10397_));
 sg13g2_buf_1 _17481_ (.A(_10552_),
    .X(_10553_));
 sg13g2_buf_1 _17482_ (.A(_10553_),
    .X(_10554_));
 sg13g2_buf_1 _17483_ (.A(net369),
    .X(_10555_));
 sg13g2_buf_1 _17484_ (.A(_10553_),
    .X(_10556_));
 sg13g2_nand2_1 _17485_ (.Y(_10557_),
    .A(\top_ihp.oisc.regs[39][10] ),
    .B(net368));
 sg13g2_o21ai_1 _17486_ (.B1(_10557_),
    .Y(_01383_),
    .A1(net39),
    .A2(net203));
 sg13g2_buf_1 _17487_ (.A(_10553_),
    .X(_10558_));
 sg13g2_nand2_1 _17488_ (.Y(_10559_),
    .A(\top_ihp.oisc.regs[39][11] ),
    .B(net367));
 sg13g2_o21ai_1 _17489_ (.B1(_10559_),
    .Y(_01384_),
    .A1(_10468_),
    .A2(_10555_));
 sg13g2_nand2_1 _17490_ (.Y(_10560_),
    .A(\top_ihp.oisc.regs[39][12] ),
    .B(net367));
 sg13g2_o21ai_1 _17491_ (.B1(_10560_),
    .Y(_01385_),
    .A1(net128),
    .A2(net203));
 sg13g2_nand2_1 _17492_ (.Y(_10561_),
    .A(\top_ihp.oisc.regs[39][13] ),
    .B(_10558_));
 sg13g2_o21ai_1 _17493_ (.B1(_10561_),
    .Y(_01386_),
    .A1(net58),
    .A2(net203));
 sg13g2_nand2_1 _17494_ (.Y(_10562_),
    .A(\top_ihp.oisc.regs[39][14] ),
    .B(net367));
 sg13g2_o21ai_1 _17495_ (.B1(_10562_),
    .Y(_01387_),
    .A1(_10416_),
    .A2(_10555_));
 sg13g2_nand2_1 _17496_ (.Y(_10563_),
    .A(\top_ihp.oisc.regs[39][15] ),
    .B(net367));
 sg13g2_o21ai_1 _17497_ (.B1(_10563_),
    .Y(_01388_),
    .A1(net120),
    .A2(net203));
 sg13g2_nand2_1 _17498_ (.Y(_10564_),
    .A(\top_ihp.oisc.regs[39][16] ),
    .B(net367));
 sg13g2_o21ai_1 _17499_ (.B1(_10564_),
    .Y(_01389_),
    .A1(net130),
    .A2(net203));
 sg13g2_nand2_1 _17500_ (.Y(_10565_),
    .A(\top_ihp.oisc.regs[39][17] ),
    .B(net367));
 sg13g2_o21ai_1 _17501_ (.B1(_10565_),
    .Y(_01390_),
    .A1(net57),
    .A2(net203));
 sg13g2_nand2_1 _17502_ (.Y(_10566_),
    .A(\top_ihp.oisc.regs[39][18] ),
    .B(_10558_));
 sg13g2_o21ai_1 _17503_ (.B1(_10566_),
    .Y(_01391_),
    .A1(net56),
    .A2(net203));
 sg13g2_nand2_1 _17504_ (.Y(_10567_),
    .A(\top_ihp.oisc.regs[39][19] ),
    .B(net367));
 sg13g2_o21ai_1 _17505_ (.B1(_10567_),
    .Y(_01392_),
    .A1(net126),
    .A2(net203));
 sg13g2_buf_1 _17506_ (.A(_10554_),
    .X(_10568_));
 sg13g2_nand2_1 _17507_ (.Y(_10569_),
    .A(\top_ihp.oisc.regs[39][1] ),
    .B(net367));
 sg13g2_o21ai_1 _17508_ (.B1(_10569_),
    .Y(_01393_),
    .A1(net380),
    .A2(net202));
 sg13g2_mux2_1 _17509_ (.A0(\top_ihp.oisc.regs[39][20] ),
    .A1(net137),
    .S(_10551_),
    .X(_01394_));
 sg13g2_buf_1 _17510_ (.A(_10553_),
    .X(_10570_));
 sg13g2_nand2_1 _17511_ (.Y(_10571_),
    .A(\top_ihp.oisc.regs[39][21] ),
    .B(net366));
 sg13g2_o21ai_1 _17512_ (.B1(_10571_),
    .Y(_01395_),
    .A1(net38),
    .A2(net202));
 sg13g2_nand2_1 _17513_ (.Y(_10572_),
    .A(\top_ihp.oisc.regs[39][22] ),
    .B(net366));
 sg13g2_o21ai_1 _17514_ (.B1(_10572_),
    .Y(_01396_),
    .A1(net129),
    .A2(net202));
 sg13g2_mux2_1 _17515_ (.A0(\top_ihp.oisc.regs[39][23] ),
    .A1(_10036_),
    .S(_10551_),
    .X(_01397_));
 sg13g2_nand2_1 _17516_ (.Y(_10573_),
    .A(\top_ihp.oisc.regs[39][24] ),
    .B(_10570_));
 sg13g2_o21ai_1 _17517_ (.B1(_10573_),
    .Y(_01398_),
    .A1(net125),
    .A2(_10568_));
 sg13g2_nand2_1 _17518_ (.Y(_10574_),
    .A(\top_ihp.oisc.regs[39][25] ),
    .B(net366));
 sg13g2_o21ai_1 _17519_ (.B1(_10574_),
    .Y(_01399_),
    .A1(net124),
    .A2(net202));
 sg13g2_nand2_1 _17520_ (.Y(_10575_),
    .A(\top_ihp.oisc.regs[39][26] ),
    .B(net366));
 sg13g2_o21ai_1 _17521_ (.B1(_10575_),
    .Y(_01400_),
    .A1(net55),
    .A2(net202));
 sg13g2_nand2_1 _17522_ (.Y(_10576_),
    .A(\top_ihp.oisc.regs[39][27] ),
    .B(_10570_));
 sg13g2_o21ai_1 _17523_ (.B1(_10576_),
    .Y(_01401_),
    .A1(net54),
    .A2(_10568_));
 sg13g2_nand2_1 _17524_ (.Y(_10577_),
    .A(\top_ihp.oisc.regs[39][28] ),
    .B(net366));
 sg13g2_o21ai_1 _17525_ (.B1(_10577_),
    .Y(_01402_),
    .A1(net37),
    .A2(net202));
 sg13g2_nand2_1 _17526_ (.Y(_10578_),
    .A(\top_ihp.oisc.regs[39][29] ),
    .B(net366));
 sg13g2_o21ai_1 _17527_ (.B1(_10578_),
    .Y(_01403_),
    .A1(net53),
    .A2(net202));
 sg13g2_nand2_1 _17528_ (.Y(_10579_),
    .A(\top_ihp.oisc.regs[39][2] ),
    .B(net366));
 sg13g2_o21ai_1 _17529_ (.B1(_10579_),
    .Y(_01404_),
    .A1(net119),
    .A2(net202));
 sg13g2_nand2_1 _17530_ (.Y(_10580_),
    .A(\top_ihp.oisc.regs[39][30] ),
    .B(net366));
 sg13g2_o21ai_1 _17531_ (.B1(_10580_),
    .Y(_01405_),
    .A1(net34),
    .A2(_10556_));
 sg13g2_nand2_1 _17532_ (.Y(_10581_),
    .A(\top_ihp.oisc.regs[39][31] ),
    .B(net369));
 sg13g2_o21ai_1 _17533_ (.B1(_10581_),
    .Y(_01406_),
    .A1(net116),
    .A2(net368));
 sg13g2_nand2_1 _17534_ (.Y(_10582_),
    .A(\top_ihp.oisc.regs[39][3] ),
    .B(net369));
 sg13g2_o21ai_1 _17535_ (.B1(_10582_),
    .Y(_01407_),
    .A1(net118),
    .A2(net368));
 sg13g2_nand2_1 _17536_ (.Y(_10583_),
    .A(\top_ihp.oisc.regs[39][4] ),
    .B(_10554_));
 sg13g2_o21ai_1 _17537_ (.B1(_10583_),
    .Y(_01408_),
    .A1(net117),
    .A2(_10556_));
 sg13g2_nand2_1 _17538_ (.Y(_10584_),
    .A(\top_ihp.oisc.regs[39][5] ),
    .B(net369));
 sg13g2_o21ai_1 _17539_ (.B1(_10584_),
    .Y(_01409_),
    .A1(net123),
    .A2(net368));
 sg13g2_nand2_1 _17540_ (.Y(_10585_),
    .A(\top_ihp.oisc.regs[39][6] ),
    .B(net369));
 sg13g2_o21ai_1 _17541_ (.B1(_10585_),
    .Y(_01410_),
    .A1(net122),
    .A2(net368));
 sg13g2_nand2_1 _17542_ (.Y(_10586_),
    .A(\top_ihp.oisc.regs[39][7] ),
    .B(net369));
 sg13g2_o21ai_1 _17543_ (.B1(_10586_),
    .Y(_01411_),
    .A1(net209),
    .A2(net368));
 sg13g2_nand2_1 _17544_ (.Y(_10587_),
    .A(\top_ihp.oisc.regs[39][8] ),
    .B(net369));
 sg13g2_o21ai_1 _17545_ (.B1(_10587_),
    .Y(_01412_),
    .A1(net36),
    .A2(net368));
 sg13g2_nand2_1 _17546_ (.Y(_10588_),
    .A(\top_ihp.oisc.regs[39][9] ),
    .B(net369));
 sg13g2_o21ai_1 _17547_ (.B1(_10588_),
    .Y(_01413_),
    .A1(_10457_),
    .A2(net368));
 sg13g2_and2_1 _17548_ (.A(_09106_),
    .B(_10009_),
    .X(_10589_));
 sg13g2_buf_1 _17549_ (.A(_10589_),
    .X(_10590_));
 sg13g2_mux2_1 _17550_ (.A0(\top_ihp.oisc.regs[3][0] ),
    .A1(_10549_),
    .S(_10590_),
    .X(_01414_));
 sg13g2_nand2_1 _17551_ (.Y(_10591_),
    .A(_09106_),
    .B(_10009_));
 sg13g2_buf_1 _17552_ (.A(_10591_),
    .X(_10592_));
 sg13g2_buf_1 _17553_ (.A(_10592_),
    .X(_10593_));
 sg13g2_buf_1 _17554_ (.A(net523),
    .X(_10594_));
 sg13g2_buf_1 _17555_ (.A(_10592_),
    .X(_10595_));
 sg13g2_nand2_1 _17556_ (.Y(_10596_),
    .A(\top_ihp.oisc.regs[3][10] ),
    .B(net522));
 sg13g2_o21ai_1 _17557_ (.B1(_10596_),
    .Y(_01415_),
    .A1(_10404_),
    .A2(net365));
 sg13g2_buf_1 _17558_ (.A(_10592_),
    .X(_10597_));
 sg13g2_nand2_1 _17559_ (.Y(_10598_),
    .A(\top_ihp.oisc.regs[3][11] ),
    .B(net521));
 sg13g2_o21ai_1 _17560_ (.B1(_10598_),
    .Y(_01416_),
    .A1(_10468_),
    .A2(net365));
 sg13g2_nand2_1 _17561_ (.Y(_10599_),
    .A(\top_ihp.oisc.regs[3][12] ),
    .B(net521));
 sg13g2_o21ai_1 _17562_ (.B1(_10599_),
    .Y(_01417_),
    .A1(net128),
    .A2(net365));
 sg13g2_nand2_1 _17563_ (.Y(_10600_),
    .A(\top_ihp.oisc.regs[3][13] ),
    .B(net521));
 sg13g2_o21ai_1 _17564_ (.B1(_10600_),
    .Y(_01418_),
    .A1(net58),
    .A2(net365));
 sg13g2_nand2_1 _17565_ (.Y(_10601_),
    .A(\top_ihp.oisc.regs[3][14] ),
    .B(net521));
 sg13g2_o21ai_1 _17566_ (.B1(_10601_),
    .Y(_01419_),
    .A1(net127),
    .A2(net365));
 sg13g2_nand2_1 _17567_ (.Y(_10602_),
    .A(\top_ihp.oisc.regs[3][15] ),
    .B(net521));
 sg13g2_o21ai_1 _17568_ (.B1(_10602_),
    .Y(_01420_),
    .A1(net120),
    .A2(net365));
 sg13g2_nand2_1 _17569_ (.Y(_10603_),
    .A(\top_ihp.oisc.regs[3][16] ),
    .B(net521));
 sg13g2_o21ai_1 _17570_ (.B1(_10603_),
    .Y(_01421_),
    .A1(_10163_),
    .A2(net365));
 sg13g2_nand2_1 _17571_ (.Y(_10604_),
    .A(\top_ihp.oisc.regs[3][17] ),
    .B(net521));
 sg13g2_o21ai_1 _17572_ (.B1(_10604_),
    .Y(_01422_),
    .A1(_10420_),
    .A2(net365));
 sg13g2_nand2_1 _17573_ (.Y(_10605_),
    .A(\top_ihp.oisc.regs[3][18] ),
    .B(_10597_));
 sg13g2_o21ai_1 _17574_ (.B1(_10605_),
    .Y(_01423_),
    .A1(_10422_),
    .A2(_10594_));
 sg13g2_nand2_1 _17575_ (.Y(_10606_),
    .A(\top_ihp.oisc.regs[3][19] ),
    .B(_10597_));
 sg13g2_o21ai_1 _17576_ (.B1(_10606_),
    .Y(_01424_),
    .A1(net126),
    .A2(_10594_));
 sg13g2_buf_1 _17577_ (.A(_10593_),
    .X(_10607_));
 sg13g2_nand2_1 _17578_ (.Y(_10608_),
    .A(\top_ihp.oisc.regs[3][1] ),
    .B(net521));
 sg13g2_o21ai_1 _17579_ (.B1(_10608_),
    .Y(_01425_),
    .A1(net380),
    .A2(net364));
 sg13g2_mux2_1 _17580_ (.A0(\top_ihp.oisc.regs[3][20] ),
    .A1(net137),
    .S(_10590_),
    .X(_01426_));
 sg13g2_buf_1 _17581_ (.A(_10592_),
    .X(_10609_));
 sg13g2_nand2_1 _17582_ (.Y(_10610_),
    .A(\top_ihp.oisc.regs[3][21] ),
    .B(net520));
 sg13g2_o21ai_1 _17583_ (.B1(_10610_),
    .Y(_01427_),
    .A1(net38),
    .A2(net364));
 sg13g2_nand2_1 _17584_ (.Y(_10611_),
    .A(\top_ihp.oisc.regs[3][22] ),
    .B(net520));
 sg13g2_o21ai_1 _17585_ (.B1(_10611_),
    .Y(_01428_),
    .A1(net129),
    .A2(net364));
 sg13g2_mux2_1 _17586_ (.A0(\top_ihp.oisc.regs[3][23] ),
    .A1(net224),
    .S(_10590_),
    .X(_01429_));
 sg13g2_nand2_1 _17587_ (.Y(_10612_),
    .A(\top_ihp.oisc.regs[3][24] ),
    .B(net520));
 sg13g2_o21ai_1 _17588_ (.B1(_10612_),
    .Y(_01430_),
    .A1(_10433_),
    .A2(_10607_));
 sg13g2_nand2_1 _17589_ (.Y(_10613_),
    .A(\top_ihp.oisc.regs[3][25] ),
    .B(_10609_));
 sg13g2_o21ai_1 _17590_ (.B1(_10613_),
    .Y(_01431_),
    .A1(net124),
    .A2(_10607_));
 sg13g2_nand2_1 _17591_ (.Y(_10614_),
    .A(\top_ihp.oisc.regs[3][26] ),
    .B(net520));
 sg13g2_o21ai_1 _17592_ (.B1(_10614_),
    .Y(_01432_),
    .A1(net55),
    .A2(net364));
 sg13g2_nand2_1 _17593_ (.Y(_10615_),
    .A(\top_ihp.oisc.regs[3][27] ),
    .B(net520));
 sg13g2_o21ai_1 _17594_ (.B1(_10615_),
    .Y(_01433_),
    .A1(_10439_),
    .A2(net364));
 sg13g2_nand2_1 _17595_ (.Y(_10616_),
    .A(\top_ihp.oisc.regs[3][28] ),
    .B(net520));
 sg13g2_o21ai_1 _17596_ (.B1(_10616_),
    .Y(_01434_),
    .A1(_10441_),
    .A2(net364));
 sg13g2_nand2_1 _17597_ (.Y(_10617_),
    .A(\top_ihp.oisc.regs[3][29] ),
    .B(_10609_));
 sg13g2_o21ai_1 _17598_ (.B1(_10617_),
    .Y(_01435_),
    .A1(net53),
    .A2(net364));
 sg13g2_nand2_1 _17599_ (.Y(_10618_),
    .A(\top_ihp.oisc.regs[3][2] ),
    .B(net520));
 sg13g2_o21ai_1 _17600_ (.B1(_10618_),
    .Y(_01436_),
    .A1(_10493_),
    .A2(net364));
 sg13g2_nand2_1 _17601_ (.Y(_10619_),
    .A(\top_ihp.oisc.regs[3][30] ),
    .B(net520));
 sg13g2_o21ai_1 _17602_ (.B1(_10619_),
    .Y(_01437_),
    .A1(_10495_),
    .A2(_10595_));
 sg13g2_nand2_1 _17603_ (.Y(_10620_),
    .A(\top_ihp.oisc.regs[3][31] ),
    .B(_10593_));
 sg13g2_o21ai_1 _17604_ (.B1(_10620_),
    .Y(_01438_),
    .A1(_10540_),
    .A2(_10595_));
 sg13g2_nand2_1 _17605_ (.Y(_10621_),
    .A(\top_ihp.oisc.regs[3][3] ),
    .B(net523));
 sg13g2_o21ai_1 _17606_ (.B1(_10621_),
    .Y(_01439_),
    .A1(net118),
    .A2(net522));
 sg13g2_nand2_1 _17607_ (.Y(_10622_),
    .A(\top_ihp.oisc.regs[3][4] ),
    .B(net523));
 sg13g2_o21ai_1 _17608_ (.B1(_10622_),
    .Y(_01440_),
    .A1(_10500_),
    .A2(net522));
 sg13g2_nand2_1 _17609_ (.Y(_10623_),
    .A(\top_ihp.oisc.regs[3][5] ),
    .B(net523));
 sg13g2_o21ai_1 _17610_ (.B1(_10623_),
    .Y(_01441_),
    .A1(_10450_),
    .A2(net522));
 sg13g2_nand2_1 _17611_ (.Y(_10624_),
    .A(\top_ihp.oisc.regs[3][6] ),
    .B(net523));
 sg13g2_o21ai_1 _17612_ (.B1(_10624_),
    .Y(_01442_),
    .A1(_10452_),
    .A2(net522));
 sg13g2_nand2_1 _17613_ (.Y(_10625_),
    .A(\top_ihp.oisc.regs[3][7] ),
    .B(net523));
 sg13g2_o21ai_1 _17614_ (.B1(_10625_),
    .Y(_01443_),
    .A1(net209),
    .A2(net522));
 sg13g2_nand2_1 _17615_ (.Y(_10626_),
    .A(\top_ihp.oisc.regs[3][8] ),
    .B(net523));
 sg13g2_o21ai_1 _17616_ (.B1(_10626_),
    .Y(_01444_),
    .A1(net36),
    .A2(net522));
 sg13g2_nand2_1 _17617_ (.Y(_10627_),
    .A(\top_ihp.oisc.regs[3][9] ),
    .B(net523));
 sg13g2_o21ai_1 _17618_ (.B1(_10627_),
    .Y(_01445_),
    .A1(_10457_),
    .A2(net522));
 sg13g2_nand2b_1 _17619_ (.Y(_10628_),
    .B(_10401_),
    .A_N(_09956_));
 sg13g2_buf_1 _17620_ (.A(_10628_),
    .X(_10629_));
 sg13g2_buf_1 _17621_ (.A(net519),
    .X(_10630_));
 sg13g2_mux2_1 _17622_ (.A0(net407),
    .A1(\top_ihp.oisc.regs[40][0] ),
    .S(net363),
    .X(_01446_));
 sg13g2_nand2_1 _17623_ (.Y(_10631_),
    .A(net545),
    .B(_10401_));
 sg13g2_buf_2 _17624_ (.A(_10631_),
    .X(_10632_));
 sg13g2_nand2_1 _17625_ (.Y(_10633_),
    .A(\top_ihp.oisc.regs[40][10] ),
    .B(net363));
 sg13g2_o21ai_1 _17626_ (.B1(_10633_),
    .Y(_01447_),
    .A1(net39),
    .A2(_10632_));
 sg13g2_buf_1 _17627_ (.A(net519),
    .X(_10634_));
 sg13g2_nand2_1 _17628_ (.Y(_10635_),
    .A(\top_ihp.oisc.regs[40][11] ),
    .B(_10634_));
 sg13g2_o21ai_1 _17629_ (.B1(_10635_),
    .Y(_01448_),
    .A1(net121),
    .A2(_10632_));
 sg13g2_buf_1 _17630_ (.A(net519),
    .X(_10636_));
 sg13g2_nand2_1 _17631_ (.Y(_10637_),
    .A(\top_ihp.oisc.regs[40][12] ),
    .B(net362));
 sg13g2_o21ai_1 _17632_ (.B1(_10637_),
    .Y(_01449_),
    .A1(_10413_),
    .A2(net361));
 sg13g2_and2_1 _17633_ (.A(net545),
    .B(_10401_),
    .X(_10638_));
 sg13g2_buf_1 _17634_ (.A(_10638_),
    .X(_10639_));
 sg13g2_nor2_1 _17635_ (.A(\top_ihp.oisc.regs[40][13] ),
    .B(net201),
    .Y(_10640_));
 sg13g2_a21oi_1 _17636_ (.A1(net59),
    .A2(net201),
    .Y(_01450_),
    .B1(_10640_));
 sg13g2_nand2_1 _17637_ (.Y(_10641_),
    .A(\top_ihp.oisc.regs[40][14] ),
    .B(_10634_));
 sg13g2_o21ai_1 _17638_ (.B1(_10641_),
    .Y(_01451_),
    .A1(net127),
    .A2(_10636_));
 sg13g2_nand2_1 _17639_ (.Y(_10642_),
    .A(\top_ihp.oisc.regs[40][15] ),
    .B(net362));
 sg13g2_o21ai_1 _17640_ (.B1(_10642_),
    .Y(_01452_),
    .A1(net120),
    .A2(net361));
 sg13g2_nor2_1 _17641_ (.A(\top_ihp.oisc.regs[40][16] ),
    .B(net201),
    .Y(_10643_));
 sg13g2_a21oi_1 _17642_ (.A1(net132),
    .A2(net201),
    .Y(_01453_),
    .B1(_10643_));
 sg13g2_nand2_1 _17643_ (.Y(_10644_),
    .A(\top_ihp.oisc.regs[40][17] ),
    .B(net362));
 sg13g2_o21ai_1 _17644_ (.B1(_10644_),
    .Y(_01454_),
    .A1(net57),
    .A2(net361));
 sg13g2_nand2_1 _17645_ (.Y(_10645_),
    .A(\top_ihp.oisc.regs[40][18] ),
    .B(net362));
 sg13g2_o21ai_1 _17646_ (.B1(_10645_),
    .Y(_01455_),
    .A1(net56),
    .A2(net361));
 sg13g2_nand2_1 _17647_ (.Y(_10646_),
    .A(\top_ihp.oisc.regs[40][19] ),
    .B(net362));
 sg13g2_o21ai_1 _17648_ (.B1(_10646_),
    .Y(_01456_),
    .A1(net126),
    .A2(net361));
 sg13g2_nand2_1 _17649_ (.Y(_10647_),
    .A(\top_ihp.oisc.regs[40][1] ),
    .B(net362));
 sg13g2_o21ai_1 _17650_ (.B1(_10647_),
    .Y(_01457_),
    .A1(net380),
    .A2(net361));
 sg13g2_nor2_1 _17651_ (.A(\top_ihp.oisc.regs[40][20] ),
    .B(_10639_),
    .Y(_10648_));
 sg13g2_a21oi_1 _17652_ (.A1(net40),
    .A2(_10639_),
    .Y(_01458_),
    .B1(_10648_));
 sg13g2_nand2_1 _17653_ (.Y(_10649_),
    .A(\top_ihp.oisc.regs[40][21] ),
    .B(net362));
 sg13g2_o21ai_1 _17654_ (.B1(_10649_),
    .Y(_01459_),
    .A1(net38),
    .A2(_10636_));
 sg13g2_nor2_1 _17655_ (.A(\top_ihp.oisc.regs[40][22] ),
    .B(net201),
    .Y(_10650_));
 sg13g2_a21oi_1 _17656_ (.A1(net131),
    .A2(net201),
    .Y(_01460_),
    .B1(_10650_));
 sg13g2_nor2_1 _17657_ (.A(\top_ihp.oisc.regs[40][23] ),
    .B(net201),
    .Y(_10651_));
 sg13g2_a21oi_1 _17658_ (.A1(net138),
    .A2(net201),
    .Y(_01461_),
    .B1(_10651_));
 sg13g2_nand2_1 _17659_ (.Y(_10652_),
    .A(\top_ihp.oisc.regs[40][24] ),
    .B(net362));
 sg13g2_o21ai_1 _17660_ (.B1(_10652_),
    .Y(_01462_),
    .A1(net125),
    .A2(_10632_));
 sg13g2_buf_1 _17661_ (.A(net519),
    .X(_10653_));
 sg13g2_nand2_1 _17662_ (.Y(_10654_),
    .A(\top_ihp.oisc.regs[40][25] ),
    .B(net360));
 sg13g2_o21ai_1 _17663_ (.B1(_10654_),
    .Y(_01463_),
    .A1(net124),
    .A2(net361));
 sg13g2_nand2_1 _17664_ (.Y(_10655_),
    .A(\top_ihp.oisc.regs[40][26] ),
    .B(net360));
 sg13g2_o21ai_1 _17665_ (.B1(_10655_),
    .Y(_01464_),
    .A1(net55),
    .A2(net361));
 sg13g2_nand2_1 _17666_ (.Y(_10656_),
    .A(\top_ihp.oisc.regs[40][27] ),
    .B(net360));
 sg13g2_o21ai_1 _17667_ (.B1(_10656_),
    .Y(_01465_),
    .A1(_10439_),
    .A2(_10632_));
 sg13g2_nand2_1 _17668_ (.Y(_10657_),
    .A(\top_ihp.oisc.regs[40][28] ),
    .B(net360));
 sg13g2_o21ai_1 _17669_ (.B1(_10657_),
    .Y(_01466_),
    .A1(net37),
    .A2(net363));
 sg13g2_nand2_1 _17670_ (.Y(_10658_),
    .A(\top_ihp.oisc.regs[40][29] ),
    .B(net360));
 sg13g2_o21ai_1 _17671_ (.B1(_10658_),
    .Y(_01467_),
    .A1(_10443_),
    .A2(_10630_));
 sg13g2_nand2_1 _17672_ (.Y(_10659_),
    .A(\top_ihp.oisc.regs[40][2] ),
    .B(net360));
 sg13g2_o21ai_1 _17673_ (.B1(_10659_),
    .Y(_01468_),
    .A1(net119),
    .A2(net363));
 sg13g2_nand2_1 _17674_ (.Y(_10660_),
    .A(\top_ihp.oisc.regs[40][30] ),
    .B(net360));
 sg13g2_o21ai_1 _17675_ (.B1(_10660_),
    .Y(_01469_),
    .A1(net34),
    .A2(_10630_));
 sg13g2_nand2_1 _17676_ (.Y(_10661_),
    .A(\top_ihp.oisc.regs[40][31] ),
    .B(net360));
 sg13g2_o21ai_1 _17677_ (.B1(_10661_),
    .Y(_01470_),
    .A1(net116),
    .A2(_10632_));
 sg13g2_nand2_1 _17678_ (.Y(_10662_),
    .A(\top_ihp.oisc.regs[40][3] ),
    .B(_10653_));
 sg13g2_o21ai_1 _17679_ (.B1(_10662_),
    .Y(_01471_),
    .A1(net118),
    .A2(net363));
 sg13g2_nand2_1 _17680_ (.Y(_10663_),
    .A(\top_ihp.oisc.regs[40][4] ),
    .B(_10653_));
 sg13g2_o21ai_1 _17681_ (.B1(_10663_),
    .Y(_01472_),
    .A1(net117),
    .A2(_10632_));
 sg13g2_nand2_1 _17682_ (.Y(_10664_),
    .A(\top_ihp.oisc.regs[40][5] ),
    .B(net519));
 sg13g2_o21ai_1 _17683_ (.B1(_10664_),
    .Y(_01473_),
    .A1(net123),
    .A2(net363));
 sg13g2_nand2_1 _17684_ (.Y(_10665_),
    .A(\top_ihp.oisc.regs[40][6] ),
    .B(net519));
 sg13g2_o21ai_1 _17685_ (.B1(_10665_),
    .Y(_01474_),
    .A1(net122),
    .A2(net363));
 sg13g2_nand2_1 _17686_ (.Y(_10666_),
    .A(\top_ihp.oisc.regs[40][7] ),
    .B(_10629_));
 sg13g2_o21ai_1 _17687_ (.B1(_10666_),
    .Y(_01475_),
    .A1(_10189_),
    .A2(net363));
 sg13g2_nand2_1 _17688_ (.Y(_10667_),
    .A(\top_ihp.oisc.regs[40][8] ),
    .B(net519));
 sg13g2_o21ai_1 _17689_ (.B1(_10667_),
    .Y(_01476_),
    .A1(net36),
    .A2(_10632_));
 sg13g2_nand2_1 _17690_ (.Y(_10668_),
    .A(\top_ihp.oisc.regs[40][9] ),
    .B(net519));
 sg13g2_o21ai_1 _17691_ (.B1(_10668_),
    .Y(_01477_),
    .A1(net35),
    .A2(_10632_));
 sg13g2_nor2_2 _17692_ (.A(_09958_),
    .B(_10276_),
    .Y(_10669_));
 sg13g2_mux2_1 _17693_ (.A0(\top_ihp.oisc.regs[41][0] ),
    .A1(net204),
    .S(_10669_),
    .X(_01478_));
 sg13g2_or2_1 _17694_ (.X(_10670_),
    .B(_10276_),
    .A(_09958_));
 sg13g2_buf_1 _17695_ (.A(_10670_),
    .X(_10671_));
 sg13g2_buf_8 _17696_ (.A(_10671_),
    .X(_10672_));
 sg13g2_buf_1 _17697_ (.A(net200),
    .X(_10673_));
 sg13g2_buf_2 _17698_ (.A(_10671_),
    .X(_10674_));
 sg13g2_nand2_1 _17699_ (.Y(_10675_),
    .A(\top_ihp.oisc.regs[41][10] ),
    .B(net199));
 sg13g2_o21ai_1 _17700_ (.B1(_10675_),
    .Y(_01479_),
    .A1(net39),
    .A2(net115));
 sg13g2_buf_1 _17701_ (.A(_10671_),
    .X(_10676_));
 sg13g2_nand2_1 _17702_ (.Y(_10677_),
    .A(\top_ihp.oisc.regs[41][11] ),
    .B(net198));
 sg13g2_o21ai_1 _17703_ (.B1(_10677_),
    .Y(_01480_),
    .A1(net121),
    .A2(net115));
 sg13g2_nand2_1 _17704_ (.Y(_10678_),
    .A(\top_ihp.oisc.regs[41][12] ),
    .B(net198));
 sg13g2_o21ai_1 _17705_ (.B1(_10678_),
    .Y(_01481_),
    .A1(net128),
    .A2(net115));
 sg13g2_nand2_1 _17706_ (.Y(_10679_),
    .A(\top_ihp.oisc.regs[41][13] ),
    .B(_10676_));
 sg13g2_o21ai_1 _17707_ (.B1(_10679_),
    .Y(_01482_),
    .A1(_10203_),
    .A2(_10673_));
 sg13g2_nand2_1 _17708_ (.Y(_10680_),
    .A(\top_ihp.oisc.regs[41][14] ),
    .B(net198));
 sg13g2_o21ai_1 _17709_ (.B1(_10680_),
    .Y(_01483_),
    .A1(net127),
    .A2(net115));
 sg13g2_nand2_1 _17710_ (.Y(_10681_),
    .A(\top_ihp.oisc.regs[41][15] ),
    .B(net198));
 sg13g2_o21ai_1 _17711_ (.B1(_10681_),
    .Y(_01484_),
    .A1(net120),
    .A2(net115));
 sg13g2_nand2_1 _17712_ (.Y(_10682_),
    .A(\top_ihp.oisc.regs[41][16] ),
    .B(net198));
 sg13g2_o21ai_1 _17713_ (.B1(_10682_),
    .Y(_01485_),
    .A1(_10163_),
    .A2(_10673_));
 sg13g2_nand2_1 _17714_ (.Y(_10683_),
    .A(\top_ihp.oisc.regs[41][17] ),
    .B(net198));
 sg13g2_o21ai_1 _17715_ (.B1(_10683_),
    .Y(_01486_),
    .A1(net57),
    .A2(net115));
 sg13g2_nand2_1 _17716_ (.Y(_10684_),
    .A(\top_ihp.oisc.regs[41][18] ),
    .B(net198));
 sg13g2_o21ai_1 _17717_ (.B1(_10684_),
    .Y(_01487_),
    .A1(net56),
    .A2(net115));
 sg13g2_nand2_1 _17718_ (.Y(_10685_),
    .A(\top_ihp.oisc.regs[41][19] ),
    .B(_10676_));
 sg13g2_o21ai_1 _17719_ (.B1(_10685_),
    .Y(_01488_),
    .A1(_10424_),
    .A2(net115));
 sg13g2_buf_1 _17720_ (.A(net200),
    .X(_10686_));
 sg13g2_nand2_1 _17721_ (.Y(_10687_),
    .A(\top_ihp.oisc.regs[41][1] ),
    .B(net198));
 sg13g2_o21ai_1 _17722_ (.B1(_10687_),
    .Y(_01489_),
    .A1(net380),
    .A2(net114));
 sg13g2_mux2_1 _17723_ (.A0(\top_ihp.oisc.regs[41][20] ),
    .A1(net137),
    .S(_10669_),
    .X(_01490_));
 sg13g2_buf_1 _17724_ (.A(_10671_),
    .X(_10688_));
 sg13g2_nand2_1 _17725_ (.Y(_10689_),
    .A(\top_ihp.oisc.regs[41][21] ),
    .B(net197));
 sg13g2_o21ai_1 _17726_ (.B1(_10689_),
    .Y(_01491_),
    .A1(net38),
    .A2(net114));
 sg13g2_nand2_1 _17727_ (.Y(_10690_),
    .A(\top_ihp.oisc.regs[41][22] ),
    .B(net197));
 sg13g2_o21ai_1 _17728_ (.B1(_10690_),
    .Y(_01492_),
    .A1(net129),
    .A2(net114));
 sg13g2_mux2_1 _17729_ (.A0(\top_ihp.oisc.regs[41][23] ),
    .A1(_10036_),
    .S(_10669_),
    .X(_01493_));
 sg13g2_nand2_1 _17730_ (.Y(_10691_),
    .A(\top_ihp.oisc.regs[41][24] ),
    .B(net197));
 sg13g2_o21ai_1 _17731_ (.B1(_10691_),
    .Y(_01494_),
    .A1(net125),
    .A2(net114));
 sg13g2_nand2_1 _17732_ (.Y(_10692_),
    .A(\top_ihp.oisc.regs[41][25] ),
    .B(net197));
 sg13g2_o21ai_1 _17733_ (.B1(_10692_),
    .Y(_01495_),
    .A1(net124),
    .A2(net114));
 sg13g2_nand2_1 _17734_ (.Y(_10693_),
    .A(\top_ihp.oisc.regs[41][26] ),
    .B(net197));
 sg13g2_o21ai_1 _17735_ (.B1(_10693_),
    .Y(_01496_),
    .A1(net55),
    .A2(net114));
 sg13g2_nand2_1 _17736_ (.Y(_10694_),
    .A(\top_ihp.oisc.regs[41][27] ),
    .B(net197));
 sg13g2_o21ai_1 _17737_ (.B1(_10694_),
    .Y(_01497_),
    .A1(net54),
    .A2(_10686_));
 sg13g2_nand2_1 _17738_ (.Y(_10695_),
    .A(\top_ihp.oisc.regs[41][28] ),
    .B(net197));
 sg13g2_o21ai_1 _17739_ (.B1(_10695_),
    .Y(_01498_),
    .A1(net37),
    .A2(_10686_));
 sg13g2_nand2_1 _17740_ (.Y(_10696_),
    .A(\top_ihp.oisc.regs[41][29] ),
    .B(net197));
 sg13g2_o21ai_1 _17741_ (.B1(_10696_),
    .Y(_01499_),
    .A1(net53),
    .A2(net114));
 sg13g2_nand2_1 _17742_ (.Y(_10697_),
    .A(\top_ihp.oisc.regs[41][2] ),
    .B(_10688_));
 sg13g2_o21ai_1 _17743_ (.B1(_10697_),
    .Y(_01500_),
    .A1(net119),
    .A2(net114));
 sg13g2_nand2_1 _17744_ (.Y(_10698_),
    .A(\top_ihp.oisc.regs[41][30] ),
    .B(_10688_));
 sg13g2_o21ai_1 _17745_ (.B1(_10698_),
    .Y(_01501_),
    .A1(net34),
    .A2(net199));
 sg13g2_nand2_1 _17746_ (.Y(_10699_),
    .A(\top_ihp.oisc.regs[41][31] ),
    .B(net200));
 sg13g2_o21ai_1 _17747_ (.B1(_10699_),
    .Y(_01502_),
    .A1(_10540_),
    .A2(net199));
 sg13g2_nand2_1 _17748_ (.Y(_10700_),
    .A(\top_ihp.oisc.regs[41][3] ),
    .B(net200));
 sg13g2_o21ai_1 _17749_ (.B1(_10700_),
    .Y(_01503_),
    .A1(_10498_),
    .A2(net199));
 sg13g2_nand2_1 _17750_ (.Y(_10701_),
    .A(\top_ihp.oisc.regs[41][4] ),
    .B(net200));
 sg13g2_o21ai_1 _17751_ (.B1(_10701_),
    .Y(_01504_),
    .A1(net117),
    .A2(net199));
 sg13g2_nand2_1 _17752_ (.Y(_10702_),
    .A(\top_ihp.oisc.regs[41][5] ),
    .B(_10672_));
 sg13g2_o21ai_1 _17753_ (.B1(_10702_),
    .Y(_01505_),
    .A1(net123),
    .A2(net199));
 sg13g2_nand2_1 _17754_ (.Y(_10703_),
    .A(\top_ihp.oisc.regs[41][6] ),
    .B(net200));
 sg13g2_o21ai_1 _17755_ (.B1(_10703_),
    .Y(_01506_),
    .A1(net122),
    .A2(_10674_));
 sg13g2_nand2_1 _17756_ (.Y(_10704_),
    .A(\top_ihp.oisc.regs[41][7] ),
    .B(_10672_));
 sg13g2_o21ai_1 _17757_ (.B1(_10704_),
    .Y(_01507_),
    .A1(net68),
    .A2(_10674_));
 sg13g2_nand2_1 _17758_ (.Y(_10705_),
    .A(\top_ihp.oisc.regs[41][8] ),
    .B(net200));
 sg13g2_o21ai_1 _17759_ (.B1(_10705_),
    .Y(_01508_),
    .A1(_10455_),
    .A2(net199));
 sg13g2_nand2_1 _17760_ (.Y(_10706_),
    .A(\top_ihp.oisc.regs[41][9] ),
    .B(net200));
 sg13g2_o21ai_1 _17761_ (.B1(_10706_),
    .Y(_01509_),
    .A1(net35),
    .A2(net199));
 sg13g2_nand2b_1 _17762_ (.Y(_10707_),
    .B(net664),
    .A_N(_09956_));
 sg13g2_buf_2 _17763_ (.A(_10707_),
    .X(_10708_));
 sg13g2_buf_2 _17764_ (.A(_10708_),
    .X(_10709_));
 sg13g2_mux2_1 _17765_ (.A0(net407),
    .A1(\top_ihp.oisc.regs[42][0] ),
    .S(_10709_),
    .X(_01510_));
 sg13g2_nand2_1 _17766_ (.Y(_10710_),
    .A(net545),
    .B(net664));
 sg13g2_buf_1 _17767_ (.A(_10710_),
    .X(_10711_));
 sg13g2_nand2_1 _17768_ (.Y(_10712_),
    .A(\top_ihp.oisc.regs[42][10] ),
    .B(net359));
 sg13g2_o21ai_1 _17769_ (.B1(_10712_),
    .Y(_01511_),
    .A1(net39),
    .A2(net196));
 sg13g2_nand2_1 _17770_ (.Y(_10713_),
    .A(\top_ihp.oisc.regs[42][11] ),
    .B(net359));
 sg13g2_o21ai_1 _17771_ (.B1(_10713_),
    .Y(_01512_),
    .A1(net121),
    .A2(net196));
 sg13g2_buf_2 _17772_ (.A(_10708_),
    .X(_10714_));
 sg13g2_buf_2 _17773_ (.A(_10708_),
    .X(_10715_));
 sg13g2_nand2_1 _17774_ (.Y(_10716_),
    .A(\top_ihp.oisc.regs[42][12] ),
    .B(net357));
 sg13g2_o21ai_1 _17775_ (.B1(_10716_),
    .Y(_01513_),
    .A1(net128),
    .A2(net358));
 sg13g2_and2_1 _17776_ (.A(net545),
    .B(net664),
    .X(_10717_));
 sg13g2_buf_1 _17777_ (.A(_10717_),
    .X(_10718_));
 sg13g2_nor2_1 _17778_ (.A(\top_ihp.oisc.regs[42][13] ),
    .B(net195),
    .Y(_10719_));
 sg13g2_a21oi_1 _17779_ (.A1(net59),
    .A2(net195),
    .Y(_01514_),
    .B1(_10719_));
 sg13g2_nand2_1 _17780_ (.Y(_10720_),
    .A(\top_ihp.oisc.regs[42][14] ),
    .B(net357));
 sg13g2_o21ai_1 _17781_ (.B1(_10720_),
    .Y(_01515_),
    .A1(net127),
    .A2(net358));
 sg13g2_nand2_1 _17782_ (.Y(_10721_),
    .A(\top_ihp.oisc.regs[42][15] ),
    .B(net357));
 sg13g2_o21ai_1 _17783_ (.B1(_10721_),
    .Y(_01516_),
    .A1(_10473_),
    .A2(net358));
 sg13g2_nor2_1 _17784_ (.A(\top_ihp.oisc.regs[42][16] ),
    .B(_10718_),
    .Y(_10722_));
 sg13g2_a21oi_1 _17785_ (.A1(net132),
    .A2(_10718_),
    .Y(_01517_),
    .B1(_10722_));
 sg13g2_nand2_1 _17786_ (.Y(_10723_),
    .A(\top_ihp.oisc.regs[42][17] ),
    .B(net357));
 sg13g2_o21ai_1 _17787_ (.B1(_10723_),
    .Y(_01518_),
    .A1(net57),
    .A2(net358));
 sg13g2_nand2_1 _17788_ (.Y(_10724_),
    .A(\top_ihp.oisc.regs[42][18] ),
    .B(net357));
 sg13g2_o21ai_1 _17789_ (.B1(_10724_),
    .Y(_01519_),
    .A1(net56),
    .A2(net358));
 sg13g2_nand2_1 _17790_ (.Y(_10725_),
    .A(\top_ihp.oisc.regs[42][19] ),
    .B(net357));
 sg13g2_o21ai_1 _17791_ (.B1(_10725_),
    .Y(_01520_),
    .A1(net126),
    .A2(net358));
 sg13g2_nand2_1 _17792_ (.Y(_10726_),
    .A(\top_ihp.oisc.regs[42][1] ),
    .B(_10715_));
 sg13g2_o21ai_1 _17793_ (.B1(_10726_),
    .Y(_01521_),
    .A1(net380),
    .A2(net358));
 sg13g2_nor2_1 _17794_ (.A(\top_ihp.oisc.regs[42][20] ),
    .B(net195),
    .Y(_10727_));
 sg13g2_a21oi_1 _17795_ (.A1(_09981_),
    .A2(net195),
    .Y(_01522_),
    .B1(_10727_));
 sg13g2_nand2_1 _17796_ (.Y(_10728_),
    .A(\top_ihp.oisc.regs[42][21] ),
    .B(net357));
 sg13g2_o21ai_1 _17797_ (.B1(_10728_),
    .Y(_01523_),
    .A1(net38),
    .A2(net358));
 sg13g2_nor2_1 _17798_ (.A(\top_ihp.oisc.regs[42][22] ),
    .B(net195),
    .Y(_10729_));
 sg13g2_a21oi_1 _17799_ (.A1(net131),
    .A2(net195),
    .Y(_01524_),
    .B1(_10729_));
 sg13g2_nor2_1 _17800_ (.A(\top_ihp.oisc.regs[42][23] ),
    .B(net195),
    .Y(_10730_));
 sg13g2_a21oi_1 _17801_ (.A1(net138),
    .A2(net195),
    .Y(_01525_),
    .B1(_10730_));
 sg13g2_nand2_1 _17802_ (.Y(_10731_),
    .A(\top_ihp.oisc.regs[42][24] ),
    .B(net357));
 sg13g2_o21ai_1 _17803_ (.B1(_10731_),
    .Y(_01526_),
    .A1(net125),
    .A2(net196));
 sg13g2_nand2_1 _17804_ (.Y(_10732_),
    .A(\top_ihp.oisc.regs[42][25] ),
    .B(_10715_));
 sg13g2_o21ai_1 _17805_ (.B1(_10732_),
    .Y(_01527_),
    .A1(net124),
    .A2(_10714_));
 sg13g2_buf_1 _17806_ (.A(_10708_),
    .X(_10733_));
 sg13g2_nand2_1 _17807_ (.Y(_10734_),
    .A(\top_ihp.oisc.regs[42][26] ),
    .B(net356));
 sg13g2_o21ai_1 _17808_ (.B1(_10734_),
    .Y(_01528_),
    .A1(_10437_),
    .A2(_10714_));
 sg13g2_nand2_1 _17809_ (.Y(_10735_),
    .A(\top_ihp.oisc.regs[42][27] ),
    .B(_10733_));
 sg13g2_o21ai_1 _17810_ (.B1(_10735_),
    .Y(_01529_),
    .A1(net54),
    .A2(_10711_));
 sg13g2_nand2_1 _17811_ (.Y(_10736_),
    .A(\top_ihp.oisc.regs[42][28] ),
    .B(net356));
 sg13g2_o21ai_1 _17812_ (.B1(_10736_),
    .Y(_01530_),
    .A1(net37),
    .A2(net359));
 sg13g2_nand2_1 _17813_ (.Y(_10737_),
    .A(\top_ihp.oisc.regs[42][29] ),
    .B(_10733_));
 sg13g2_o21ai_1 _17814_ (.B1(_10737_),
    .Y(_01531_),
    .A1(net53),
    .A2(net359));
 sg13g2_nand2_1 _17815_ (.Y(_10738_),
    .A(\top_ihp.oisc.regs[42][2] ),
    .B(net356));
 sg13g2_o21ai_1 _17816_ (.B1(_10738_),
    .Y(_01532_),
    .A1(net119),
    .A2(net359));
 sg13g2_nand2_1 _17817_ (.Y(_10739_),
    .A(\top_ihp.oisc.regs[42][30] ),
    .B(net356));
 sg13g2_o21ai_1 _17818_ (.B1(_10739_),
    .Y(_01533_),
    .A1(net34),
    .A2(_10709_));
 sg13g2_nand2_1 _17819_ (.Y(_10740_),
    .A(\top_ihp.oisc.regs[42][31] ),
    .B(net356));
 sg13g2_o21ai_1 _17820_ (.B1(_10740_),
    .Y(_01534_),
    .A1(net116),
    .A2(net196));
 sg13g2_nand2_1 _17821_ (.Y(_10741_),
    .A(\top_ihp.oisc.regs[42][3] ),
    .B(net356));
 sg13g2_o21ai_1 _17822_ (.B1(_10741_),
    .Y(_01535_),
    .A1(net118),
    .A2(net359));
 sg13g2_nand2_1 _17823_ (.Y(_10742_),
    .A(\top_ihp.oisc.regs[42][4] ),
    .B(net356));
 sg13g2_o21ai_1 _17824_ (.B1(_10742_),
    .Y(_01536_),
    .A1(net117),
    .A2(net196));
 sg13g2_nand2_1 _17825_ (.Y(_10743_),
    .A(\top_ihp.oisc.regs[42][5] ),
    .B(net356));
 sg13g2_o21ai_1 _17826_ (.B1(_10743_),
    .Y(_01537_),
    .A1(_10450_),
    .A2(net359));
 sg13g2_nand2_1 _17827_ (.Y(_10744_),
    .A(\top_ihp.oisc.regs[42][6] ),
    .B(_10708_));
 sg13g2_o21ai_1 _17828_ (.B1(_10744_),
    .Y(_01538_),
    .A1(net122),
    .A2(net359));
 sg13g2_nand2_1 _17829_ (.Y(_10745_),
    .A(\top_ihp.oisc.regs[42][7] ),
    .B(_10708_));
 sg13g2_o21ai_1 _17830_ (.B1(_10745_),
    .Y(_01539_),
    .A1(_09914_),
    .A2(net196));
 sg13g2_nand2_1 _17831_ (.Y(_10746_),
    .A(\top_ihp.oisc.regs[42][8] ),
    .B(_10708_));
 sg13g2_o21ai_1 _17832_ (.B1(_10746_),
    .Y(_01540_),
    .A1(net36),
    .A2(net196));
 sg13g2_nand2_1 _17833_ (.Y(_10747_),
    .A(\top_ihp.oisc.regs[42][9] ),
    .B(_10708_));
 sg13g2_o21ai_1 _17834_ (.B1(_10747_),
    .Y(_01541_),
    .A1(net35),
    .A2(net196));
 sg13g2_and2_1 _17835_ (.A(_10029_),
    .B(_10358_),
    .X(_10748_));
 sg13g2_buf_1 _17836_ (.A(_10748_),
    .X(_10749_));
 sg13g2_mux2_1 _17837_ (.A0(\top_ihp.oisc.regs[43][0] ),
    .A1(net204),
    .S(_10749_),
    .X(_01542_));
 sg13g2_nand2_1 _17838_ (.Y(_10750_),
    .A(_10007_),
    .B(_10358_));
 sg13g2_buf_1 _17839_ (.A(_10750_),
    .X(_10751_));
 sg13g2_buf_1 _17840_ (.A(_10751_),
    .X(_10752_));
 sg13g2_buf_1 _17841_ (.A(_10752_),
    .X(_10753_));
 sg13g2_buf_1 _17842_ (.A(_10751_),
    .X(_10754_));
 sg13g2_nand2_1 _17843_ (.Y(_10755_),
    .A(\top_ihp.oisc.regs[43][10] ),
    .B(net193));
 sg13g2_o21ai_1 _17844_ (.B1(_10755_),
    .Y(_01543_),
    .A1(net39),
    .A2(_10753_));
 sg13g2_buf_1 _17845_ (.A(_10751_),
    .X(_10756_));
 sg13g2_nand2_1 _17846_ (.Y(_10757_),
    .A(\top_ihp.oisc.regs[43][11] ),
    .B(_10756_));
 sg13g2_o21ai_1 _17847_ (.B1(_10757_),
    .Y(_01544_),
    .A1(net121),
    .A2(net113));
 sg13g2_nand2_1 _17848_ (.Y(_10758_),
    .A(\top_ihp.oisc.regs[43][12] ),
    .B(_10756_));
 sg13g2_o21ai_1 _17849_ (.B1(_10758_),
    .Y(_01545_),
    .A1(_10413_),
    .A2(net113));
 sg13g2_nand2_1 _17850_ (.Y(_10759_),
    .A(\top_ihp.oisc.regs[43][13] ),
    .B(net192));
 sg13g2_o21ai_1 _17851_ (.B1(_10759_),
    .Y(_01546_),
    .A1(_10203_),
    .A2(net113));
 sg13g2_nand2_1 _17852_ (.Y(_10760_),
    .A(\top_ihp.oisc.regs[43][14] ),
    .B(net192));
 sg13g2_o21ai_1 _17853_ (.B1(_10760_),
    .Y(_01547_),
    .A1(net127),
    .A2(net113));
 sg13g2_nand2_1 _17854_ (.Y(_10761_),
    .A(\top_ihp.oisc.regs[43][15] ),
    .B(net192));
 sg13g2_o21ai_1 _17855_ (.B1(_10761_),
    .Y(_01548_),
    .A1(net120),
    .A2(net113));
 sg13g2_buf_2 _17856_ (.A(_09435_),
    .X(_10762_));
 sg13g2_nand2_1 _17857_ (.Y(_10763_),
    .A(\top_ihp.oisc.regs[43][16] ),
    .B(net192));
 sg13g2_o21ai_1 _17858_ (.B1(_10763_),
    .Y(_01549_),
    .A1(net191),
    .A2(_10753_));
 sg13g2_nand2_1 _17859_ (.Y(_10764_),
    .A(\top_ihp.oisc.regs[43][17] ),
    .B(net192));
 sg13g2_o21ai_1 _17860_ (.B1(_10764_),
    .Y(_01550_),
    .A1(net57),
    .A2(net113));
 sg13g2_nand2_1 _17861_ (.Y(_10765_),
    .A(\top_ihp.oisc.regs[43][18] ),
    .B(net192));
 sg13g2_o21ai_1 _17862_ (.B1(_10765_),
    .Y(_01551_),
    .A1(net56),
    .A2(net113));
 sg13g2_nand2_1 _17863_ (.Y(_10766_),
    .A(\top_ihp.oisc.regs[43][19] ),
    .B(net192));
 sg13g2_o21ai_1 _17864_ (.B1(_10766_),
    .Y(_01552_),
    .A1(net126),
    .A2(net113));
 sg13g2_buf_1 _17865_ (.A(net194),
    .X(_10767_));
 sg13g2_nand2_1 _17866_ (.Y(_10768_),
    .A(\top_ihp.oisc.regs[43][1] ),
    .B(net192));
 sg13g2_o21ai_1 _17867_ (.B1(_10768_),
    .Y(_01553_),
    .A1(net380),
    .A2(net112));
 sg13g2_mux2_1 _17868_ (.A0(\top_ihp.oisc.regs[43][20] ),
    .A1(_10032_),
    .S(_10749_),
    .X(_01554_));
 sg13g2_buf_1 _17869_ (.A(_10751_),
    .X(_10769_));
 sg13g2_nand2_1 _17870_ (.Y(_10770_),
    .A(\top_ihp.oisc.regs[43][21] ),
    .B(net190));
 sg13g2_o21ai_1 _17871_ (.B1(_10770_),
    .Y(_01555_),
    .A1(net38),
    .A2(net112));
 sg13g2_nand2_1 _17872_ (.Y(_10771_),
    .A(\top_ihp.oisc.regs[43][22] ),
    .B(net190));
 sg13g2_o21ai_1 _17873_ (.B1(_10771_),
    .Y(_01556_),
    .A1(net129),
    .A2(net112));
 sg13g2_mux2_1 _17874_ (.A0(\top_ihp.oisc.regs[43][23] ),
    .A1(net406),
    .S(_10749_),
    .X(_01557_));
 sg13g2_nand2_1 _17875_ (.Y(_10772_),
    .A(\top_ihp.oisc.regs[43][24] ),
    .B(net190));
 sg13g2_o21ai_1 _17876_ (.B1(_10772_),
    .Y(_01558_),
    .A1(net125),
    .A2(net112));
 sg13g2_nand2_1 _17877_ (.Y(_10773_),
    .A(\top_ihp.oisc.regs[43][25] ),
    .B(net190));
 sg13g2_o21ai_1 _17878_ (.B1(_10773_),
    .Y(_01559_),
    .A1(_10435_),
    .A2(net112));
 sg13g2_nand2_1 _17879_ (.Y(_10774_),
    .A(\top_ihp.oisc.regs[43][26] ),
    .B(net190));
 sg13g2_o21ai_1 _17880_ (.B1(_10774_),
    .Y(_01560_),
    .A1(net55),
    .A2(_10767_));
 sg13g2_nand2_1 _17881_ (.Y(_10775_),
    .A(\top_ihp.oisc.regs[43][27] ),
    .B(net190));
 sg13g2_o21ai_1 _17882_ (.B1(_10775_),
    .Y(_01561_),
    .A1(net54),
    .A2(_10767_));
 sg13g2_nand2_1 _17883_ (.Y(_10776_),
    .A(\top_ihp.oisc.regs[43][28] ),
    .B(_10769_));
 sg13g2_o21ai_1 _17884_ (.B1(_10776_),
    .Y(_01562_),
    .A1(net37),
    .A2(net112));
 sg13g2_nand2_1 _17885_ (.Y(_10777_),
    .A(\top_ihp.oisc.regs[43][29] ),
    .B(net190));
 sg13g2_o21ai_1 _17886_ (.B1(_10777_),
    .Y(_01563_),
    .A1(_10443_),
    .A2(net112));
 sg13g2_nand2_1 _17887_ (.Y(_10778_),
    .A(\top_ihp.oisc.regs[43][2] ),
    .B(net190));
 sg13g2_o21ai_1 _17888_ (.B1(_10778_),
    .Y(_01564_),
    .A1(net119),
    .A2(net112));
 sg13g2_nand2_1 _17889_ (.Y(_10779_),
    .A(\top_ihp.oisc.regs[43][30] ),
    .B(_10769_));
 sg13g2_o21ai_1 _17890_ (.B1(_10779_),
    .Y(_01565_),
    .A1(net34),
    .A2(_10754_));
 sg13g2_nand2_1 _17891_ (.Y(_10780_),
    .A(\top_ihp.oisc.regs[43][31] ),
    .B(net194));
 sg13g2_o21ai_1 _17892_ (.B1(_10780_),
    .Y(_01566_),
    .A1(net116),
    .A2(net193));
 sg13g2_nand2_1 _17893_ (.Y(_10781_),
    .A(\top_ihp.oisc.regs[43][3] ),
    .B(net194));
 sg13g2_o21ai_1 _17894_ (.B1(_10781_),
    .Y(_01567_),
    .A1(net118),
    .A2(_10754_));
 sg13g2_nand2_1 _17895_ (.Y(_10782_),
    .A(\top_ihp.oisc.regs[43][4] ),
    .B(net194));
 sg13g2_o21ai_1 _17896_ (.B1(_10782_),
    .Y(_01568_),
    .A1(net117),
    .A2(net193));
 sg13g2_nand2_1 _17897_ (.Y(_10783_),
    .A(\top_ihp.oisc.regs[43][5] ),
    .B(_10752_));
 sg13g2_o21ai_1 _17898_ (.B1(_10783_),
    .Y(_01569_),
    .A1(net123),
    .A2(net193));
 sg13g2_nand2_1 _17899_ (.Y(_10784_),
    .A(\top_ihp.oisc.regs[43][6] ),
    .B(net194));
 sg13g2_o21ai_1 _17900_ (.B1(_10784_),
    .Y(_01570_),
    .A1(net122),
    .A2(net193));
 sg13g2_nand2_1 _17901_ (.Y(_10785_),
    .A(\top_ihp.oisc.regs[43][7] ),
    .B(net194));
 sg13g2_o21ai_1 _17902_ (.B1(_10785_),
    .Y(_01571_),
    .A1(_09914_),
    .A2(net193));
 sg13g2_nand2_1 _17903_ (.Y(_10786_),
    .A(\top_ihp.oisc.regs[43][8] ),
    .B(net194));
 sg13g2_o21ai_1 _17904_ (.B1(_10786_),
    .Y(_01572_),
    .A1(net36),
    .A2(net193));
 sg13g2_nand2_1 _17905_ (.Y(_10787_),
    .A(\top_ihp.oisc.regs[43][9] ),
    .B(net194));
 sg13g2_o21ai_1 _17906_ (.B1(_10787_),
    .Y(_01573_),
    .A1(net35),
    .A2(net193));
 sg13g2_and2_1 _17907_ (.A(net665),
    .B(_10401_),
    .X(_10788_));
 sg13g2_buf_1 _17908_ (.A(_10788_),
    .X(_10789_));
 sg13g2_mux2_1 _17909_ (.A0(\top_ihp.oisc.regs[44][0] ),
    .A1(net204),
    .S(_10789_),
    .X(_01574_));
 sg13g2_nand2_1 _17910_ (.Y(_10790_),
    .A(_10055_),
    .B(_10401_));
 sg13g2_buf_1 _17911_ (.A(_10790_),
    .X(_10791_));
 sg13g2_buf_1 _17912_ (.A(_10791_),
    .X(_10792_));
 sg13g2_buf_1 _17913_ (.A(net355),
    .X(_10793_));
 sg13g2_buf_2 _17914_ (.A(_10791_),
    .X(_10794_));
 sg13g2_nand2_1 _17915_ (.Y(_10795_),
    .A(\top_ihp.oisc.regs[44][10] ),
    .B(net354));
 sg13g2_o21ai_1 _17916_ (.B1(_10795_),
    .Y(_01575_),
    .A1(net39),
    .A2(net189));
 sg13g2_buf_1 _17917_ (.A(_10791_),
    .X(_10796_));
 sg13g2_nand2_1 _17918_ (.Y(_10797_),
    .A(\top_ihp.oisc.regs[44][11] ),
    .B(_10796_));
 sg13g2_o21ai_1 _17919_ (.B1(_10797_),
    .Y(_01576_),
    .A1(net121),
    .A2(_10793_));
 sg13g2_nand2_1 _17920_ (.Y(_10798_),
    .A(\top_ihp.oisc.regs[44][12] ),
    .B(net353));
 sg13g2_o21ai_1 _17921_ (.B1(_10798_),
    .Y(_01577_),
    .A1(net128),
    .A2(net189));
 sg13g2_buf_2 _17922_ (.A(_09373_),
    .X(_10799_));
 sg13g2_nand2_1 _17923_ (.Y(_10800_),
    .A(\top_ihp.oisc.regs[44][13] ),
    .B(net353));
 sg13g2_o21ai_1 _17924_ (.B1(_10800_),
    .Y(_01578_),
    .A1(net111),
    .A2(net189));
 sg13g2_nand2_1 _17925_ (.Y(_10801_),
    .A(\top_ihp.oisc.regs[44][14] ),
    .B(_10796_));
 sg13g2_o21ai_1 _17926_ (.B1(_10801_),
    .Y(_01579_),
    .A1(net127),
    .A2(_10793_));
 sg13g2_nand2_1 _17927_ (.Y(_10802_),
    .A(\top_ihp.oisc.regs[44][15] ),
    .B(net353));
 sg13g2_o21ai_1 _17928_ (.B1(_10802_),
    .Y(_01580_),
    .A1(_10473_),
    .A2(net189));
 sg13g2_nand2_1 _17929_ (.Y(_10803_),
    .A(\top_ihp.oisc.regs[44][16] ),
    .B(net353));
 sg13g2_o21ai_1 _17930_ (.B1(_10803_),
    .Y(_01581_),
    .A1(net191),
    .A2(net189));
 sg13g2_nand2_1 _17931_ (.Y(_10804_),
    .A(\top_ihp.oisc.regs[44][17] ),
    .B(net353));
 sg13g2_o21ai_1 _17932_ (.B1(_10804_),
    .Y(_01582_),
    .A1(net57),
    .A2(net189));
 sg13g2_nand2_1 _17933_ (.Y(_10805_),
    .A(\top_ihp.oisc.regs[44][18] ),
    .B(net353));
 sg13g2_o21ai_1 _17934_ (.B1(_10805_),
    .Y(_01583_),
    .A1(net56),
    .A2(net189));
 sg13g2_nand2_1 _17935_ (.Y(_10806_),
    .A(\top_ihp.oisc.regs[44][19] ),
    .B(net353));
 sg13g2_o21ai_1 _17936_ (.B1(_10806_),
    .Y(_01584_),
    .A1(_10424_),
    .A2(net189));
 sg13g2_buf_1 _17937_ (.A(net355),
    .X(_10807_));
 sg13g2_nand2_1 _17938_ (.Y(_10808_),
    .A(\top_ihp.oisc.regs[44][1] ),
    .B(net353));
 sg13g2_o21ai_1 _17939_ (.B1(_10808_),
    .Y(_01585_),
    .A1(_10426_),
    .A2(net188));
 sg13g2_mux2_1 _17940_ (.A0(\top_ihp.oisc.regs[44][20] ),
    .A1(_10032_),
    .S(_10789_),
    .X(_01586_));
 sg13g2_buf_1 _17941_ (.A(_10791_),
    .X(_10809_));
 sg13g2_nand2_1 _17942_ (.Y(_10810_),
    .A(\top_ihp.oisc.regs[44][21] ),
    .B(net352));
 sg13g2_o21ai_1 _17943_ (.B1(_10810_),
    .Y(_01587_),
    .A1(_10429_),
    .A2(net188));
 sg13g2_buf_2 _17944_ (.A(net244),
    .X(_10811_));
 sg13g2_nand2_1 _17945_ (.Y(_10812_),
    .A(\top_ihp.oisc.regs[44][22] ),
    .B(net352));
 sg13g2_o21ai_1 _17946_ (.B1(_10812_),
    .Y(_01588_),
    .A1(net110),
    .A2(net188));
 sg13g2_mux2_1 _17947_ (.A0(\top_ihp.oisc.regs[44][23] ),
    .A1(net406),
    .S(_10789_),
    .X(_01589_));
 sg13g2_nand2_1 _17948_ (.Y(_10813_),
    .A(\top_ihp.oisc.regs[44][24] ),
    .B(_10809_));
 sg13g2_o21ai_1 _17949_ (.B1(_10813_),
    .Y(_01590_),
    .A1(net125),
    .A2(net188));
 sg13g2_nand2_1 _17950_ (.Y(_10814_),
    .A(\top_ihp.oisc.regs[44][25] ),
    .B(net352));
 sg13g2_o21ai_1 _17951_ (.B1(_10814_),
    .Y(_01591_),
    .A1(_10435_),
    .A2(net188));
 sg13g2_nand2_1 _17952_ (.Y(_10815_),
    .A(\top_ihp.oisc.regs[44][26] ),
    .B(net352));
 sg13g2_o21ai_1 _17953_ (.B1(_10815_),
    .Y(_01592_),
    .A1(_10437_),
    .A2(net188));
 sg13g2_nand2_1 _17954_ (.Y(_10816_),
    .A(\top_ihp.oisc.regs[44][27] ),
    .B(net352));
 sg13g2_o21ai_1 _17955_ (.B1(_10816_),
    .Y(_01593_),
    .A1(net54),
    .A2(_10807_));
 sg13g2_nand2_1 _17956_ (.Y(_10817_),
    .A(\top_ihp.oisc.regs[44][28] ),
    .B(_10809_));
 sg13g2_o21ai_1 _17957_ (.B1(_10817_),
    .Y(_01594_),
    .A1(net37),
    .A2(_10807_));
 sg13g2_nand2_1 _17958_ (.Y(_10818_),
    .A(\top_ihp.oisc.regs[44][29] ),
    .B(net352));
 sg13g2_o21ai_1 _17959_ (.B1(_10818_),
    .Y(_01595_),
    .A1(net53),
    .A2(net188));
 sg13g2_nand2_1 _17960_ (.Y(_10819_),
    .A(\top_ihp.oisc.regs[44][2] ),
    .B(net352));
 sg13g2_o21ai_1 _17961_ (.B1(_10819_),
    .Y(_01596_),
    .A1(net119),
    .A2(net188));
 sg13g2_nand2_1 _17962_ (.Y(_10820_),
    .A(\top_ihp.oisc.regs[44][30] ),
    .B(net352));
 sg13g2_o21ai_1 _17963_ (.B1(_10820_),
    .Y(_01597_),
    .A1(net34),
    .A2(net354));
 sg13g2_nand2_1 _17964_ (.Y(_10821_),
    .A(\top_ihp.oisc.regs[44][31] ),
    .B(net355));
 sg13g2_o21ai_1 _17965_ (.B1(_10821_),
    .Y(_01598_),
    .A1(net116),
    .A2(_10794_));
 sg13g2_nand2_1 _17966_ (.Y(_10822_),
    .A(\top_ihp.oisc.regs[44][3] ),
    .B(net355));
 sg13g2_o21ai_1 _17967_ (.B1(_10822_),
    .Y(_01599_),
    .A1(_10498_),
    .A2(net354));
 sg13g2_nand2_1 _17968_ (.Y(_10823_),
    .A(\top_ihp.oisc.regs[44][4] ),
    .B(net355));
 sg13g2_o21ai_1 _17969_ (.B1(_10823_),
    .Y(_01600_),
    .A1(net117),
    .A2(net354));
 sg13g2_nand2_1 _17970_ (.Y(_10824_),
    .A(\top_ihp.oisc.regs[44][5] ),
    .B(net355));
 sg13g2_o21ai_1 _17971_ (.B1(_10824_),
    .Y(_01601_),
    .A1(net123),
    .A2(net354));
 sg13g2_nand2_1 _17972_ (.Y(_10825_),
    .A(\top_ihp.oisc.regs[44][6] ),
    .B(net355));
 sg13g2_o21ai_1 _17973_ (.B1(_10825_),
    .Y(_01602_),
    .A1(_10452_),
    .A2(net354));
 sg13g2_nand2_1 _17974_ (.Y(_10826_),
    .A(\top_ihp.oisc.regs[44][7] ),
    .B(_10792_));
 sg13g2_o21ai_1 _17975_ (.B1(_10826_),
    .Y(_01603_),
    .A1(_10189_),
    .A2(_10794_));
 sg13g2_nand2_1 _17976_ (.Y(_10827_),
    .A(\top_ihp.oisc.regs[44][8] ),
    .B(_10792_));
 sg13g2_o21ai_1 _17977_ (.B1(_10827_),
    .Y(_01604_),
    .A1(_10455_),
    .A2(net354));
 sg13g2_nand2_1 _17978_ (.Y(_10828_),
    .A(\top_ihp.oisc.regs[44][9] ),
    .B(net355));
 sg13g2_o21ai_1 _17979_ (.B1(_10828_),
    .Y(_01605_),
    .A1(net35),
    .A2(net354));
 sg13g2_nor2_1 _17980_ (.A(_10090_),
    .B(_10276_),
    .Y(_10829_));
 sg13g2_buf_1 _17981_ (.A(_10829_),
    .X(_10830_));
 sg13g2_mux2_1 _17982_ (.A0(\top_ihp.oisc.regs[45][0] ),
    .A1(net204),
    .S(_10830_),
    .X(_01606_));
 sg13g2_buf_8 _17983_ (.A(_10063_),
    .X(_10831_));
 sg13g2_nand3_1 _17984_ (.B(_10092_),
    .C(_10274_),
    .A(net665),
    .Y(_10832_));
 sg13g2_buf_2 _17985_ (.A(_10832_),
    .X(_10833_));
 sg13g2_buf_2 _17986_ (.A(_10833_),
    .X(_10834_));
 sg13g2_buf_1 _17987_ (.A(_10833_),
    .X(_10835_));
 sg13g2_nand2_1 _17988_ (.Y(_10836_),
    .A(\top_ihp.oisc.regs[45][10] ),
    .B(net350));
 sg13g2_o21ai_1 _17989_ (.B1(_10836_),
    .Y(_01607_),
    .A1(net33),
    .A2(net351));
 sg13g2_nand2_1 _17990_ (.Y(_10837_),
    .A(\top_ihp.oisc.regs[45][11] ),
    .B(net350));
 sg13g2_o21ai_1 _17991_ (.B1(_10837_),
    .Y(_01608_),
    .A1(net121),
    .A2(net351));
 sg13g2_buf_1 _17992_ (.A(_10064_),
    .X(_10838_));
 sg13g2_nand2_1 _17993_ (.Y(_10839_),
    .A(\top_ihp.oisc.regs[45][12] ),
    .B(net350));
 sg13g2_o21ai_1 _17994_ (.B1(_10839_),
    .Y(_01609_),
    .A1(net109),
    .A2(net351));
 sg13g2_nor2_1 _17995_ (.A(\top_ihp.oisc.regs[45][13] ),
    .B(net518),
    .Y(_10840_));
 sg13g2_a21oi_1 _17996_ (.A1(net59),
    .A2(net518),
    .Y(_01610_),
    .B1(_10840_));
 sg13g2_buf_1 _17997_ (.A(net217),
    .X(_10841_));
 sg13g2_nand2_1 _17998_ (.Y(_10842_),
    .A(\top_ihp.oisc.regs[45][14] ),
    .B(net350));
 sg13g2_o21ai_1 _17999_ (.B1(_10842_),
    .Y(_01611_),
    .A1(net108),
    .A2(net351));
 sg13g2_buf_1 _18000_ (.A(_10833_),
    .X(_10843_));
 sg13g2_nand2_1 _18001_ (.Y(_10844_),
    .A(\top_ihp.oisc.regs[45][15] ),
    .B(net349));
 sg13g2_o21ai_1 _18002_ (.B1(_10844_),
    .Y(_01612_),
    .A1(net120),
    .A2(net351));
 sg13g2_nor2_1 _18003_ (.A(\top_ihp.oisc.regs[45][16] ),
    .B(net518),
    .Y(_10845_));
 sg13g2_a21oi_1 _18004_ (.A1(net132),
    .A2(net518),
    .Y(_01613_),
    .B1(_10845_));
 sg13g2_buf_1 _18005_ (.A(_10070_),
    .X(_10846_));
 sg13g2_nand2_1 _18006_ (.Y(_10847_),
    .A(\top_ihp.oisc.regs[45][17] ),
    .B(net349));
 sg13g2_o21ai_1 _18007_ (.B1(_10847_),
    .Y(_01614_),
    .A1(net52),
    .A2(net351));
 sg13g2_buf_1 _18008_ (.A(_10071_),
    .X(_10848_));
 sg13g2_nand2_1 _18009_ (.Y(_10849_),
    .A(\top_ihp.oisc.regs[45][18] ),
    .B(net349));
 sg13g2_o21ai_1 _18010_ (.B1(_10849_),
    .Y(_01615_),
    .A1(net51),
    .A2(net351));
 sg13g2_buf_1 _18011_ (.A(net215),
    .X(_10850_));
 sg13g2_nand2_1 _18012_ (.Y(_10851_),
    .A(\top_ihp.oisc.regs[45][19] ),
    .B(net349));
 sg13g2_o21ai_1 _18013_ (.B1(_10851_),
    .Y(_01616_),
    .A1(net107),
    .A2(_10834_));
 sg13g2_buf_1 _18014_ (.A(_09552_),
    .X(_10852_));
 sg13g2_nand2_1 _18015_ (.Y(_10853_),
    .A(\top_ihp.oisc.regs[45][1] ),
    .B(net349));
 sg13g2_o21ai_1 _18016_ (.B1(_10853_),
    .Y(_01617_),
    .A1(net517),
    .A2(net351));
 sg13g2_nor2_1 _18017_ (.A(\top_ihp.oisc.regs[45][20] ),
    .B(net518),
    .Y(_10854_));
 sg13g2_a21oi_1 _18018_ (.A1(_09981_),
    .A2(net518),
    .Y(_01618_),
    .B1(_10854_));
 sg13g2_buf_8 _18019_ (.A(net64),
    .X(_10855_));
 sg13g2_nand2_1 _18020_ (.Y(_10856_),
    .A(\top_ihp.oisc.regs[45][21] ),
    .B(net349));
 sg13g2_o21ai_1 _18021_ (.B1(_10856_),
    .Y(_01619_),
    .A1(net32),
    .A2(_10834_));
 sg13g2_nor2_1 _18022_ (.A(\top_ihp.oisc.regs[45][22] ),
    .B(_10830_),
    .Y(_10857_));
 sg13g2_a21oi_1 _18023_ (.A1(net131),
    .A2(net518),
    .Y(_01620_),
    .B1(_10857_));
 sg13g2_nor2_1 _18024_ (.A(\top_ihp.oisc.regs[45][23] ),
    .B(_10829_),
    .Y(_10858_));
 sg13g2_a21oi_1 _18025_ (.A1(net138),
    .A2(net518),
    .Y(_01621_),
    .B1(_10858_));
 sg13g2_buf_1 _18026_ (.A(net214),
    .X(_10859_));
 sg13g2_buf_2 _18027_ (.A(_10833_),
    .X(_10860_));
 sg13g2_nand2_1 _18028_ (.Y(_10861_),
    .A(\top_ihp.oisc.regs[45][24] ),
    .B(_10843_));
 sg13g2_o21ai_1 _18029_ (.B1(_10861_),
    .Y(_01622_),
    .A1(net106),
    .A2(net348));
 sg13g2_buf_2 _18030_ (.A(net213),
    .X(_10862_));
 sg13g2_nand2_1 _18031_ (.Y(_10863_),
    .A(\top_ihp.oisc.regs[45][25] ),
    .B(net349));
 sg13g2_o21ai_1 _18032_ (.B1(_10863_),
    .Y(_01623_),
    .A1(net105),
    .A2(net348));
 sg13g2_buf_8 _18033_ (.A(net134),
    .X(_02648_));
 sg13g2_nand2_1 _18034_ (.Y(_02649_),
    .A(\top_ihp.oisc.regs[45][26] ),
    .B(_10843_));
 sg13g2_o21ai_1 _18035_ (.B1(_02649_),
    .Y(_01624_),
    .A1(net50),
    .A2(net348));
 sg13g2_buf_8 _18036_ (.A(net141),
    .X(_02650_));
 sg13g2_nand2_1 _18037_ (.Y(_02651_),
    .A(\top_ihp.oisc.regs[45][27] ),
    .B(net349));
 sg13g2_o21ai_1 _18038_ (.B1(_02651_),
    .Y(_01625_),
    .A1(net49),
    .A2(net348));
 sg13g2_buf_8 _18039_ (.A(net63),
    .X(_02652_));
 sg13g2_buf_1 _18040_ (.A(_10833_),
    .X(_02653_));
 sg13g2_nand2_1 _18041_ (.Y(_02654_),
    .A(\top_ihp.oisc.regs[45][28] ),
    .B(net347));
 sg13g2_o21ai_1 _18042_ (.B1(_02654_),
    .Y(_01626_),
    .A1(net31),
    .A2(_10860_));
 sg13g2_buf_2 _18043_ (.A(net133),
    .X(_02655_));
 sg13g2_nand2_1 _18044_ (.Y(_02656_),
    .A(\top_ihp.oisc.regs[45][29] ),
    .B(net347));
 sg13g2_o21ai_1 _18045_ (.B1(_02656_),
    .Y(_01627_),
    .A1(net48),
    .A2(net348));
 sg13g2_nand2_1 _18046_ (.Y(_02657_),
    .A(\top_ihp.oisc.regs[45][2] ),
    .B(net347));
 sg13g2_o21ai_1 _18047_ (.B1(_02657_),
    .Y(_01628_),
    .A1(_10493_),
    .A2(_10860_));
 sg13g2_nand2_1 _18048_ (.Y(_02658_),
    .A(\top_ihp.oisc.regs[45][30] ),
    .B(net347));
 sg13g2_o21ai_1 _18049_ (.B1(_02658_),
    .Y(_01629_),
    .A1(_10495_),
    .A2(net348));
 sg13g2_nand2_1 _18050_ (.Y(_02659_),
    .A(\top_ihp.oisc.regs[45][31] ),
    .B(net347));
 sg13g2_o21ai_1 _18051_ (.B1(_02659_),
    .Y(_01630_),
    .A1(net116),
    .A2(net348));
 sg13g2_nand2_1 _18052_ (.Y(_02660_),
    .A(\top_ihp.oisc.regs[45][3] ),
    .B(net347));
 sg13g2_o21ai_1 _18053_ (.B1(_02660_),
    .Y(_01631_),
    .A1(net118),
    .A2(net348));
 sg13g2_nand2_1 _18054_ (.Y(_02661_),
    .A(\top_ihp.oisc.regs[45][4] ),
    .B(net347));
 sg13g2_o21ai_1 _18055_ (.B1(_02661_),
    .Y(_01632_),
    .A1(net117),
    .A2(net350));
 sg13g2_buf_2 _18056_ (.A(_10085_),
    .X(_02662_));
 sg13g2_nand2_1 _18057_ (.Y(_02663_),
    .A(\top_ihp.oisc.regs[45][5] ),
    .B(net347));
 sg13g2_o21ai_1 _18058_ (.B1(_02663_),
    .Y(_01633_),
    .A1(net104),
    .A2(net350));
 sg13g2_buf_1 _18059_ (.A(net211),
    .X(_02664_));
 sg13g2_nand2_1 _18060_ (.Y(_02665_),
    .A(\top_ihp.oisc.regs[45][6] ),
    .B(_02653_));
 sg13g2_o21ai_1 _18061_ (.B1(_02665_),
    .Y(_01634_),
    .A1(net103),
    .A2(net350));
 sg13g2_buf_2 _18062_ (.A(net408),
    .X(_02666_));
 sg13g2_nand2_1 _18063_ (.Y(_02667_),
    .A(\top_ihp.oisc.regs[45][7] ),
    .B(_02653_));
 sg13g2_o21ai_1 _18064_ (.B1(_02667_),
    .Y(_01635_),
    .A1(net187),
    .A2(net350));
 sg13g2_buf_1 _18065_ (.A(net61),
    .X(_02668_));
 sg13g2_nand2_1 _18066_ (.Y(_02669_),
    .A(\top_ihp.oisc.regs[45][8] ),
    .B(_10833_));
 sg13g2_o21ai_1 _18067_ (.B1(_02669_),
    .Y(_01636_),
    .A1(net30),
    .A2(_10835_));
 sg13g2_buf_8 _18068_ (.A(net60),
    .X(_02670_));
 sg13g2_nand2_1 _18069_ (.Y(_02671_),
    .A(\top_ihp.oisc.regs[45][9] ),
    .B(_10833_));
 sg13g2_o21ai_1 _18070_ (.B1(_02671_),
    .Y(_01637_),
    .A1(net29),
    .A2(_10835_));
 sg13g2_and2_1 _18071_ (.A(net665),
    .B(net664),
    .X(_02672_));
 sg13g2_buf_1 _18072_ (.A(_02672_),
    .X(_02673_));
 sg13g2_buf_1 _18073_ (.A(_02673_),
    .X(_02674_));
 sg13g2_mux2_1 _18074_ (.A0(\top_ihp.oisc.regs[46][0] ),
    .A1(_10549_),
    .S(net346),
    .X(_01638_));
 sg13g2_nand2_1 _18075_ (.Y(_02675_),
    .A(net665),
    .B(net664));
 sg13g2_buf_2 _18076_ (.A(_02675_),
    .X(_02676_));
 sg13g2_buf_2 _18077_ (.A(_02676_),
    .X(_02677_));
 sg13g2_buf_1 _18078_ (.A(_02676_),
    .X(_02678_));
 sg13g2_nand2_1 _18079_ (.Y(_02679_),
    .A(\top_ihp.oisc.regs[46][10] ),
    .B(net344));
 sg13g2_o21ai_1 _18080_ (.B1(_02679_),
    .Y(_01639_),
    .A1(net33),
    .A2(net345));
 sg13g2_buf_1 _18081_ (.A(net251),
    .X(_02680_));
 sg13g2_nand2_1 _18082_ (.Y(_02681_),
    .A(\top_ihp.oisc.regs[46][11] ),
    .B(net344));
 sg13g2_o21ai_1 _18083_ (.B1(_02681_),
    .Y(_01640_),
    .A1(net102),
    .A2(net345));
 sg13g2_nand2_1 _18084_ (.Y(_02682_),
    .A(\top_ihp.oisc.regs[46][12] ),
    .B(net344));
 sg13g2_o21ai_1 _18085_ (.B1(_02682_),
    .Y(_01641_),
    .A1(net109),
    .A2(net345));
 sg13g2_nor2_1 _18086_ (.A(\top_ihp.oisc.regs[46][13] ),
    .B(net346),
    .Y(_02683_));
 sg13g2_a21oi_1 _18087_ (.A1(net59),
    .A2(net346),
    .Y(_01642_),
    .B1(_02683_));
 sg13g2_nand2_1 _18088_ (.Y(_02684_),
    .A(\top_ihp.oisc.regs[46][14] ),
    .B(net344));
 sg13g2_o21ai_1 _18089_ (.B1(_02684_),
    .Y(_01643_),
    .A1(net108),
    .A2(net345));
 sg13g2_buf_1 _18090_ (.A(_10068_),
    .X(_02685_));
 sg13g2_buf_1 _18091_ (.A(_02676_),
    .X(_02686_));
 sg13g2_nand2_1 _18092_ (.Y(_02687_),
    .A(\top_ihp.oisc.regs[46][15] ),
    .B(net343));
 sg13g2_o21ai_1 _18093_ (.B1(_02687_),
    .Y(_01644_),
    .A1(net101),
    .A2(net345));
 sg13g2_nor2_1 _18094_ (.A(\top_ihp.oisc.regs[46][16] ),
    .B(net346),
    .Y(_02688_));
 sg13g2_a21oi_1 _18095_ (.A1(net132),
    .A2(net346),
    .Y(_01645_),
    .B1(_02688_));
 sg13g2_nand2_1 _18096_ (.Y(_02689_),
    .A(\top_ihp.oisc.regs[46][17] ),
    .B(net343));
 sg13g2_o21ai_1 _18097_ (.B1(_02689_),
    .Y(_01646_),
    .A1(net52),
    .A2(net345));
 sg13g2_nand2_1 _18098_ (.Y(_02690_),
    .A(\top_ihp.oisc.regs[46][18] ),
    .B(net343));
 sg13g2_o21ai_1 _18099_ (.B1(_02690_),
    .Y(_01647_),
    .A1(net51),
    .A2(_02677_));
 sg13g2_nand2_1 _18100_ (.Y(_02691_),
    .A(\top_ihp.oisc.regs[46][19] ),
    .B(net343));
 sg13g2_o21ai_1 _18101_ (.B1(_02691_),
    .Y(_01648_),
    .A1(net107),
    .A2(net345));
 sg13g2_nand2_1 _18102_ (.Y(_02692_),
    .A(\top_ihp.oisc.regs[46][1] ),
    .B(_02686_));
 sg13g2_o21ai_1 _18103_ (.B1(_02692_),
    .Y(_01649_),
    .A1(net517),
    .A2(net345));
 sg13g2_buf_8 _18104_ (.A(_09581_),
    .X(_02693_));
 sg13g2_nor2_1 _18105_ (.A(\top_ihp.oisc.regs[46][20] ),
    .B(net346),
    .Y(_02694_));
 sg13g2_a21oi_1 _18106_ (.A1(net28),
    .A2(net346),
    .Y(_01650_),
    .B1(_02694_));
 sg13g2_nand2_1 _18107_ (.Y(_02695_),
    .A(\top_ihp.oisc.regs[46][21] ),
    .B(net343));
 sg13g2_o21ai_1 _18108_ (.B1(_02695_),
    .Y(_01651_),
    .A1(_10855_),
    .A2(_02677_));
 sg13g2_nor2_1 _18109_ (.A(\top_ihp.oisc.regs[46][22] ),
    .B(net346),
    .Y(_02696_));
 sg13g2_a21oi_1 _18110_ (.A1(net131),
    .A2(_02674_),
    .Y(_01652_),
    .B1(_02696_));
 sg13g2_buf_1 _18111_ (.A(net243),
    .X(_02697_));
 sg13g2_nor2_1 _18112_ (.A(\top_ihp.oisc.regs[46][23] ),
    .B(_02673_),
    .Y(_02698_));
 sg13g2_a21oi_1 _18113_ (.A1(net100),
    .A2(_02674_),
    .Y(_01653_),
    .B1(_02698_));
 sg13g2_buf_1 _18114_ (.A(_02676_),
    .X(_02699_));
 sg13g2_nand2_1 _18115_ (.Y(_02700_),
    .A(\top_ihp.oisc.regs[46][24] ),
    .B(net343));
 sg13g2_o21ai_1 _18116_ (.B1(_02700_),
    .Y(_01654_),
    .A1(net106),
    .A2(net342));
 sg13g2_nand2_1 _18117_ (.Y(_02701_),
    .A(\top_ihp.oisc.regs[46][25] ),
    .B(net343));
 sg13g2_o21ai_1 _18118_ (.B1(_02701_),
    .Y(_01655_),
    .A1(net105),
    .A2(net342));
 sg13g2_nand2_1 _18119_ (.Y(_02702_),
    .A(\top_ihp.oisc.regs[46][26] ),
    .B(_02686_));
 sg13g2_o21ai_1 _18120_ (.B1(_02702_),
    .Y(_01656_),
    .A1(net50),
    .A2(net342));
 sg13g2_nand2_1 _18121_ (.Y(_02703_),
    .A(\top_ihp.oisc.regs[46][27] ),
    .B(net343));
 sg13g2_o21ai_1 _18122_ (.B1(_02703_),
    .Y(_01657_),
    .A1(net49),
    .A2(net342));
 sg13g2_buf_1 _18123_ (.A(_02676_),
    .X(_02704_));
 sg13g2_nand2_1 _18124_ (.Y(_02705_),
    .A(\top_ihp.oisc.regs[46][28] ),
    .B(net341));
 sg13g2_o21ai_1 _18125_ (.B1(_02705_),
    .Y(_01658_),
    .A1(net31),
    .A2(_02699_));
 sg13g2_nand2_1 _18126_ (.Y(_02706_),
    .A(\top_ihp.oisc.regs[46][29] ),
    .B(net341));
 sg13g2_o21ai_1 _18127_ (.B1(_02706_),
    .Y(_01659_),
    .A1(net48),
    .A2(_02699_));
 sg13g2_buf_2 _18128_ (.A(_10044_),
    .X(_02707_));
 sg13g2_nand2_1 _18129_ (.Y(_02708_),
    .A(\top_ihp.oisc.regs[46][2] ),
    .B(net341));
 sg13g2_o21ai_1 _18130_ (.B1(_02708_),
    .Y(_01660_),
    .A1(net99),
    .A2(net342));
 sg13g2_buf_1 _18131_ (.A(net62),
    .X(_02709_));
 sg13g2_nand2_1 _18132_ (.Y(_02710_),
    .A(\top_ihp.oisc.regs[46][30] ),
    .B(net341));
 sg13g2_o21ai_1 _18133_ (.B1(_02710_),
    .Y(_01661_),
    .A1(net27),
    .A2(net342));
 sg13g2_nand2_1 _18134_ (.Y(_02711_),
    .A(\top_ihp.oisc.regs[46][31] ),
    .B(_02704_));
 sg13g2_o21ai_1 _18135_ (.B1(_02711_),
    .Y(_01662_),
    .A1(net116),
    .A2(net342));
 sg13g2_buf_2 _18136_ (.A(net221),
    .X(_02712_));
 sg13g2_nand2_1 _18137_ (.Y(_02713_),
    .A(\top_ihp.oisc.regs[46][3] ),
    .B(_02704_));
 sg13g2_o21ai_1 _18138_ (.B1(_02713_),
    .Y(_01663_),
    .A1(net98),
    .A2(net342));
 sg13g2_buf_2 _18139_ (.A(net220),
    .X(_02714_));
 sg13g2_nand2_1 _18140_ (.Y(_02715_),
    .A(\top_ihp.oisc.regs[46][4] ),
    .B(net341));
 sg13g2_o21ai_1 _18141_ (.B1(_02715_),
    .Y(_01664_),
    .A1(net97),
    .A2(net344));
 sg13g2_nand2_1 _18142_ (.Y(_02716_),
    .A(\top_ihp.oisc.regs[46][5] ),
    .B(net341));
 sg13g2_o21ai_1 _18143_ (.B1(_02716_),
    .Y(_01665_),
    .A1(net104),
    .A2(net344));
 sg13g2_nand2_1 _18144_ (.Y(_02717_),
    .A(\top_ihp.oisc.regs[46][6] ),
    .B(net341));
 sg13g2_o21ai_1 _18145_ (.B1(_02717_),
    .Y(_01666_),
    .A1(net103),
    .A2(net344));
 sg13g2_buf_2 _18146_ (.A(_09913_),
    .X(_02718_));
 sg13g2_nand2_1 _18147_ (.Y(_02719_),
    .A(\top_ihp.oisc.regs[46][7] ),
    .B(net341));
 sg13g2_o21ai_1 _18148_ (.B1(_02719_),
    .Y(_01667_),
    .A1(net47),
    .A2(_02678_));
 sg13g2_nand2_1 _18149_ (.Y(_02720_),
    .A(\top_ihp.oisc.regs[46][8] ),
    .B(_02676_));
 sg13g2_o21ai_1 _18150_ (.B1(_02720_),
    .Y(_01668_),
    .A1(net30),
    .A2(net344));
 sg13g2_nand2_1 _18151_ (.Y(_02721_),
    .A(\top_ihp.oisc.regs[46][9] ),
    .B(_02676_));
 sg13g2_o21ai_1 _18152_ (.B1(_02721_),
    .Y(_01669_),
    .A1(_02670_),
    .A2(_02678_));
 sg13g2_and2_1 _18153_ (.A(_10151_),
    .B(_10358_),
    .X(_02722_));
 sg13g2_buf_1 _18154_ (.A(_02722_),
    .X(_02723_));
 sg13g2_mux2_1 _18155_ (.A0(\top_ihp.oisc.regs[47][0] ),
    .A1(net204),
    .S(_02723_),
    .X(_01670_));
 sg13g2_nand2_1 _18156_ (.Y(_02724_),
    .A(_10055_),
    .B(_10358_));
 sg13g2_buf_1 _18157_ (.A(_02724_),
    .X(_02725_));
 sg13g2_buf_2 _18158_ (.A(_02725_),
    .X(_02726_));
 sg13g2_buf_2 _18159_ (.A(net340),
    .X(_02727_));
 sg13g2_buf_1 _18160_ (.A(_02725_),
    .X(_02728_));
 sg13g2_nand2_1 _18161_ (.Y(_02729_),
    .A(\top_ihp.oisc.regs[47][10] ),
    .B(net339));
 sg13g2_o21ai_1 _18162_ (.B1(_02729_),
    .Y(_01671_),
    .A1(net33),
    .A2(net186));
 sg13g2_buf_1 _18163_ (.A(_02725_),
    .X(_02730_));
 sg13g2_nand2_1 _18164_ (.Y(_02731_),
    .A(\top_ihp.oisc.regs[47][11] ),
    .B(net338));
 sg13g2_o21ai_1 _18165_ (.B1(_02731_),
    .Y(_01672_),
    .A1(net102),
    .A2(net186));
 sg13g2_nand2_1 _18166_ (.Y(_02732_),
    .A(\top_ihp.oisc.regs[47][12] ),
    .B(net338));
 sg13g2_o21ai_1 _18167_ (.B1(_02732_),
    .Y(_01673_),
    .A1(net109),
    .A2(net186));
 sg13g2_nand2_1 _18168_ (.Y(_02733_),
    .A(\top_ihp.oisc.regs[47][13] ),
    .B(net338));
 sg13g2_o21ai_1 _18169_ (.B1(_02733_),
    .Y(_01674_),
    .A1(net111),
    .A2(_02727_));
 sg13g2_nand2_1 _18170_ (.Y(_02734_),
    .A(\top_ihp.oisc.regs[47][14] ),
    .B(net338));
 sg13g2_o21ai_1 _18171_ (.B1(_02734_),
    .Y(_01675_),
    .A1(net108),
    .A2(net186));
 sg13g2_nand2_1 _18172_ (.Y(_02735_),
    .A(\top_ihp.oisc.regs[47][15] ),
    .B(net338));
 sg13g2_o21ai_1 _18173_ (.B1(_02735_),
    .Y(_01676_),
    .A1(net101),
    .A2(net186));
 sg13g2_nand2_1 _18174_ (.Y(_02736_),
    .A(\top_ihp.oisc.regs[47][16] ),
    .B(net338));
 sg13g2_o21ai_1 _18175_ (.B1(_02736_),
    .Y(_01677_),
    .A1(net191),
    .A2(net186));
 sg13g2_nand2_1 _18176_ (.Y(_02737_),
    .A(\top_ihp.oisc.regs[47][17] ),
    .B(net338));
 sg13g2_o21ai_1 _18177_ (.B1(_02737_),
    .Y(_01678_),
    .A1(net52),
    .A2(net186));
 sg13g2_nand2_1 _18178_ (.Y(_02738_),
    .A(\top_ihp.oisc.regs[47][18] ),
    .B(net338));
 sg13g2_o21ai_1 _18179_ (.B1(_02738_),
    .Y(_01679_),
    .A1(net51),
    .A2(net186));
 sg13g2_nand2_1 _18180_ (.Y(_02739_),
    .A(\top_ihp.oisc.regs[47][19] ),
    .B(_02730_));
 sg13g2_o21ai_1 _18181_ (.B1(_02739_),
    .Y(_01680_),
    .A1(_10850_),
    .A2(_02727_));
 sg13g2_buf_1 _18182_ (.A(net340),
    .X(_02740_));
 sg13g2_nand2_1 _18183_ (.Y(_02741_),
    .A(\top_ihp.oisc.regs[47][1] ),
    .B(_02730_));
 sg13g2_o21ai_1 _18184_ (.B1(_02741_),
    .Y(_01681_),
    .A1(net517),
    .A2(net185));
 sg13g2_mux2_1 _18185_ (.A0(\top_ihp.oisc.regs[47][20] ),
    .A1(net245),
    .S(_02723_),
    .X(_01682_));
 sg13g2_buf_1 _18186_ (.A(_02725_),
    .X(_02742_));
 sg13g2_nand2_1 _18187_ (.Y(_02743_),
    .A(\top_ihp.oisc.regs[47][21] ),
    .B(net337));
 sg13g2_o21ai_1 _18188_ (.B1(_02743_),
    .Y(_01683_),
    .A1(net32),
    .A2(net185));
 sg13g2_nand2_1 _18189_ (.Y(_02744_),
    .A(\top_ihp.oisc.regs[47][22] ),
    .B(net337));
 sg13g2_o21ai_1 _18190_ (.B1(_02744_),
    .Y(_01684_),
    .A1(net110),
    .A2(net185));
 sg13g2_mux2_1 _18191_ (.A0(\top_ihp.oisc.regs[47][23] ),
    .A1(net406),
    .S(_02723_),
    .X(_01685_));
 sg13g2_nand2_1 _18192_ (.Y(_02745_),
    .A(\top_ihp.oisc.regs[47][24] ),
    .B(net337));
 sg13g2_o21ai_1 _18193_ (.B1(_02745_),
    .Y(_01686_),
    .A1(net106),
    .A2(net185));
 sg13g2_nand2_1 _18194_ (.Y(_02746_),
    .A(\top_ihp.oisc.regs[47][25] ),
    .B(net337));
 sg13g2_o21ai_1 _18195_ (.B1(_02746_),
    .Y(_01687_),
    .A1(net105),
    .A2(net185));
 sg13g2_nand2_1 _18196_ (.Y(_02747_),
    .A(\top_ihp.oisc.regs[47][26] ),
    .B(net337));
 sg13g2_o21ai_1 _18197_ (.B1(_02747_),
    .Y(_01688_),
    .A1(net50),
    .A2(net185));
 sg13g2_nand2_1 _18198_ (.Y(_02748_),
    .A(\top_ihp.oisc.regs[47][27] ),
    .B(net337));
 sg13g2_o21ai_1 _18199_ (.B1(_02748_),
    .Y(_01689_),
    .A1(net49),
    .A2(_02740_));
 sg13g2_nand2_1 _18200_ (.Y(_02749_),
    .A(\top_ihp.oisc.regs[47][28] ),
    .B(_02742_));
 sg13g2_o21ai_1 _18201_ (.B1(_02749_),
    .Y(_01690_),
    .A1(net31),
    .A2(_02740_));
 sg13g2_nand2_1 _18202_ (.Y(_02750_),
    .A(\top_ihp.oisc.regs[47][29] ),
    .B(net337));
 sg13g2_o21ai_1 _18203_ (.B1(_02750_),
    .Y(_01691_),
    .A1(net48),
    .A2(net185));
 sg13g2_nand2_1 _18204_ (.Y(_02751_),
    .A(\top_ihp.oisc.regs[47][2] ),
    .B(net337));
 sg13g2_o21ai_1 _18205_ (.B1(_02751_),
    .Y(_01692_),
    .A1(_02707_),
    .A2(net185));
 sg13g2_nand2_1 _18206_ (.Y(_02752_),
    .A(\top_ihp.oisc.regs[47][30] ),
    .B(_02742_));
 sg13g2_o21ai_1 _18207_ (.B1(_02752_),
    .Y(_01693_),
    .A1(net27),
    .A2(_02728_));
 sg13g2_buf_8 _18208_ (.A(net239),
    .X(_02753_));
 sg13g2_nand2_1 _18209_ (.Y(_02754_),
    .A(\top_ihp.oisc.regs[47][31] ),
    .B(net340));
 sg13g2_o21ai_1 _18210_ (.B1(_02754_),
    .Y(_01694_),
    .A1(net96),
    .A2(net339));
 sg13g2_nand2_1 _18211_ (.Y(_02755_),
    .A(\top_ihp.oisc.regs[47][3] ),
    .B(net340));
 sg13g2_o21ai_1 _18212_ (.B1(_02755_),
    .Y(_01695_),
    .A1(net98),
    .A2(net339));
 sg13g2_nand2_1 _18213_ (.Y(_02756_),
    .A(\top_ihp.oisc.regs[47][4] ),
    .B(net340));
 sg13g2_o21ai_1 _18214_ (.B1(_02756_),
    .Y(_01696_),
    .A1(net97),
    .A2(net339));
 sg13g2_nand2_1 _18215_ (.Y(_02757_),
    .A(\top_ihp.oisc.regs[47][5] ),
    .B(net340));
 sg13g2_o21ai_1 _18216_ (.B1(_02757_),
    .Y(_01697_),
    .A1(net104),
    .A2(net339));
 sg13g2_nand2_1 _18217_ (.Y(_02758_),
    .A(\top_ihp.oisc.regs[47][6] ),
    .B(net340));
 sg13g2_o21ai_1 _18218_ (.B1(_02758_),
    .Y(_01698_),
    .A1(net103),
    .A2(net339));
 sg13g2_nand2_1 _18219_ (.Y(_02759_),
    .A(\top_ihp.oisc.regs[47][7] ),
    .B(_02726_));
 sg13g2_o21ai_1 _18220_ (.B1(_02759_),
    .Y(_01699_),
    .A1(net187),
    .A2(net339));
 sg13g2_nand2_1 _18221_ (.Y(_02760_),
    .A(\top_ihp.oisc.regs[47][8] ),
    .B(_02726_));
 sg13g2_o21ai_1 _18222_ (.B1(_02760_),
    .Y(_01700_),
    .A1(net30),
    .A2(_02728_));
 sg13g2_nand2_1 _18223_ (.Y(_02761_),
    .A(\top_ihp.oisc.regs[47][9] ),
    .B(net340));
 sg13g2_o21ai_1 _18224_ (.B1(_02761_),
    .Y(_01701_),
    .A1(net29),
    .A2(net339));
 sg13g2_nor2b_1 _18225_ (.A(_09088_),
    .B_N(_09092_),
    .Y(_02762_));
 sg13g2_buf_4 _18226_ (.X(_02763_),
    .A(_02762_));
 sg13g2_and2_1 _18227_ (.A(_09104_),
    .B(_02763_),
    .X(_02764_));
 sg13g2_buf_2 _18228_ (.A(_02764_),
    .X(_02765_));
 sg13g2_nor2b_1 _18229_ (.A(_09082_),
    .B_N(_02765_),
    .Y(_02766_));
 sg13g2_buf_1 _18230_ (.A(_02766_),
    .X(_02767_));
 sg13g2_mux2_1 _18231_ (.A0(\top_ihp.oisc.regs[48][0] ),
    .A1(net204),
    .S(net632),
    .X(_01702_));
 sg13g2_nand2b_1 _18232_ (.Y(_02768_),
    .B(_02765_),
    .A_N(_09082_));
 sg13g2_buf_2 _18233_ (.A(_02768_),
    .X(_02769_));
 sg13g2_buf_2 _18234_ (.A(_02769_),
    .X(_02770_));
 sg13g2_buf_1 _18235_ (.A(_02769_),
    .X(_02771_));
 sg13g2_nand2_1 _18236_ (.Y(_02772_),
    .A(\top_ihp.oisc.regs[48][10] ),
    .B(net515));
 sg13g2_o21ai_1 _18237_ (.B1(_02772_),
    .Y(_01703_),
    .A1(net33),
    .A2(net516));
 sg13g2_nand2_1 _18238_ (.Y(_02773_),
    .A(\top_ihp.oisc.regs[48][11] ),
    .B(net515));
 sg13g2_o21ai_1 _18239_ (.B1(_02773_),
    .Y(_01704_),
    .A1(net102),
    .A2(net516));
 sg13g2_nand2_1 _18240_ (.Y(_02774_),
    .A(\top_ihp.oisc.regs[48][12] ),
    .B(net515));
 sg13g2_o21ai_1 _18241_ (.B1(_02774_),
    .Y(_01705_),
    .A1(net109),
    .A2(net516));
 sg13g2_nor2_1 _18242_ (.A(\top_ihp.oisc.regs[48][13] ),
    .B(net632),
    .Y(_02775_));
 sg13g2_a21oi_1 _18243_ (.A1(net59),
    .A2(net632),
    .Y(_01706_),
    .B1(_02775_));
 sg13g2_nand2_1 _18244_ (.Y(_02776_),
    .A(\top_ihp.oisc.regs[48][14] ),
    .B(net515));
 sg13g2_o21ai_1 _18245_ (.B1(_02776_),
    .Y(_01707_),
    .A1(net108),
    .A2(net516));
 sg13g2_buf_2 _18246_ (.A(_02769_),
    .X(_02777_));
 sg13g2_nand2_1 _18247_ (.Y(_02778_),
    .A(\top_ihp.oisc.regs[48][15] ),
    .B(net514));
 sg13g2_o21ai_1 _18248_ (.B1(_02778_),
    .Y(_01708_),
    .A1(net101),
    .A2(net516));
 sg13g2_nor2_1 _18249_ (.A(\top_ihp.oisc.regs[48][16] ),
    .B(net632),
    .Y(_02779_));
 sg13g2_a21oi_1 _18250_ (.A1(net132),
    .A2(net632),
    .Y(_01709_),
    .B1(_02779_));
 sg13g2_nand2_1 _18251_ (.Y(_02780_),
    .A(\top_ihp.oisc.regs[48][17] ),
    .B(net514));
 sg13g2_o21ai_1 _18252_ (.B1(_02780_),
    .Y(_01710_),
    .A1(net52),
    .A2(net516));
 sg13g2_nand2_1 _18253_ (.Y(_02781_),
    .A(\top_ihp.oisc.regs[48][18] ),
    .B(net514));
 sg13g2_o21ai_1 _18254_ (.B1(_02781_),
    .Y(_01711_),
    .A1(net51),
    .A2(_02770_));
 sg13g2_nand2_1 _18255_ (.Y(_02782_),
    .A(\top_ihp.oisc.regs[48][19] ),
    .B(net514));
 sg13g2_o21ai_1 _18256_ (.B1(_02782_),
    .Y(_01712_),
    .A1(net107),
    .A2(net516));
 sg13g2_nand2_1 _18257_ (.Y(_02783_),
    .A(\top_ihp.oisc.regs[48][1] ),
    .B(net514));
 sg13g2_o21ai_1 _18258_ (.B1(_02783_),
    .Y(_01713_),
    .A1(net517),
    .A2(_02770_));
 sg13g2_nor2_1 _18259_ (.A(\top_ihp.oisc.regs[48][20] ),
    .B(net632),
    .Y(_02784_));
 sg13g2_a21oi_1 _18260_ (.A1(net28),
    .A2(net632),
    .Y(_01714_),
    .B1(_02784_));
 sg13g2_nand2_1 _18261_ (.Y(_02785_),
    .A(\top_ihp.oisc.regs[48][21] ),
    .B(net514));
 sg13g2_o21ai_1 _18262_ (.B1(_02785_),
    .Y(_01715_),
    .A1(net32),
    .A2(net516));
 sg13g2_nor2_1 _18263_ (.A(\top_ihp.oisc.regs[48][22] ),
    .B(_02767_),
    .Y(_02786_));
 sg13g2_a21oi_1 _18264_ (.A1(net131),
    .A2(_02767_),
    .Y(_01716_),
    .B1(_02786_));
 sg13g2_nor2_1 _18265_ (.A(\top_ihp.oisc.regs[48][23] ),
    .B(_02766_),
    .Y(_02787_));
 sg13g2_a21oi_1 _18266_ (.A1(net100),
    .A2(net632),
    .Y(_01717_),
    .B1(_02787_));
 sg13g2_buf_1 _18267_ (.A(_02769_),
    .X(_02788_));
 sg13g2_nand2_1 _18268_ (.Y(_02789_),
    .A(\top_ihp.oisc.regs[48][24] ),
    .B(net514));
 sg13g2_o21ai_1 _18269_ (.B1(_02789_),
    .Y(_01718_),
    .A1(net106),
    .A2(net513));
 sg13g2_nand2_1 _18270_ (.Y(_02790_),
    .A(\top_ihp.oisc.regs[48][25] ),
    .B(net514));
 sg13g2_o21ai_1 _18271_ (.B1(_02790_),
    .Y(_01719_),
    .A1(net105),
    .A2(net513));
 sg13g2_nand2_1 _18272_ (.Y(_02791_),
    .A(\top_ihp.oisc.regs[48][26] ),
    .B(_02777_));
 sg13g2_o21ai_1 _18273_ (.B1(_02791_),
    .Y(_01720_),
    .A1(net50),
    .A2(net513));
 sg13g2_nand2_1 _18274_ (.Y(_02792_),
    .A(\top_ihp.oisc.regs[48][27] ),
    .B(_02777_));
 sg13g2_o21ai_1 _18275_ (.B1(_02792_),
    .Y(_01721_),
    .A1(net49),
    .A2(net513));
 sg13g2_buf_1 _18276_ (.A(_02769_),
    .X(_02793_));
 sg13g2_nand2_1 _18277_ (.Y(_02794_),
    .A(\top_ihp.oisc.regs[48][28] ),
    .B(net512));
 sg13g2_o21ai_1 _18278_ (.B1(_02794_),
    .Y(_01722_),
    .A1(net31),
    .A2(_02788_));
 sg13g2_nand2_1 _18279_ (.Y(_02795_),
    .A(\top_ihp.oisc.regs[48][29] ),
    .B(net512));
 sg13g2_o21ai_1 _18280_ (.B1(_02795_),
    .Y(_01723_),
    .A1(net48),
    .A2(_02788_));
 sg13g2_nand2_1 _18281_ (.Y(_02796_),
    .A(\top_ihp.oisc.regs[48][2] ),
    .B(_02793_));
 sg13g2_o21ai_1 _18282_ (.B1(_02796_),
    .Y(_01724_),
    .A1(net99),
    .A2(net513));
 sg13g2_nand2_1 _18283_ (.Y(_02797_),
    .A(\top_ihp.oisc.regs[48][30] ),
    .B(net512));
 sg13g2_o21ai_1 _18284_ (.B1(_02797_),
    .Y(_01725_),
    .A1(net27),
    .A2(net513));
 sg13g2_nand2_1 _18285_ (.Y(_02798_),
    .A(\top_ihp.oisc.regs[48][31] ),
    .B(net512));
 sg13g2_o21ai_1 _18286_ (.B1(_02798_),
    .Y(_01726_),
    .A1(net96),
    .A2(net513));
 sg13g2_nand2_1 _18287_ (.Y(_02799_),
    .A(\top_ihp.oisc.regs[48][3] ),
    .B(_02793_));
 sg13g2_o21ai_1 _18288_ (.B1(_02799_),
    .Y(_01727_),
    .A1(net98),
    .A2(net513));
 sg13g2_nand2_1 _18289_ (.Y(_02800_),
    .A(\top_ihp.oisc.regs[48][4] ),
    .B(net512));
 sg13g2_o21ai_1 _18290_ (.B1(_02800_),
    .Y(_01728_),
    .A1(net97),
    .A2(net515));
 sg13g2_nand2_1 _18291_ (.Y(_02801_),
    .A(\top_ihp.oisc.regs[48][5] ),
    .B(net512));
 sg13g2_o21ai_1 _18292_ (.B1(_02801_),
    .Y(_01729_),
    .A1(net104),
    .A2(net515));
 sg13g2_nand2_1 _18293_ (.Y(_02802_),
    .A(\top_ihp.oisc.regs[48][6] ),
    .B(net512));
 sg13g2_o21ai_1 _18294_ (.B1(_02802_),
    .Y(_01730_),
    .A1(net103),
    .A2(_02771_));
 sg13g2_nand2_1 _18295_ (.Y(_02803_),
    .A(\top_ihp.oisc.regs[48][7] ),
    .B(net512));
 sg13g2_o21ai_1 _18296_ (.B1(_02803_),
    .Y(_01731_),
    .A1(net187),
    .A2(_02771_));
 sg13g2_nand2_1 _18297_ (.Y(_02804_),
    .A(\top_ihp.oisc.regs[48][8] ),
    .B(_02769_));
 sg13g2_o21ai_1 _18298_ (.B1(_02804_),
    .Y(_01732_),
    .A1(_02668_),
    .A2(net515));
 sg13g2_nand2_1 _18299_ (.Y(_02805_),
    .A(\top_ihp.oisc.regs[48][9] ),
    .B(_02769_));
 sg13g2_o21ai_1 _18300_ (.B1(_02805_),
    .Y(_01733_),
    .A1(net29),
    .A2(net515));
 sg13g2_and2_1 _18301_ (.A(net710),
    .B(_02765_),
    .X(_02806_));
 sg13g2_buf_1 _18302_ (.A(_02806_),
    .X(_02807_));
 sg13g2_mux2_1 _18303_ (.A0(\top_ihp.oisc.regs[49][0] ),
    .A1(net204),
    .S(_02807_),
    .X(_01734_));
 sg13g2_nand2_1 _18304_ (.Y(_02808_),
    .A(net710),
    .B(_02765_));
 sg13g2_buf_1 _18305_ (.A(_02808_),
    .X(_02809_));
 sg13g2_buf_1 _18306_ (.A(_02809_),
    .X(_02810_));
 sg13g2_buf_2 _18307_ (.A(net511),
    .X(_02811_));
 sg13g2_buf_1 _18308_ (.A(_02809_),
    .X(_02812_));
 sg13g2_nand2_1 _18309_ (.Y(_02813_),
    .A(\top_ihp.oisc.regs[49][10] ),
    .B(net510));
 sg13g2_o21ai_1 _18310_ (.B1(_02813_),
    .Y(_01735_),
    .A1(net33),
    .A2(_02811_));
 sg13g2_buf_1 _18311_ (.A(_02809_),
    .X(_02814_));
 sg13g2_nand2_1 _18312_ (.Y(_02815_),
    .A(\top_ihp.oisc.regs[49][11] ),
    .B(net509));
 sg13g2_o21ai_1 _18313_ (.B1(_02815_),
    .Y(_01736_),
    .A1(net102),
    .A2(net336));
 sg13g2_nand2_1 _18314_ (.Y(_02816_),
    .A(\top_ihp.oisc.regs[49][12] ),
    .B(net509));
 sg13g2_o21ai_1 _18315_ (.B1(_02816_),
    .Y(_01737_),
    .A1(net109),
    .A2(net336));
 sg13g2_nand2_1 _18316_ (.Y(_02817_),
    .A(\top_ihp.oisc.regs[49][13] ),
    .B(net509));
 sg13g2_o21ai_1 _18317_ (.B1(_02817_),
    .Y(_01738_),
    .A1(net111),
    .A2(_02811_));
 sg13g2_nand2_1 _18318_ (.Y(_02818_),
    .A(\top_ihp.oisc.regs[49][14] ),
    .B(net509));
 sg13g2_o21ai_1 _18319_ (.B1(_02818_),
    .Y(_01739_),
    .A1(_10841_),
    .A2(net336));
 sg13g2_nand2_1 _18320_ (.Y(_02819_),
    .A(\top_ihp.oisc.regs[49][15] ),
    .B(net509));
 sg13g2_o21ai_1 _18321_ (.B1(_02819_),
    .Y(_01740_),
    .A1(net101),
    .A2(net336));
 sg13g2_nand2_1 _18322_ (.Y(_02820_),
    .A(\top_ihp.oisc.regs[49][16] ),
    .B(net509));
 sg13g2_o21ai_1 _18323_ (.B1(_02820_),
    .Y(_01741_),
    .A1(net191),
    .A2(net336));
 sg13g2_nand2_1 _18324_ (.Y(_02821_),
    .A(\top_ihp.oisc.regs[49][17] ),
    .B(net509));
 sg13g2_o21ai_1 _18325_ (.B1(_02821_),
    .Y(_01742_),
    .A1(_10846_),
    .A2(net336));
 sg13g2_nand2_1 _18326_ (.Y(_02822_),
    .A(\top_ihp.oisc.regs[49][18] ),
    .B(_02814_));
 sg13g2_o21ai_1 _18327_ (.B1(_02822_),
    .Y(_01743_),
    .A1(_10848_),
    .A2(net336));
 sg13g2_nand2_1 _18328_ (.Y(_02823_),
    .A(\top_ihp.oisc.regs[49][19] ),
    .B(_02814_));
 sg13g2_o21ai_1 _18329_ (.B1(_02823_),
    .Y(_01744_),
    .A1(net107),
    .A2(net336));
 sg13g2_buf_1 _18330_ (.A(_02810_),
    .X(_02824_));
 sg13g2_nand2_1 _18331_ (.Y(_02825_),
    .A(\top_ihp.oisc.regs[49][1] ),
    .B(net509));
 sg13g2_o21ai_1 _18332_ (.B1(_02825_),
    .Y(_01745_),
    .A1(net517),
    .A2(net335));
 sg13g2_mux2_1 _18333_ (.A0(\top_ihp.oisc.regs[49][20] ),
    .A1(net245),
    .S(_02807_),
    .X(_01746_));
 sg13g2_buf_1 _18334_ (.A(_02809_),
    .X(_02826_));
 sg13g2_nand2_1 _18335_ (.Y(_02827_),
    .A(\top_ihp.oisc.regs[49][21] ),
    .B(net508));
 sg13g2_o21ai_1 _18336_ (.B1(_02827_),
    .Y(_01747_),
    .A1(net32),
    .A2(net335));
 sg13g2_nand2_1 _18337_ (.Y(_02828_),
    .A(\top_ihp.oisc.regs[49][22] ),
    .B(net508));
 sg13g2_o21ai_1 _18338_ (.B1(_02828_),
    .Y(_01748_),
    .A1(net110),
    .A2(net335));
 sg13g2_mux2_1 _18339_ (.A0(\top_ihp.oisc.regs[49][23] ),
    .A1(net406),
    .S(_02807_),
    .X(_01749_));
 sg13g2_nand2_1 _18340_ (.Y(_02829_),
    .A(\top_ihp.oisc.regs[49][24] ),
    .B(net508));
 sg13g2_o21ai_1 _18341_ (.B1(_02829_),
    .Y(_01750_),
    .A1(net106),
    .A2(net335));
 sg13g2_nand2_1 _18342_ (.Y(_02830_),
    .A(\top_ihp.oisc.regs[49][25] ),
    .B(net508));
 sg13g2_o21ai_1 _18343_ (.B1(_02830_),
    .Y(_01751_),
    .A1(net105),
    .A2(net335));
 sg13g2_nand2_1 _18344_ (.Y(_02831_),
    .A(\top_ihp.oisc.regs[49][26] ),
    .B(net508));
 sg13g2_o21ai_1 _18345_ (.B1(_02831_),
    .Y(_01752_),
    .A1(net50),
    .A2(net335));
 sg13g2_nand2_1 _18346_ (.Y(_02832_),
    .A(\top_ihp.oisc.regs[49][27] ),
    .B(net508));
 sg13g2_o21ai_1 _18347_ (.B1(_02832_),
    .Y(_01753_),
    .A1(net49),
    .A2(net335));
 sg13g2_nand2_1 _18348_ (.Y(_02833_),
    .A(\top_ihp.oisc.regs[49][28] ),
    .B(_02826_));
 sg13g2_o21ai_1 _18349_ (.B1(_02833_),
    .Y(_01754_),
    .A1(net31),
    .A2(_02824_));
 sg13g2_nand2_1 _18350_ (.Y(_02834_),
    .A(\top_ihp.oisc.regs[49][29] ),
    .B(_02826_));
 sg13g2_o21ai_1 _18351_ (.B1(_02834_),
    .Y(_01755_),
    .A1(net48),
    .A2(_02824_));
 sg13g2_nand2_1 _18352_ (.Y(_02835_),
    .A(\top_ihp.oisc.regs[49][2] ),
    .B(net508));
 sg13g2_o21ai_1 _18353_ (.B1(_02835_),
    .Y(_01756_),
    .A1(net99),
    .A2(net335));
 sg13g2_nand2_1 _18354_ (.Y(_02836_),
    .A(\top_ihp.oisc.regs[49][30] ),
    .B(net508));
 sg13g2_o21ai_1 _18355_ (.B1(_02836_),
    .Y(_01757_),
    .A1(net27),
    .A2(_02812_));
 sg13g2_nand2_1 _18356_ (.Y(_02837_),
    .A(\top_ihp.oisc.regs[49][31] ),
    .B(net511));
 sg13g2_o21ai_1 _18357_ (.B1(_02837_),
    .Y(_01758_),
    .A1(net96),
    .A2(net510));
 sg13g2_nand2_1 _18358_ (.Y(_02838_),
    .A(\top_ihp.oisc.regs[49][3] ),
    .B(_02810_));
 sg13g2_o21ai_1 _18359_ (.B1(_02838_),
    .Y(_01759_),
    .A1(net98),
    .A2(_02812_));
 sg13g2_nand2_1 _18360_ (.Y(_02839_),
    .A(\top_ihp.oisc.regs[49][4] ),
    .B(net511));
 sg13g2_o21ai_1 _18361_ (.B1(_02839_),
    .Y(_01760_),
    .A1(net97),
    .A2(net510));
 sg13g2_nand2_1 _18362_ (.Y(_02840_),
    .A(\top_ihp.oisc.regs[49][5] ),
    .B(net511));
 sg13g2_o21ai_1 _18363_ (.B1(_02840_),
    .Y(_01761_),
    .A1(_02662_),
    .A2(net510));
 sg13g2_nand2_1 _18364_ (.Y(_02841_),
    .A(\top_ihp.oisc.regs[49][6] ),
    .B(net511));
 sg13g2_o21ai_1 _18365_ (.B1(_02841_),
    .Y(_01762_),
    .A1(net103),
    .A2(net510));
 sg13g2_nand2_1 _18366_ (.Y(_02842_),
    .A(\top_ihp.oisc.regs[49][7] ),
    .B(net511));
 sg13g2_o21ai_1 _18367_ (.B1(_02842_),
    .Y(_01763_),
    .A1(net187),
    .A2(net510));
 sg13g2_nand2_1 _18368_ (.Y(_02843_),
    .A(\top_ihp.oisc.regs[49][8] ),
    .B(net511));
 sg13g2_o21ai_1 _18369_ (.B1(_02843_),
    .Y(_01764_),
    .A1(net30),
    .A2(net510));
 sg13g2_nand2_1 _18370_ (.Y(_02844_),
    .A(\top_ihp.oisc.regs[49][9] ),
    .B(net511));
 sg13g2_o21ai_1 _18371_ (.B1(_02844_),
    .Y(_01765_),
    .A1(net29),
    .A2(net510));
 sg13g2_buf_1 _18372_ (.A(_09198_),
    .X(_02845_));
 sg13g2_and2_1 _18373_ (.A(_10057_),
    .B(net663),
    .X(_02846_));
 sg13g2_buf_1 _18374_ (.A(_02846_),
    .X(_02847_));
 sg13g2_mux2_1 _18375_ (.A0(\top_ihp.oisc.regs[4][0] ),
    .A1(net334),
    .S(_02847_),
    .X(_01766_));
 sg13g2_nand2_1 _18376_ (.Y(_02848_),
    .A(_10057_),
    .B(_10397_));
 sg13g2_buf_1 _18377_ (.A(_02848_),
    .X(_02849_));
 sg13g2_buf_1 _18378_ (.A(_02849_),
    .X(_02850_));
 sg13g2_buf_1 _18379_ (.A(net333),
    .X(_02851_));
 sg13g2_buf_1 _18380_ (.A(_02849_),
    .X(_02852_));
 sg13g2_nand2_1 _18381_ (.Y(_02853_),
    .A(\top_ihp.oisc.regs[4][10] ),
    .B(net332));
 sg13g2_o21ai_1 _18382_ (.B1(_02853_),
    .Y(_01767_),
    .A1(_10831_),
    .A2(net184));
 sg13g2_buf_1 _18383_ (.A(_02849_),
    .X(_02854_));
 sg13g2_nand2_1 _18384_ (.Y(_02855_),
    .A(\top_ihp.oisc.regs[4][11] ),
    .B(net331));
 sg13g2_o21ai_1 _18385_ (.B1(_02855_),
    .Y(_01768_),
    .A1(_02680_),
    .A2(net184));
 sg13g2_nand2_1 _18386_ (.Y(_02856_),
    .A(\top_ihp.oisc.regs[4][12] ),
    .B(net331));
 sg13g2_o21ai_1 _18387_ (.B1(_02856_),
    .Y(_01769_),
    .A1(net109),
    .A2(net184));
 sg13g2_nand2_1 _18388_ (.Y(_02857_),
    .A(\top_ihp.oisc.regs[4][13] ),
    .B(net331));
 sg13g2_o21ai_1 _18389_ (.B1(_02857_),
    .Y(_01770_),
    .A1(_10799_),
    .A2(net184));
 sg13g2_nand2_1 _18390_ (.Y(_02858_),
    .A(\top_ihp.oisc.regs[4][14] ),
    .B(net331));
 sg13g2_o21ai_1 _18391_ (.B1(_02858_),
    .Y(_01771_),
    .A1(net108),
    .A2(net184));
 sg13g2_nand2_1 _18392_ (.Y(_02859_),
    .A(\top_ihp.oisc.regs[4][15] ),
    .B(net331));
 sg13g2_o21ai_1 _18393_ (.B1(_02859_),
    .Y(_01772_),
    .A1(net101),
    .A2(net184));
 sg13g2_nand2_1 _18394_ (.Y(_02860_),
    .A(\top_ihp.oisc.regs[4][16] ),
    .B(net331));
 sg13g2_o21ai_1 _18395_ (.B1(_02860_),
    .Y(_01773_),
    .A1(net191),
    .A2(net184));
 sg13g2_nand2_1 _18396_ (.Y(_02861_),
    .A(\top_ihp.oisc.regs[4][17] ),
    .B(net331));
 sg13g2_o21ai_1 _18397_ (.B1(_02861_),
    .Y(_01774_),
    .A1(_10846_),
    .A2(net184));
 sg13g2_nand2_1 _18398_ (.Y(_02862_),
    .A(\top_ihp.oisc.regs[4][18] ),
    .B(_02854_));
 sg13g2_o21ai_1 _18399_ (.B1(_02862_),
    .Y(_01775_),
    .A1(net51),
    .A2(_02851_));
 sg13g2_nand2_1 _18400_ (.Y(_02863_),
    .A(\top_ihp.oisc.regs[4][19] ),
    .B(_02854_));
 sg13g2_o21ai_1 _18401_ (.B1(_02863_),
    .Y(_01776_),
    .A1(net107),
    .A2(_02851_));
 sg13g2_buf_1 _18402_ (.A(_02850_),
    .X(_02864_));
 sg13g2_nand2_1 _18403_ (.Y(_02865_),
    .A(\top_ihp.oisc.regs[4][1] ),
    .B(net331));
 sg13g2_o21ai_1 _18404_ (.B1(_02865_),
    .Y(_01777_),
    .A1(net517),
    .A2(net183));
 sg13g2_nor2_1 _18405_ (.A(\top_ihp.oisc.regs[4][20] ),
    .B(_02847_),
    .Y(_02866_));
 sg13g2_a21oi_1 _18406_ (.A1(_02693_),
    .A2(_02847_),
    .Y(_01778_),
    .B1(_02866_));
 sg13g2_buf_1 _18407_ (.A(_02849_),
    .X(_02867_));
 sg13g2_nand2_1 _18408_ (.Y(_02868_),
    .A(\top_ihp.oisc.regs[4][21] ),
    .B(net330));
 sg13g2_o21ai_1 _18409_ (.B1(_02868_),
    .Y(_01779_),
    .A1(net32),
    .A2(net183));
 sg13g2_nand2_1 _18410_ (.Y(_02869_),
    .A(\top_ihp.oisc.regs[4][22] ),
    .B(net330));
 sg13g2_o21ai_1 _18411_ (.B1(_02869_),
    .Y(_01780_),
    .A1(_10811_),
    .A2(net183));
 sg13g2_nor2_1 _18412_ (.A(\top_ihp.oisc.regs[4][23] ),
    .B(_02847_),
    .Y(_02870_));
 sg13g2_a21oi_1 _18413_ (.A1(net100),
    .A2(_02847_),
    .Y(_01781_),
    .B1(_02870_));
 sg13g2_nand2_1 _18414_ (.Y(_02871_),
    .A(\top_ihp.oisc.regs[4][24] ),
    .B(net330));
 sg13g2_o21ai_1 _18415_ (.B1(_02871_),
    .Y(_01782_),
    .A1(_10859_),
    .A2(net183));
 sg13g2_nand2_1 _18416_ (.Y(_02872_),
    .A(\top_ihp.oisc.regs[4][25] ),
    .B(_02867_));
 sg13g2_o21ai_1 _18417_ (.B1(_02872_),
    .Y(_01783_),
    .A1(net105),
    .A2(_02864_));
 sg13g2_nand2_1 _18418_ (.Y(_02873_),
    .A(\top_ihp.oisc.regs[4][26] ),
    .B(_02867_));
 sg13g2_o21ai_1 _18419_ (.B1(_02873_),
    .Y(_01784_),
    .A1(_02648_),
    .A2(net183));
 sg13g2_nand2_1 _18420_ (.Y(_02874_),
    .A(\top_ihp.oisc.regs[4][27] ),
    .B(net330));
 sg13g2_o21ai_1 _18421_ (.B1(_02874_),
    .Y(_01785_),
    .A1(net49),
    .A2(net183));
 sg13g2_nand2_1 _18422_ (.Y(_02875_),
    .A(\top_ihp.oisc.regs[4][28] ),
    .B(net330));
 sg13g2_o21ai_1 _18423_ (.B1(_02875_),
    .Y(_01786_),
    .A1(_02652_),
    .A2(net183));
 sg13g2_nand2_1 _18424_ (.Y(_02876_),
    .A(\top_ihp.oisc.regs[4][29] ),
    .B(net330));
 sg13g2_o21ai_1 _18425_ (.B1(_02876_),
    .Y(_01787_),
    .A1(net48),
    .A2(_02864_));
 sg13g2_nand2_1 _18426_ (.Y(_02877_),
    .A(\top_ihp.oisc.regs[4][2] ),
    .B(net330));
 sg13g2_o21ai_1 _18427_ (.B1(_02877_),
    .Y(_01788_),
    .A1(_02707_),
    .A2(net183));
 sg13g2_nand2_1 _18428_ (.Y(_02878_),
    .A(\top_ihp.oisc.regs[4][30] ),
    .B(net330));
 sg13g2_o21ai_1 _18429_ (.B1(_02878_),
    .Y(_01789_),
    .A1(_02709_),
    .A2(net332));
 sg13g2_nand2_1 _18430_ (.Y(_02879_),
    .A(\top_ihp.oisc.regs[4][31] ),
    .B(net333));
 sg13g2_o21ai_1 _18431_ (.B1(_02879_),
    .Y(_01790_),
    .A1(_02753_),
    .A2(net332));
 sg13g2_nand2_1 _18432_ (.Y(_02880_),
    .A(\top_ihp.oisc.regs[4][3] ),
    .B(net333));
 sg13g2_o21ai_1 _18433_ (.B1(_02880_),
    .Y(_01791_),
    .A1(_02712_),
    .A2(net332));
 sg13g2_nand2_1 _18434_ (.Y(_02881_),
    .A(\top_ihp.oisc.regs[4][4] ),
    .B(_02850_));
 sg13g2_o21ai_1 _18435_ (.B1(_02881_),
    .Y(_01792_),
    .A1(_02714_),
    .A2(_02852_));
 sg13g2_nand2_1 _18436_ (.Y(_02882_),
    .A(\top_ihp.oisc.regs[4][5] ),
    .B(net333));
 sg13g2_o21ai_1 _18437_ (.B1(_02882_),
    .Y(_01793_),
    .A1(_02662_),
    .A2(_02852_));
 sg13g2_nand2_1 _18438_ (.Y(_02883_),
    .A(\top_ihp.oisc.regs[4][6] ),
    .B(net333));
 sg13g2_o21ai_1 _18439_ (.B1(_02883_),
    .Y(_01794_),
    .A1(_02664_),
    .A2(net332));
 sg13g2_nand2_1 _18440_ (.Y(_02884_),
    .A(\top_ihp.oisc.regs[4][7] ),
    .B(net333));
 sg13g2_o21ai_1 _18441_ (.B1(_02884_),
    .Y(_01795_),
    .A1(net47),
    .A2(net332));
 sg13g2_nand2_1 _18442_ (.Y(_02885_),
    .A(\top_ihp.oisc.regs[4][8] ),
    .B(net333));
 sg13g2_o21ai_1 _18443_ (.B1(_02885_),
    .Y(_01796_),
    .A1(_02668_),
    .A2(net332));
 sg13g2_nand2_1 _18444_ (.Y(_02886_),
    .A(\top_ihp.oisc.regs[4][9] ),
    .B(net333));
 sg13g2_o21ai_1 _18445_ (.B1(_02886_),
    .Y(_01797_),
    .A1(_02670_),
    .A2(net332));
 sg13g2_and2_1 _18446_ (.A(net711),
    .B(_02765_),
    .X(_02887_));
 sg13g2_buf_1 _18447_ (.A(_02887_),
    .X(_02888_));
 sg13g2_mux2_1 _18448_ (.A0(\top_ihp.oisc.regs[50][0] ),
    .A1(net334),
    .S(_02888_),
    .X(_01798_));
 sg13g2_nand2_1 _18449_ (.Y(_02889_),
    .A(net711),
    .B(_02765_));
 sg13g2_buf_1 _18450_ (.A(_02889_),
    .X(_02890_));
 sg13g2_buf_1 _18451_ (.A(_02890_),
    .X(_02891_));
 sg13g2_buf_1 _18452_ (.A(net507),
    .X(_02892_));
 sg13g2_buf_1 _18453_ (.A(_02890_),
    .X(_02893_));
 sg13g2_nand2_1 _18454_ (.Y(_02894_),
    .A(\top_ihp.oisc.regs[50][10] ),
    .B(net506));
 sg13g2_o21ai_1 _18455_ (.B1(_02894_),
    .Y(_01799_),
    .A1(_10831_),
    .A2(_02892_));
 sg13g2_buf_1 _18456_ (.A(_02890_),
    .X(_02895_));
 sg13g2_nand2_1 _18457_ (.Y(_02896_),
    .A(\top_ihp.oisc.regs[50][11] ),
    .B(_02895_));
 sg13g2_o21ai_1 _18458_ (.B1(_02896_),
    .Y(_01800_),
    .A1(net102),
    .A2(_02892_));
 sg13g2_nand2_1 _18459_ (.Y(_02897_),
    .A(\top_ihp.oisc.regs[50][12] ),
    .B(net505));
 sg13g2_o21ai_1 _18460_ (.B1(_02897_),
    .Y(_01801_),
    .A1(net109),
    .A2(net329));
 sg13g2_nand2_1 _18461_ (.Y(_02898_),
    .A(\top_ihp.oisc.regs[50][13] ),
    .B(net505));
 sg13g2_o21ai_1 _18462_ (.B1(_02898_),
    .Y(_01802_),
    .A1(net111),
    .A2(net329));
 sg13g2_nand2_1 _18463_ (.Y(_02899_),
    .A(\top_ihp.oisc.regs[50][14] ),
    .B(_02895_));
 sg13g2_o21ai_1 _18464_ (.B1(_02899_),
    .Y(_01803_),
    .A1(net108),
    .A2(net329));
 sg13g2_nand2_1 _18465_ (.Y(_02900_),
    .A(\top_ihp.oisc.regs[50][15] ),
    .B(net505));
 sg13g2_o21ai_1 _18466_ (.B1(_02900_),
    .Y(_01804_),
    .A1(_02685_),
    .A2(net329));
 sg13g2_nand2_1 _18467_ (.Y(_02901_),
    .A(\top_ihp.oisc.regs[50][16] ),
    .B(net505));
 sg13g2_o21ai_1 _18468_ (.B1(_02901_),
    .Y(_01805_),
    .A1(net191),
    .A2(net329));
 sg13g2_nand2_1 _18469_ (.Y(_02902_),
    .A(\top_ihp.oisc.regs[50][17] ),
    .B(net505));
 sg13g2_o21ai_1 _18470_ (.B1(_02902_),
    .Y(_01806_),
    .A1(net52),
    .A2(net329));
 sg13g2_nand2_1 _18471_ (.Y(_02903_),
    .A(\top_ihp.oisc.regs[50][18] ),
    .B(net505));
 sg13g2_o21ai_1 _18472_ (.B1(_02903_),
    .Y(_01807_),
    .A1(net51),
    .A2(net329));
 sg13g2_nand2_1 _18473_ (.Y(_02904_),
    .A(\top_ihp.oisc.regs[50][19] ),
    .B(net505));
 sg13g2_o21ai_1 _18474_ (.B1(_02904_),
    .Y(_01808_),
    .A1(_10850_),
    .A2(net329));
 sg13g2_buf_1 _18475_ (.A(net507),
    .X(_02905_));
 sg13g2_nand2_1 _18476_ (.Y(_02906_),
    .A(\top_ihp.oisc.regs[50][1] ),
    .B(net505));
 sg13g2_o21ai_1 _18477_ (.B1(_02906_),
    .Y(_01809_),
    .A1(net517),
    .A2(net328));
 sg13g2_nor2_1 _18478_ (.A(\top_ihp.oisc.regs[50][20] ),
    .B(_02888_),
    .Y(_02907_));
 sg13g2_a21oi_1 _18479_ (.A1(net28),
    .A2(_02888_),
    .Y(_01810_),
    .B1(_02907_));
 sg13g2_buf_1 _18480_ (.A(_02890_),
    .X(_02908_));
 sg13g2_nand2_1 _18481_ (.Y(_02909_),
    .A(\top_ihp.oisc.regs[50][21] ),
    .B(net504));
 sg13g2_o21ai_1 _18482_ (.B1(_02909_),
    .Y(_01811_),
    .A1(net32),
    .A2(net328));
 sg13g2_nand2_1 _18483_ (.Y(_02910_),
    .A(\top_ihp.oisc.regs[50][22] ),
    .B(net504));
 sg13g2_o21ai_1 _18484_ (.B1(_02910_),
    .Y(_01812_),
    .A1(net110),
    .A2(net328));
 sg13g2_nor2_1 _18485_ (.A(\top_ihp.oisc.regs[50][23] ),
    .B(_02888_),
    .Y(_02911_));
 sg13g2_a21oi_1 _18486_ (.A1(net100),
    .A2(_02888_),
    .Y(_01813_),
    .B1(_02911_));
 sg13g2_nand2_1 _18487_ (.Y(_02912_),
    .A(\top_ihp.oisc.regs[50][24] ),
    .B(net504));
 sg13g2_o21ai_1 _18488_ (.B1(_02912_),
    .Y(_01814_),
    .A1(net106),
    .A2(net328));
 sg13g2_nand2_1 _18489_ (.Y(_02913_),
    .A(\top_ihp.oisc.regs[50][25] ),
    .B(net504));
 sg13g2_o21ai_1 _18490_ (.B1(_02913_),
    .Y(_01815_),
    .A1(net105),
    .A2(net328));
 sg13g2_nand2_1 _18491_ (.Y(_02914_),
    .A(\top_ihp.oisc.regs[50][26] ),
    .B(net504));
 sg13g2_o21ai_1 _18492_ (.B1(_02914_),
    .Y(_01816_),
    .A1(net50),
    .A2(net328));
 sg13g2_nand2_1 _18493_ (.Y(_02915_),
    .A(\top_ihp.oisc.regs[50][27] ),
    .B(net504));
 sg13g2_o21ai_1 _18494_ (.B1(_02915_),
    .Y(_01817_),
    .A1(net49),
    .A2(_02905_));
 sg13g2_nand2_1 _18495_ (.Y(_02916_),
    .A(\top_ihp.oisc.regs[50][28] ),
    .B(_02908_));
 sg13g2_o21ai_1 _18496_ (.B1(_02916_),
    .Y(_01818_),
    .A1(net31),
    .A2(net328));
 sg13g2_nand2_1 _18497_ (.Y(_02917_),
    .A(\top_ihp.oisc.regs[50][29] ),
    .B(net504));
 sg13g2_o21ai_1 _18498_ (.B1(_02917_),
    .Y(_01819_),
    .A1(net48),
    .A2(net328));
 sg13g2_nand2_1 _18499_ (.Y(_02918_),
    .A(\top_ihp.oisc.regs[50][2] ),
    .B(net504));
 sg13g2_o21ai_1 _18500_ (.B1(_02918_),
    .Y(_01820_),
    .A1(net99),
    .A2(_02905_));
 sg13g2_nand2_1 _18501_ (.Y(_02919_),
    .A(\top_ihp.oisc.regs[50][30] ),
    .B(_02908_));
 sg13g2_o21ai_1 _18502_ (.B1(_02919_),
    .Y(_01821_),
    .A1(net27),
    .A2(_02893_));
 sg13g2_nand2_1 _18503_ (.Y(_02920_),
    .A(\top_ihp.oisc.regs[50][31] ),
    .B(net507));
 sg13g2_o21ai_1 _18504_ (.B1(_02920_),
    .Y(_01822_),
    .A1(net96),
    .A2(_02893_));
 sg13g2_nand2_1 _18505_ (.Y(_02921_),
    .A(\top_ihp.oisc.regs[50][3] ),
    .B(net507));
 sg13g2_o21ai_1 _18506_ (.B1(_02921_),
    .Y(_01823_),
    .A1(_02712_),
    .A2(net506));
 sg13g2_nand2_1 _18507_ (.Y(_02922_),
    .A(\top_ihp.oisc.regs[50][4] ),
    .B(net507));
 sg13g2_o21ai_1 _18508_ (.B1(_02922_),
    .Y(_01824_),
    .A1(net97),
    .A2(net506));
 sg13g2_nand2_1 _18509_ (.Y(_02923_),
    .A(\top_ihp.oisc.regs[50][5] ),
    .B(net507));
 sg13g2_o21ai_1 _18510_ (.B1(_02923_),
    .Y(_01825_),
    .A1(net104),
    .A2(net506));
 sg13g2_nand2_1 _18511_ (.Y(_02924_),
    .A(\top_ihp.oisc.regs[50][6] ),
    .B(_02891_));
 sg13g2_o21ai_1 _18512_ (.B1(_02924_),
    .Y(_01826_),
    .A1(_02664_),
    .A2(net506));
 sg13g2_nand2_1 _18513_ (.Y(_02925_),
    .A(\top_ihp.oisc.regs[50][7] ),
    .B(_02891_));
 sg13g2_o21ai_1 _18514_ (.B1(_02925_),
    .Y(_01827_),
    .A1(net47),
    .A2(net506));
 sg13g2_nand2_1 _18515_ (.Y(_02926_),
    .A(\top_ihp.oisc.regs[50][8] ),
    .B(net507));
 sg13g2_o21ai_1 _18516_ (.B1(_02926_),
    .Y(_01828_),
    .A1(net30),
    .A2(net506));
 sg13g2_nand2_1 _18517_ (.Y(_02927_),
    .A(\top_ihp.oisc.regs[50][9] ),
    .B(net507));
 sg13g2_o21ai_1 _18518_ (.B1(_02927_),
    .Y(_01829_),
    .A1(net29),
    .A2(net506));
 sg13g2_and2_1 _18519_ (.A(_10009_),
    .B(_02765_),
    .X(_02928_));
 sg13g2_buf_1 _18520_ (.A(_02928_),
    .X(_02929_));
 sg13g2_mux2_1 _18521_ (.A0(\top_ihp.oisc.regs[51][0] ),
    .A1(net334),
    .S(_02929_),
    .X(_01830_));
 sg13g2_nand2_1 _18522_ (.Y(_02930_),
    .A(_10009_),
    .B(_02765_));
 sg13g2_buf_1 _18523_ (.A(_02930_),
    .X(_02931_));
 sg13g2_buf_1 _18524_ (.A(_02931_),
    .X(_02932_));
 sg13g2_buf_2 _18525_ (.A(net503),
    .X(_02933_));
 sg13g2_buf_1 _18526_ (.A(_02931_),
    .X(_02934_));
 sg13g2_nand2_1 _18527_ (.Y(_02935_),
    .A(\top_ihp.oisc.regs[51][10] ),
    .B(net502));
 sg13g2_o21ai_1 _18528_ (.B1(_02935_),
    .Y(_01831_),
    .A1(net33),
    .A2(_02933_));
 sg13g2_buf_1 _18529_ (.A(_02931_),
    .X(_02936_));
 sg13g2_nand2_1 _18530_ (.Y(_02937_),
    .A(\top_ihp.oisc.regs[51][11] ),
    .B(net501));
 sg13g2_o21ai_1 _18531_ (.B1(_02937_),
    .Y(_01832_),
    .A1(net102),
    .A2(net327));
 sg13g2_nand2_1 _18532_ (.Y(_02938_),
    .A(\top_ihp.oisc.regs[51][12] ),
    .B(net501));
 sg13g2_o21ai_1 _18533_ (.B1(_02938_),
    .Y(_01833_),
    .A1(net109),
    .A2(net327));
 sg13g2_nand2_1 _18534_ (.Y(_02939_),
    .A(\top_ihp.oisc.regs[51][13] ),
    .B(net501));
 sg13g2_o21ai_1 _18535_ (.B1(_02939_),
    .Y(_01834_),
    .A1(net111),
    .A2(net327));
 sg13g2_nand2_1 _18536_ (.Y(_02940_),
    .A(\top_ihp.oisc.regs[51][14] ),
    .B(net501));
 sg13g2_o21ai_1 _18537_ (.B1(_02940_),
    .Y(_01835_),
    .A1(net108),
    .A2(net327));
 sg13g2_nand2_1 _18538_ (.Y(_02941_),
    .A(\top_ihp.oisc.regs[51][15] ),
    .B(net501));
 sg13g2_o21ai_1 _18539_ (.B1(_02941_),
    .Y(_01836_),
    .A1(net101),
    .A2(net327));
 sg13g2_nand2_1 _18540_ (.Y(_02942_),
    .A(\top_ihp.oisc.regs[51][16] ),
    .B(net501));
 sg13g2_o21ai_1 _18541_ (.B1(_02942_),
    .Y(_01837_),
    .A1(net191),
    .A2(net327));
 sg13g2_nand2_1 _18542_ (.Y(_02943_),
    .A(\top_ihp.oisc.regs[51][17] ),
    .B(net501));
 sg13g2_o21ai_1 _18543_ (.B1(_02943_),
    .Y(_01838_),
    .A1(net52),
    .A2(net327));
 sg13g2_nand2_1 _18544_ (.Y(_02944_),
    .A(\top_ihp.oisc.regs[51][18] ),
    .B(_02936_));
 sg13g2_o21ai_1 _18545_ (.B1(_02944_),
    .Y(_01839_),
    .A1(net51),
    .A2(net327));
 sg13g2_nand2_1 _18546_ (.Y(_02945_),
    .A(\top_ihp.oisc.regs[51][19] ),
    .B(_02936_));
 sg13g2_o21ai_1 _18547_ (.B1(_02945_),
    .Y(_01840_),
    .A1(net107),
    .A2(_02933_));
 sg13g2_buf_1 _18548_ (.A(_02932_),
    .X(_02946_));
 sg13g2_nand2_1 _18549_ (.Y(_02947_),
    .A(\top_ihp.oisc.regs[51][1] ),
    .B(net501));
 sg13g2_o21ai_1 _18550_ (.B1(_02947_),
    .Y(_01841_),
    .A1(_10852_),
    .A2(net326));
 sg13g2_mux2_1 _18551_ (.A0(\top_ihp.oisc.regs[51][20] ),
    .A1(net245),
    .S(_02929_),
    .X(_01842_));
 sg13g2_buf_1 _18552_ (.A(_02931_),
    .X(_02948_));
 sg13g2_nand2_1 _18553_ (.Y(_02949_),
    .A(\top_ihp.oisc.regs[51][21] ),
    .B(net500));
 sg13g2_o21ai_1 _18554_ (.B1(_02949_),
    .Y(_01843_),
    .A1(net32),
    .A2(net326));
 sg13g2_nand2_1 _18555_ (.Y(_02950_),
    .A(\top_ihp.oisc.regs[51][22] ),
    .B(net500));
 sg13g2_o21ai_1 _18556_ (.B1(_02950_),
    .Y(_01844_),
    .A1(net110),
    .A2(net326));
 sg13g2_mux2_1 _18557_ (.A0(\top_ihp.oisc.regs[51][23] ),
    .A1(net406),
    .S(_02929_),
    .X(_01845_));
 sg13g2_nand2_1 _18558_ (.Y(_02951_),
    .A(\top_ihp.oisc.regs[51][24] ),
    .B(net500));
 sg13g2_o21ai_1 _18559_ (.B1(_02951_),
    .Y(_01846_),
    .A1(net106),
    .A2(net326));
 sg13g2_nand2_1 _18560_ (.Y(_02952_),
    .A(\top_ihp.oisc.regs[51][25] ),
    .B(net500));
 sg13g2_o21ai_1 _18561_ (.B1(_02952_),
    .Y(_01847_),
    .A1(_10862_),
    .A2(net326));
 sg13g2_nand2_1 _18562_ (.Y(_02953_),
    .A(\top_ihp.oisc.regs[51][26] ),
    .B(net500));
 sg13g2_o21ai_1 _18563_ (.B1(_02953_),
    .Y(_01848_),
    .A1(net50),
    .A2(net326));
 sg13g2_nand2_1 _18564_ (.Y(_02954_),
    .A(\top_ihp.oisc.regs[51][27] ),
    .B(net500));
 sg13g2_o21ai_1 _18565_ (.B1(_02954_),
    .Y(_01849_),
    .A1(net49),
    .A2(net326));
 sg13g2_nand2_1 _18566_ (.Y(_02955_),
    .A(\top_ihp.oisc.regs[51][28] ),
    .B(net500));
 sg13g2_o21ai_1 _18567_ (.B1(_02955_),
    .Y(_01850_),
    .A1(net31),
    .A2(_02946_));
 sg13g2_nand2_1 _18568_ (.Y(_02956_),
    .A(\top_ihp.oisc.regs[51][29] ),
    .B(_02948_));
 sg13g2_o21ai_1 _18569_ (.B1(_02956_),
    .Y(_01851_),
    .A1(_02655_),
    .A2(_02946_));
 sg13g2_nand2_1 _18570_ (.Y(_02957_),
    .A(\top_ihp.oisc.regs[51][2] ),
    .B(net500));
 sg13g2_o21ai_1 _18571_ (.B1(_02957_),
    .Y(_01852_),
    .A1(net99),
    .A2(net326));
 sg13g2_nand2_1 _18572_ (.Y(_02958_),
    .A(\top_ihp.oisc.regs[51][30] ),
    .B(_02948_));
 sg13g2_o21ai_1 _18573_ (.B1(_02958_),
    .Y(_01853_),
    .A1(_02709_),
    .A2(net502));
 sg13g2_nand2_1 _18574_ (.Y(_02959_),
    .A(\top_ihp.oisc.regs[51][31] ),
    .B(net503));
 sg13g2_o21ai_1 _18575_ (.B1(_02959_),
    .Y(_01854_),
    .A1(net96),
    .A2(_02934_));
 sg13g2_nand2_1 _18576_ (.Y(_02960_),
    .A(\top_ihp.oisc.regs[51][3] ),
    .B(_02932_));
 sg13g2_o21ai_1 _18577_ (.B1(_02960_),
    .Y(_01855_),
    .A1(net98),
    .A2(_02934_));
 sg13g2_nand2_1 _18578_ (.Y(_02961_),
    .A(\top_ihp.oisc.regs[51][4] ),
    .B(net503));
 sg13g2_o21ai_1 _18579_ (.B1(_02961_),
    .Y(_01856_),
    .A1(net97),
    .A2(net502));
 sg13g2_nand2_1 _18580_ (.Y(_02962_),
    .A(\top_ihp.oisc.regs[51][5] ),
    .B(net503));
 sg13g2_o21ai_1 _18581_ (.B1(_02962_),
    .Y(_01857_),
    .A1(net104),
    .A2(net502));
 sg13g2_nand2_1 _18582_ (.Y(_02963_),
    .A(\top_ihp.oisc.regs[51][6] ),
    .B(net503));
 sg13g2_o21ai_1 _18583_ (.B1(_02963_),
    .Y(_01858_),
    .A1(net103),
    .A2(net502));
 sg13g2_nand2_1 _18584_ (.Y(_02964_),
    .A(\top_ihp.oisc.regs[51][7] ),
    .B(net503));
 sg13g2_o21ai_1 _18585_ (.B1(_02964_),
    .Y(_01859_),
    .A1(net187),
    .A2(net502));
 sg13g2_nand2_1 _18586_ (.Y(_02965_),
    .A(\top_ihp.oisc.regs[51][8] ),
    .B(net503));
 sg13g2_o21ai_1 _18587_ (.B1(_02965_),
    .Y(_01860_),
    .A1(net30),
    .A2(net502));
 sg13g2_nand2_1 _18588_ (.Y(_02966_),
    .A(\top_ihp.oisc.regs[51][9] ),
    .B(net503));
 sg13g2_o21ai_1 _18589_ (.B1(_02966_),
    .Y(_01861_),
    .A1(net29),
    .A2(net502));
 sg13g2_nor2b_1 _18590_ (.A(_09082_),
    .B_N(_02763_),
    .Y(_02967_));
 sg13g2_buf_2 _18591_ (.A(_02967_),
    .X(_02968_));
 sg13g2_and2_1 _18592_ (.A(_10398_),
    .B(_02968_),
    .X(_02969_));
 sg13g2_buf_1 _18593_ (.A(_02969_),
    .X(_02970_));
 sg13g2_mux2_1 _18594_ (.A0(\top_ihp.oisc.regs[52][0] ),
    .A1(net334),
    .S(_02970_),
    .X(_01862_));
 sg13g2_nand2_1 _18595_ (.Y(_02971_),
    .A(_10397_),
    .B(_02968_));
 sg13g2_buf_1 _18596_ (.A(_02971_),
    .X(_02972_));
 sg13g2_buf_1 _18597_ (.A(_02972_),
    .X(_02973_));
 sg13g2_buf_2 _18598_ (.A(net325),
    .X(_02974_));
 sg13g2_buf_1 _18599_ (.A(_02972_),
    .X(_02975_));
 sg13g2_nand2_1 _18600_ (.Y(_02976_),
    .A(\top_ihp.oisc.regs[52][10] ),
    .B(net324));
 sg13g2_o21ai_1 _18601_ (.B1(_02976_),
    .Y(_01863_),
    .A1(net33),
    .A2(_02974_));
 sg13g2_buf_1 _18602_ (.A(_02972_),
    .X(_02977_));
 sg13g2_nand2_1 _18603_ (.Y(_02978_),
    .A(\top_ihp.oisc.regs[52][11] ),
    .B(net323));
 sg13g2_o21ai_1 _18604_ (.B1(_02978_),
    .Y(_01864_),
    .A1(net102),
    .A2(net182));
 sg13g2_nand2_1 _18605_ (.Y(_02979_),
    .A(\top_ihp.oisc.regs[52][12] ),
    .B(net323));
 sg13g2_o21ai_1 _18606_ (.B1(_02979_),
    .Y(_01865_),
    .A1(_10838_),
    .A2(net182));
 sg13g2_nand2_1 _18607_ (.Y(_02980_),
    .A(\top_ihp.oisc.regs[52][13] ),
    .B(_02977_));
 sg13g2_o21ai_1 _18608_ (.B1(_02980_),
    .Y(_01866_),
    .A1(net111),
    .A2(net182));
 sg13g2_nand2_1 _18609_ (.Y(_02981_),
    .A(\top_ihp.oisc.regs[52][14] ),
    .B(net323));
 sg13g2_o21ai_1 _18610_ (.B1(_02981_),
    .Y(_01867_),
    .A1(net108),
    .A2(net182));
 sg13g2_nand2_1 _18611_ (.Y(_02982_),
    .A(\top_ihp.oisc.regs[52][15] ),
    .B(net323));
 sg13g2_o21ai_1 _18612_ (.B1(_02982_),
    .Y(_01868_),
    .A1(_02685_),
    .A2(net182));
 sg13g2_nand2_1 _18613_ (.Y(_02983_),
    .A(\top_ihp.oisc.regs[52][16] ),
    .B(net323));
 sg13g2_o21ai_1 _18614_ (.B1(_02983_),
    .Y(_01869_),
    .A1(_10762_),
    .A2(net182));
 sg13g2_nand2_1 _18615_ (.Y(_02984_),
    .A(\top_ihp.oisc.regs[52][17] ),
    .B(net323));
 sg13g2_o21ai_1 _18616_ (.B1(_02984_),
    .Y(_01870_),
    .A1(net52),
    .A2(net182));
 sg13g2_nand2_1 _18617_ (.Y(_02985_),
    .A(\top_ihp.oisc.regs[52][18] ),
    .B(net323));
 sg13g2_o21ai_1 _18618_ (.B1(_02985_),
    .Y(_01871_),
    .A1(net51),
    .A2(net182));
 sg13g2_nand2_1 _18619_ (.Y(_02986_),
    .A(\top_ihp.oisc.regs[52][19] ),
    .B(_02977_));
 sg13g2_o21ai_1 _18620_ (.B1(_02986_),
    .Y(_01872_),
    .A1(net107),
    .A2(_02974_));
 sg13g2_buf_1 _18621_ (.A(net325),
    .X(_02987_));
 sg13g2_nand2_1 _18622_ (.Y(_02988_),
    .A(\top_ihp.oisc.regs[52][1] ),
    .B(net323));
 sg13g2_o21ai_1 _18623_ (.B1(_02988_),
    .Y(_01873_),
    .A1(net517),
    .A2(net181));
 sg13g2_mux2_1 _18624_ (.A0(\top_ihp.oisc.regs[52][20] ),
    .A1(net245),
    .S(_02970_),
    .X(_01874_));
 sg13g2_buf_1 _18625_ (.A(_02972_),
    .X(_02989_));
 sg13g2_nand2_1 _18626_ (.Y(_02990_),
    .A(\top_ihp.oisc.regs[52][21] ),
    .B(net322));
 sg13g2_o21ai_1 _18627_ (.B1(_02990_),
    .Y(_01875_),
    .A1(net32),
    .A2(net181));
 sg13g2_nand2_1 _18628_ (.Y(_02991_),
    .A(\top_ihp.oisc.regs[52][22] ),
    .B(net322));
 sg13g2_o21ai_1 _18629_ (.B1(_02991_),
    .Y(_01876_),
    .A1(net110),
    .A2(net181));
 sg13g2_mux2_1 _18630_ (.A0(\top_ihp.oisc.regs[52][23] ),
    .A1(net406),
    .S(_02970_),
    .X(_01877_));
 sg13g2_nand2_1 _18631_ (.Y(_02992_),
    .A(\top_ihp.oisc.regs[52][24] ),
    .B(net322));
 sg13g2_o21ai_1 _18632_ (.B1(_02992_),
    .Y(_01878_),
    .A1(_10859_),
    .A2(_02987_));
 sg13g2_nand2_1 _18633_ (.Y(_02993_),
    .A(\top_ihp.oisc.regs[52][25] ),
    .B(net322));
 sg13g2_o21ai_1 _18634_ (.B1(_02993_),
    .Y(_01879_),
    .A1(net105),
    .A2(net181));
 sg13g2_nand2_1 _18635_ (.Y(_02994_),
    .A(\top_ihp.oisc.regs[52][26] ),
    .B(net322));
 sg13g2_o21ai_1 _18636_ (.B1(_02994_),
    .Y(_01880_),
    .A1(net50),
    .A2(net181));
 sg13g2_nand2_1 _18637_ (.Y(_02995_),
    .A(\top_ihp.oisc.regs[52][27] ),
    .B(net322));
 sg13g2_o21ai_1 _18638_ (.B1(_02995_),
    .Y(_01881_),
    .A1(_02650_),
    .A2(_02987_));
 sg13g2_nand2_1 _18639_ (.Y(_02996_),
    .A(\top_ihp.oisc.regs[52][28] ),
    .B(_02989_));
 sg13g2_o21ai_1 _18640_ (.B1(_02996_),
    .Y(_01882_),
    .A1(net31),
    .A2(net181));
 sg13g2_nand2_1 _18641_ (.Y(_02997_),
    .A(\top_ihp.oisc.regs[52][29] ),
    .B(net322));
 sg13g2_o21ai_1 _18642_ (.B1(_02997_),
    .Y(_01883_),
    .A1(net48),
    .A2(net181));
 sg13g2_nand2_1 _18643_ (.Y(_02998_),
    .A(\top_ihp.oisc.regs[52][2] ),
    .B(net322));
 sg13g2_o21ai_1 _18644_ (.B1(_02998_),
    .Y(_01884_),
    .A1(net99),
    .A2(net181));
 sg13g2_nand2_1 _18645_ (.Y(_02999_),
    .A(\top_ihp.oisc.regs[52][30] ),
    .B(_02989_));
 sg13g2_o21ai_1 _18646_ (.B1(_02999_),
    .Y(_01885_),
    .A1(net27),
    .A2(_02975_));
 sg13g2_nand2_1 _18647_ (.Y(_03000_),
    .A(\top_ihp.oisc.regs[52][31] ),
    .B(_02973_));
 sg13g2_o21ai_1 _18648_ (.B1(_03000_),
    .Y(_01886_),
    .A1(net96),
    .A2(net324));
 sg13g2_nand2_1 _18649_ (.Y(_03001_),
    .A(\top_ihp.oisc.regs[52][3] ),
    .B(net325));
 sg13g2_o21ai_1 _18650_ (.B1(_03001_),
    .Y(_01887_),
    .A1(net98),
    .A2(net324));
 sg13g2_nand2_1 _18651_ (.Y(_03002_),
    .A(\top_ihp.oisc.regs[52][4] ),
    .B(net325));
 sg13g2_o21ai_1 _18652_ (.B1(_03002_),
    .Y(_01888_),
    .A1(_02714_),
    .A2(_02975_));
 sg13g2_nand2_1 _18653_ (.Y(_03003_),
    .A(\top_ihp.oisc.regs[52][5] ),
    .B(_02973_));
 sg13g2_o21ai_1 _18654_ (.B1(_03003_),
    .Y(_01889_),
    .A1(net104),
    .A2(net324));
 sg13g2_nand2_1 _18655_ (.Y(_03004_),
    .A(\top_ihp.oisc.regs[52][6] ),
    .B(net325));
 sg13g2_o21ai_1 _18656_ (.B1(_03004_),
    .Y(_01890_),
    .A1(net103),
    .A2(net324));
 sg13g2_nand2_1 _18657_ (.Y(_03005_),
    .A(\top_ihp.oisc.regs[52][7] ),
    .B(net325));
 sg13g2_o21ai_1 _18658_ (.B1(_03005_),
    .Y(_01891_),
    .A1(net187),
    .A2(net324));
 sg13g2_nand2_1 _18659_ (.Y(_03006_),
    .A(\top_ihp.oisc.regs[52][8] ),
    .B(net325));
 sg13g2_o21ai_1 _18660_ (.B1(_03006_),
    .Y(_01892_),
    .A1(net30),
    .A2(net324));
 sg13g2_nand2_1 _18661_ (.Y(_03007_),
    .A(\top_ihp.oisc.regs[52][9] ),
    .B(net325));
 sg13g2_o21ai_1 _18662_ (.B1(_03007_),
    .Y(_01893_),
    .A1(net29),
    .A2(net324));
 sg13g2_nand2_1 _18663_ (.Y(_03008_),
    .A(net710),
    .B(_02763_));
 sg13g2_buf_1 _18664_ (.A(_03008_),
    .X(_03009_));
 sg13g2_nor2_1 _18665_ (.A(net682),
    .B(_03009_),
    .Y(_03010_));
 sg13g2_buf_1 _18666_ (.A(_03010_),
    .X(_03011_));
 sg13g2_mux2_1 _18667_ (.A0(\top_ihp.oisc.regs[53][0] ),
    .A1(net334),
    .S(net499),
    .X(_01894_));
 sg13g2_or2_1 _18668_ (.X(_03012_),
    .B(_03009_),
    .A(net682));
 sg13g2_buf_2 _18669_ (.A(_03012_),
    .X(_03013_));
 sg13g2_buf_2 _18670_ (.A(_03013_),
    .X(_03014_));
 sg13g2_buf_1 _18671_ (.A(_03013_),
    .X(_03015_));
 sg13g2_nand2_1 _18672_ (.Y(_03016_),
    .A(\top_ihp.oisc.regs[53][10] ),
    .B(net320));
 sg13g2_o21ai_1 _18673_ (.B1(_03016_),
    .Y(_01895_),
    .A1(net33),
    .A2(net321));
 sg13g2_nand2_1 _18674_ (.Y(_03017_),
    .A(\top_ihp.oisc.regs[53][11] ),
    .B(net320));
 sg13g2_o21ai_1 _18675_ (.B1(_03017_),
    .Y(_01896_),
    .A1(net102),
    .A2(net321));
 sg13g2_nand2_1 _18676_ (.Y(_03018_),
    .A(\top_ihp.oisc.regs[53][12] ),
    .B(net320));
 sg13g2_o21ai_1 _18677_ (.B1(_03018_),
    .Y(_01897_),
    .A1(_10838_),
    .A2(net321));
 sg13g2_nor2_1 _18678_ (.A(\top_ihp.oisc.regs[53][13] ),
    .B(net499),
    .Y(_03019_));
 sg13g2_a21oi_1 _18679_ (.A1(_10117_),
    .A2(net499),
    .Y(_01898_),
    .B1(_03019_));
 sg13g2_nand2_1 _18680_ (.Y(_03020_),
    .A(\top_ihp.oisc.regs[53][14] ),
    .B(net320));
 sg13g2_o21ai_1 _18681_ (.B1(_03020_),
    .Y(_01899_),
    .A1(_10841_),
    .A2(net321));
 sg13g2_buf_2 _18682_ (.A(_03013_),
    .X(_03021_));
 sg13g2_nand2_1 _18683_ (.Y(_03022_),
    .A(\top_ihp.oisc.regs[53][15] ),
    .B(net319));
 sg13g2_o21ai_1 _18684_ (.B1(_03022_),
    .Y(_01900_),
    .A1(net101),
    .A2(net321));
 sg13g2_nor2_1 _18685_ (.A(\top_ihp.oisc.regs[53][16] ),
    .B(net499),
    .Y(_03023_));
 sg13g2_a21oi_1 _18686_ (.A1(net132),
    .A2(net499),
    .Y(_01901_),
    .B1(_03023_));
 sg13g2_nand2_1 _18687_ (.Y(_03024_),
    .A(\top_ihp.oisc.regs[53][17] ),
    .B(net319));
 sg13g2_o21ai_1 _18688_ (.B1(_03024_),
    .Y(_01902_),
    .A1(net52),
    .A2(net321));
 sg13g2_nand2_1 _18689_ (.Y(_03025_),
    .A(\top_ihp.oisc.regs[53][18] ),
    .B(net319));
 sg13g2_o21ai_1 _18690_ (.B1(_03025_),
    .Y(_01903_),
    .A1(_10848_),
    .A2(net321));
 sg13g2_nand2_1 _18691_ (.Y(_03026_),
    .A(\top_ihp.oisc.regs[53][19] ),
    .B(net319));
 sg13g2_o21ai_1 _18692_ (.B1(_03026_),
    .Y(_01904_),
    .A1(net107),
    .A2(_03014_));
 sg13g2_nand2_1 _18693_ (.Y(_03027_),
    .A(\top_ihp.oisc.regs[53][1] ),
    .B(net319));
 sg13g2_o21ai_1 _18694_ (.B1(_03027_),
    .Y(_01905_),
    .A1(_10852_),
    .A2(net321));
 sg13g2_nor2_1 _18695_ (.A(\top_ihp.oisc.regs[53][20] ),
    .B(_03011_),
    .Y(_03028_));
 sg13g2_a21oi_1 _18696_ (.A1(_02693_),
    .A2(_03011_),
    .Y(_01906_),
    .B1(_03028_));
 sg13g2_nand2_1 _18697_ (.Y(_03029_),
    .A(\top_ihp.oisc.regs[53][21] ),
    .B(_03021_));
 sg13g2_o21ai_1 _18698_ (.B1(_03029_),
    .Y(_01907_),
    .A1(_10855_),
    .A2(_03014_));
 sg13g2_nor2_1 _18699_ (.A(\top_ihp.oisc.regs[53][22] ),
    .B(net499),
    .Y(_03030_));
 sg13g2_a21oi_1 _18700_ (.A1(_10130_),
    .A2(net499),
    .Y(_01908_),
    .B1(_03030_));
 sg13g2_nor2_1 _18701_ (.A(\top_ihp.oisc.regs[53][23] ),
    .B(_03010_),
    .Y(_03031_));
 sg13g2_a21oi_1 _18702_ (.A1(net100),
    .A2(net499),
    .Y(_01909_),
    .B1(_03031_));
 sg13g2_buf_1 _18703_ (.A(_03013_),
    .X(_03032_));
 sg13g2_nand2_1 _18704_ (.Y(_03033_),
    .A(\top_ihp.oisc.regs[53][24] ),
    .B(net319));
 sg13g2_o21ai_1 _18705_ (.B1(_03033_),
    .Y(_01910_),
    .A1(net106),
    .A2(net318));
 sg13g2_nand2_1 _18706_ (.Y(_03034_),
    .A(\top_ihp.oisc.regs[53][25] ),
    .B(net319));
 sg13g2_o21ai_1 _18707_ (.B1(_03034_),
    .Y(_01911_),
    .A1(_10862_),
    .A2(_03032_));
 sg13g2_nand2_1 _18708_ (.Y(_03035_),
    .A(\top_ihp.oisc.regs[53][26] ),
    .B(net319));
 sg13g2_o21ai_1 _18709_ (.B1(_03035_),
    .Y(_01912_),
    .A1(_02648_),
    .A2(_03032_));
 sg13g2_nand2_1 _18710_ (.Y(_03036_),
    .A(\top_ihp.oisc.regs[53][27] ),
    .B(_03021_));
 sg13g2_o21ai_1 _18711_ (.B1(_03036_),
    .Y(_01913_),
    .A1(_02650_),
    .A2(net318));
 sg13g2_buf_2 _18712_ (.A(_03013_),
    .X(_03037_));
 sg13g2_nand2_1 _18713_ (.Y(_03038_),
    .A(\top_ihp.oisc.regs[53][28] ),
    .B(net317));
 sg13g2_o21ai_1 _18714_ (.B1(_03038_),
    .Y(_01914_),
    .A1(_02652_),
    .A2(net318));
 sg13g2_nand2_1 _18715_ (.Y(_03039_),
    .A(\top_ihp.oisc.regs[53][29] ),
    .B(net317));
 sg13g2_o21ai_1 _18716_ (.B1(_03039_),
    .Y(_01915_),
    .A1(_02655_),
    .A2(net318));
 sg13g2_nand2_1 _18717_ (.Y(_03040_),
    .A(\top_ihp.oisc.regs[53][2] ),
    .B(_03037_));
 sg13g2_o21ai_1 _18718_ (.B1(_03040_),
    .Y(_01916_),
    .A1(net99),
    .A2(net318));
 sg13g2_nand2_1 _18719_ (.Y(_03041_),
    .A(\top_ihp.oisc.regs[53][30] ),
    .B(net317));
 sg13g2_o21ai_1 _18720_ (.B1(_03041_),
    .Y(_01917_),
    .A1(net27),
    .A2(net318));
 sg13g2_nand2_1 _18721_ (.Y(_03042_),
    .A(\top_ihp.oisc.regs[53][31] ),
    .B(_03037_));
 sg13g2_o21ai_1 _18722_ (.B1(_03042_),
    .Y(_01918_),
    .A1(net96),
    .A2(net318));
 sg13g2_nand2_1 _18723_ (.Y(_03043_),
    .A(\top_ihp.oisc.regs[53][3] ),
    .B(net317));
 sg13g2_o21ai_1 _18724_ (.B1(_03043_),
    .Y(_01919_),
    .A1(net98),
    .A2(net318));
 sg13g2_nand2_1 _18725_ (.Y(_03044_),
    .A(\top_ihp.oisc.regs[53][4] ),
    .B(net317));
 sg13g2_o21ai_1 _18726_ (.B1(_03044_),
    .Y(_01920_),
    .A1(net97),
    .A2(net320));
 sg13g2_nand2_1 _18727_ (.Y(_03045_),
    .A(\top_ihp.oisc.regs[53][5] ),
    .B(net317));
 sg13g2_o21ai_1 _18728_ (.B1(_03045_),
    .Y(_01921_),
    .A1(net104),
    .A2(net320));
 sg13g2_nand2_1 _18729_ (.Y(_03046_),
    .A(\top_ihp.oisc.regs[53][6] ),
    .B(net317));
 sg13g2_o21ai_1 _18730_ (.B1(_03046_),
    .Y(_01922_),
    .A1(net103),
    .A2(_03015_));
 sg13g2_nand2_1 _18731_ (.Y(_03047_),
    .A(\top_ihp.oisc.regs[53][7] ),
    .B(net317));
 sg13g2_o21ai_1 _18732_ (.B1(_03047_),
    .Y(_01923_),
    .A1(net187),
    .A2(net320));
 sg13g2_nand2_1 _18733_ (.Y(_03048_),
    .A(\top_ihp.oisc.regs[53][8] ),
    .B(_03013_));
 sg13g2_o21ai_1 _18734_ (.B1(_03048_),
    .Y(_01924_),
    .A1(net30),
    .A2(_03015_));
 sg13g2_nand2_1 _18735_ (.Y(_03049_),
    .A(\top_ihp.oisc.regs[53][9] ),
    .B(_03013_));
 sg13g2_o21ai_1 _18736_ (.B1(_03049_),
    .Y(_01925_),
    .A1(net29),
    .A2(net320));
 sg13g2_nand2_2 _18737_ (.Y(_03050_),
    .A(net711),
    .B(_02763_));
 sg13g2_nor2_1 _18738_ (.A(net682),
    .B(_03050_),
    .Y(_03051_));
 sg13g2_buf_2 _18739_ (.A(_03051_),
    .X(_03052_));
 sg13g2_mux2_1 _18740_ (.A0(\top_ihp.oisc.regs[54][0] ),
    .A1(net334),
    .S(_03052_),
    .X(_01926_));
 sg13g2_buf_8 _18741_ (.A(net65),
    .X(_03053_));
 sg13g2_or2_1 _18742_ (.X(_03054_),
    .B(_03050_),
    .A(net682));
 sg13g2_buf_1 _18743_ (.A(_03054_),
    .X(_03055_));
 sg13g2_buf_1 _18744_ (.A(_03055_),
    .X(_03056_));
 sg13g2_buf_1 _18745_ (.A(net498),
    .X(_03057_));
 sg13g2_buf_1 _18746_ (.A(_03055_),
    .X(_03058_));
 sg13g2_nand2_1 _18747_ (.Y(_03059_),
    .A(\top_ihp.oisc.regs[54][10] ),
    .B(net497));
 sg13g2_o21ai_1 _18748_ (.B1(_03059_),
    .Y(_01927_),
    .A1(net26),
    .A2(net316));
 sg13g2_nand2_1 _18749_ (.Y(_03060_),
    .A(\top_ihp.oisc.regs[54][11] ),
    .B(net497));
 sg13g2_o21ai_1 _18750_ (.B1(_03060_),
    .Y(_01928_),
    .A1(_02680_),
    .A2(net316));
 sg13g2_buf_2 _18751_ (.A(_09347_),
    .X(_03061_));
 sg13g2_buf_1 _18752_ (.A(net498),
    .X(_03062_));
 sg13g2_nand2_1 _18753_ (.Y(_03063_),
    .A(\top_ihp.oisc.regs[54][12] ),
    .B(net315));
 sg13g2_o21ai_1 _18754_ (.B1(_03063_),
    .Y(_01929_),
    .A1(net180),
    .A2(_03057_));
 sg13g2_nand2_1 _18755_ (.Y(_03064_),
    .A(\top_ihp.oisc.regs[54][13] ),
    .B(net315));
 sg13g2_o21ai_1 _18756_ (.B1(_03064_),
    .Y(_01930_),
    .A1(net111),
    .A2(net316));
 sg13g2_buf_1 _18757_ (.A(_10066_),
    .X(_03065_));
 sg13g2_nand2_1 _18758_ (.Y(_03066_),
    .A(\top_ihp.oisc.regs[54][14] ),
    .B(net315));
 sg13g2_o21ai_1 _18759_ (.B1(_03066_),
    .Y(_01931_),
    .A1(net95),
    .A2(net316));
 sg13g2_nand2_1 _18760_ (.Y(_03067_),
    .A(\top_ihp.oisc.regs[54][15] ),
    .B(net315));
 sg13g2_o21ai_1 _18761_ (.B1(_03067_),
    .Y(_01932_),
    .A1(net101),
    .A2(net316));
 sg13g2_nor2_1 _18762_ (.A(\top_ihp.oisc.regs[54][16] ),
    .B(_03052_),
    .Y(_03068_));
 sg13g2_a21oi_1 _18763_ (.A1(net132),
    .A2(_03052_),
    .Y(_01933_),
    .B1(_03068_));
 sg13g2_buf_1 _18764_ (.A(_09461_),
    .X(_03069_));
 sg13g2_nand2_1 _18765_ (.Y(_03070_),
    .A(\top_ihp.oisc.regs[54][17] ),
    .B(net315));
 sg13g2_o21ai_1 _18766_ (.B1(_03070_),
    .Y(_01934_),
    .A1(net94),
    .A2(_03057_));
 sg13g2_buf_1 _18767_ (.A(_09482_),
    .X(_03071_));
 sg13g2_nand2_1 _18768_ (.Y(_03072_),
    .A(\top_ihp.oisc.regs[54][18] ),
    .B(_03062_));
 sg13g2_o21ai_1 _18769_ (.B1(_03072_),
    .Y(_01935_),
    .A1(net93),
    .A2(net316));
 sg13g2_buf_1 _18770_ (.A(_10072_),
    .X(_03073_));
 sg13g2_nand2_1 _18771_ (.Y(_03074_),
    .A(\top_ihp.oisc.regs[54][19] ),
    .B(net315));
 sg13g2_o21ai_1 _18772_ (.B1(_03074_),
    .Y(_01936_),
    .A1(net92),
    .A2(net316));
 sg13g2_buf_1 _18773_ (.A(_09552_),
    .X(_03075_));
 sg13g2_nand2_1 _18774_ (.Y(_03076_),
    .A(\top_ihp.oisc.regs[54][1] ),
    .B(_03062_));
 sg13g2_o21ai_1 _18775_ (.B1(_03076_),
    .Y(_01937_),
    .A1(_03075_),
    .A2(net316));
 sg13g2_nor2_1 _18776_ (.A(\top_ihp.oisc.regs[54][20] ),
    .B(_03052_),
    .Y(_03077_));
 sg13g2_a21oi_1 _18777_ (.A1(net28),
    .A2(_03052_),
    .Y(_01938_),
    .B1(_03077_));
 sg13g2_buf_1 _18778_ (.A(_09598_),
    .X(_03078_));
 sg13g2_buf_1 _18779_ (.A(net498),
    .X(_03079_));
 sg13g2_nand2_1 _18780_ (.Y(_03080_),
    .A(\top_ihp.oisc.regs[54][21] ),
    .B(net315));
 sg13g2_o21ai_1 _18781_ (.B1(_03080_),
    .Y(_01939_),
    .A1(net46),
    .A2(net314));
 sg13g2_nand2_1 _18782_ (.Y(_03081_),
    .A(\top_ihp.oisc.regs[54][22] ),
    .B(net315));
 sg13g2_o21ai_1 _18783_ (.B1(_03081_),
    .Y(_01940_),
    .A1(net110),
    .A2(net314));
 sg13g2_nor2_1 _18784_ (.A(\top_ihp.oisc.regs[54][23] ),
    .B(_03052_),
    .Y(_03082_));
 sg13g2_a21oi_1 _18785_ (.A1(net100),
    .A2(_03052_),
    .Y(_01941_),
    .B1(_03082_));
 sg13g2_buf_1 _18786_ (.A(_10077_),
    .X(_03083_));
 sg13g2_buf_1 _18787_ (.A(net498),
    .X(_03084_));
 sg13g2_nand2_1 _18788_ (.Y(_03085_),
    .A(\top_ihp.oisc.regs[54][24] ),
    .B(net313));
 sg13g2_o21ai_1 _18789_ (.B1(_03085_),
    .Y(_01942_),
    .A1(_03083_),
    .A2(net314));
 sg13g2_buf_1 _18790_ (.A(_09668_),
    .X(_03086_));
 sg13g2_nand2_1 _18791_ (.Y(_03087_),
    .A(\top_ihp.oisc.regs[54][25] ),
    .B(net313));
 sg13g2_o21ai_1 _18792_ (.B1(_03087_),
    .Y(_01943_),
    .A1(net179),
    .A2(net314));
 sg13g2_buf_1 _18793_ (.A(_09678_),
    .X(_03088_));
 sg13g2_nand2_1 _18794_ (.Y(_03089_),
    .A(\top_ihp.oisc.regs[54][26] ),
    .B(net313));
 sg13g2_o21ai_1 _18795_ (.B1(_03089_),
    .Y(_01944_),
    .A1(net90),
    .A2(net314));
 sg13g2_buf_8 _18796_ (.A(_09702_),
    .X(_03090_));
 sg13g2_nand2_1 _18797_ (.Y(_03091_),
    .A(\top_ihp.oisc.regs[54][27] ),
    .B(net313));
 sg13g2_o21ai_1 _18798_ (.B1(_03091_),
    .Y(_01945_),
    .A1(net45),
    .A2(net314));
 sg13g2_buf_8 _18799_ (.A(_09713_),
    .X(_03092_));
 sg13g2_nand2_1 _18800_ (.Y(_03093_),
    .A(\top_ihp.oisc.regs[54][28] ),
    .B(net313));
 sg13g2_o21ai_1 _18801_ (.B1(_03093_),
    .Y(_01946_),
    .A1(net44),
    .A2(net314));
 sg13g2_buf_2 _18802_ (.A(_10083_),
    .X(_03094_));
 sg13g2_nand2_1 _18803_ (.Y(_03095_),
    .A(\top_ihp.oisc.regs[54][29] ),
    .B(net313));
 sg13g2_o21ai_1 _18804_ (.B1(_03095_),
    .Y(_01947_),
    .A1(net43),
    .A2(net314));
 sg13g2_nand2_1 _18805_ (.Y(_03096_),
    .A(\top_ihp.oisc.regs[54][2] ),
    .B(_03084_));
 sg13g2_o21ai_1 _18806_ (.B1(_03096_),
    .Y(_01948_),
    .A1(net99),
    .A2(_03079_));
 sg13g2_nand2_1 _18807_ (.Y(_03097_),
    .A(\top_ihp.oisc.regs[54][30] ),
    .B(_03084_));
 sg13g2_o21ai_1 _18808_ (.B1(_03097_),
    .Y(_01949_),
    .A1(net27),
    .A2(_03079_));
 sg13g2_nand2_1 _18809_ (.Y(_03098_),
    .A(\top_ihp.oisc.regs[54][31] ),
    .B(net313));
 sg13g2_o21ai_1 _18810_ (.B1(_03098_),
    .Y(_01950_),
    .A1(net96),
    .A2(net497));
 sg13g2_nand2_1 _18811_ (.Y(_03099_),
    .A(\top_ihp.oisc.regs[54][3] ),
    .B(net313));
 sg13g2_o21ai_1 _18812_ (.B1(_03099_),
    .Y(_01951_),
    .A1(net98),
    .A2(net497));
 sg13g2_nand2_1 _18813_ (.Y(_03100_),
    .A(\top_ihp.oisc.regs[54][4] ),
    .B(net498));
 sg13g2_o21ai_1 _18814_ (.B1(_03100_),
    .Y(_01952_),
    .A1(net97),
    .A2(net497));
 sg13g2_buf_2 _18815_ (.A(_09871_),
    .X(_03101_));
 sg13g2_nand2_1 _18816_ (.Y(_03102_),
    .A(\top_ihp.oisc.regs[54][5] ),
    .B(net498));
 sg13g2_o21ai_1 _18817_ (.B1(_03102_),
    .Y(_01953_),
    .A1(net178),
    .A2(net497));
 sg13g2_buf_2 _18818_ (.A(_09894_),
    .X(_03103_));
 sg13g2_nand2_1 _18819_ (.Y(_03104_),
    .A(\top_ihp.oisc.regs[54][6] ),
    .B(net498));
 sg13g2_o21ai_1 _18820_ (.B1(_03104_),
    .Y(_01954_),
    .A1(net177),
    .A2(net497));
 sg13g2_nand2_1 _18821_ (.Y(_03105_),
    .A(\top_ihp.oisc.regs[54][7] ),
    .B(_03056_));
 sg13g2_o21ai_1 _18822_ (.B1(_03105_),
    .Y(_01955_),
    .A1(net47),
    .A2(_03058_));
 sg13g2_buf_2 _18823_ (.A(_09929_),
    .X(_03106_));
 sg13g2_nand2_1 _18824_ (.Y(_03107_),
    .A(\top_ihp.oisc.regs[54][8] ),
    .B(_03056_));
 sg13g2_o21ai_1 _18825_ (.B1(_03107_),
    .Y(_01956_),
    .A1(net42),
    .A2(_03058_));
 sg13g2_buf_8 _18826_ (.A(net60),
    .X(_03108_));
 sg13g2_nand2_1 _18827_ (.Y(_03109_),
    .A(\top_ihp.oisc.regs[54][9] ),
    .B(net498));
 sg13g2_o21ai_1 _18828_ (.B1(_03109_),
    .Y(_01957_),
    .A1(net25),
    .A2(net497));
 sg13g2_nand2_2 _18829_ (.Y(_03110_),
    .A(_10009_),
    .B(_02763_));
 sg13g2_nor2_1 _18830_ (.A(net682),
    .B(_03110_),
    .Y(_03111_));
 sg13g2_buf_1 _18831_ (.A(_03111_),
    .X(_03112_));
 sg13g2_mux2_1 _18832_ (.A0(\top_ihp.oisc.regs[55][0] ),
    .A1(net334),
    .S(net631),
    .X(_01958_));
 sg13g2_or2_1 _18833_ (.X(_03113_),
    .B(_03110_),
    .A(_10460_));
 sg13g2_buf_2 _18834_ (.A(_03113_),
    .X(_03114_));
 sg13g2_buf_2 _18835_ (.A(_03114_),
    .X(_03115_));
 sg13g2_buf_1 _18836_ (.A(_03114_),
    .X(_03116_));
 sg13g2_nand2_1 _18837_ (.Y(_03117_),
    .A(\top_ihp.oisc.regs[55][10] ),
    .B(net494));
 sg13g2_o21ai_1 _18838_ (.B1(_03117_),
    .Y(_01959_),
    .A1(net26),
    .A2(net495));
 sg13g2_buf_1 _18839_ (.A(net251),
    .X(_03118_));
 sg13g2_nand2_1 _18840_ (.Y(_03119_),
    .A(\top_ihp.oisc.regs[55][11] ),
    .B(net494));
 sg13g2_o21ai_1 _18841_ (.B1(_03119_),
    .Y(_01960_),
    .A1(net89),
    .A2(net495));
 sg13g2_nand2_1 _18842_ (.Y(_03120_),
    .A(\top_ihp.oisc.regs[55][12] ),
    .B(net494));
 sg13g2_o21ai_1 _18843_ (.B1(_03120_),
    .Y(_01961_),
    .A1(net180),
    .A2(net495));
 sg13g2_nor2_1 _18844_ (.A(\top_ihp.oisc.regs[55][13] ),
    .B(net631),
    .Y(_03121_));
 sg13g2_a21oi_1 _18845_ (.A1(_10117_),
    .A2(net631),
    .Y(_01962_),
    .B1(_03121_));
 sg13g2_nand2_1 _18846_ (.Y(_03122_),
    .A(\top_ihp.oisc.regs[55][14] ),
    .B(net494));
 sg13g2_o21ai_1 _18847_ (.B1(_03122_),
    .Y(_01963_),
    .A1(net95),
    .A2(net495));
 sg13g2_buf_1 _18848_ (.A(_09418_),
    .X(_03123_));
 sg13g2_buf_1 _18849_ (.A(_03114_),
    .X(_03124_));
 sg13g2_nand2_1 _18850_ (.Y(_03125_),
    .A(\top_ihp.oisc.regs[55][15] ),
    .B(net493));
 sg13g2_o21ai_1 _18851_ (.B1(_03125_),
    .Y(_01964_),
    .A1(net176),
    .A2(net495));
 sg13g2_nor2_1 _18852_ (.A(\top_ihp.oisc.regs[55][16] ),
    .B(net631),
    .Y(_03126_));
 sg13g2_a21oi_1 _18853_ (.A1(net146),
    .A2(net631),
    .Y(_01965_),
    .B1(_03126_));
 sg13g2_nand2_1 _18854_ (.Y(_03127_),
    .A(\top_ihp.oisc.regs[55][17] ),
    .B(net493));
 sg13g2_o21ai_1 _18855_ (.B1(_03127_),
    .Y(_01966_),
    .A1(net94),
    .A2(net495));
 sg13g2_nand2_1 _18856_ (.Y(_03128_),
    .A(\top_ihp.oisc.regs[55][18] ),
    .B(net493));
 sg13g2_o21ai_1 _18857_ (.B1(_03128_),
    .Y(_01967_),
    .A1(_03071_),
    .A2(_03115_));
 sg13g2_nand2_1 _18858_ (.Y(_03129_),
    .A(\top_ihp.oisc.regs[55][19] ),
    .B(net493));
 sg13g2_o21ai_1 _18859_ (.B1(_03129_),
    .Y(_01968_),
    .A1(_03073_),
    .A2(net495));
 sg13g2_nand2_1 _18860_ (.Y(_03130_),
    .A(\top_ihp.oisc.regs[55][1] ),
    .B(net493));
 sg13g2_o21ai_1 _18861_ (.B1(_03130_),
    .Y(_01969_),
    .A1(net496),
    .A2(net495));
 sg13g2_nor2_1 _18862_ (.A(\top_ihp.oisc.regs[55][20] ),
    .B(net631),
    .Y(_03131_));
 sg13g2_a21oi_1 _18863_ (.A1(net28),
    .A2(net631),
    .Y(_01970_),
    .B1(_03131_));
 sg13g2_nand2_1 _18864_ (.Y(_03132_),
    .A(\top_ihp.oisc.regs[55][21] ),
    .B(net493));
 sg13g2_o21ai_1 _18865_ (.B1(_03132_),
    .Y(_01971_),
    .A1(net46),
    .A2(_03115_));
 sg13g2_nor2_1 _18866_ (.A(\top_ihp.oisc.regs[55][22] ),
    .B(_03112_),
    .Y(_03133_));
 sg13g2_a21oi_1 _18867_ (.A1(_10130_),
    .A2(_03112_),
    .Y(_01972_),
    .B1(_03133_));
 sg13g2_nor2_1 _18868_ (.A(\top_ihp.oisc.regs[55][23] ),
    .B(_03111_),
    .Y(_03134_));
 sg13g2_a21oi_1 _18869_ (.A1(net100),
    .A2(net631),
    .Y(_01973_),
    .B1(_03134_));
 sg13g2_buf_1 _18870_ (.A(_03114_),
    .X(_03135_));
 sg13g2_nand2_1 _18871_ (.Y(_03136_),
    .A(\top_ihp.oisc.regs[55][24] ),
    .B(_03124_));
 sg13g2_o21ai_1 _18872_ (.B1(_03136_),
    .Y(_01974_),
    .A1(net91),
    .A2(net492));
 sg13g2_nand2_1 _18873_ (.Y(_03137_),
    .A(\top_ihp.oisc.regs[55][25] ),
    .B(net493));
 sg13g2_o21ai_1 _18874_ (.B1(_03137_),
    .Y(_01975_),
    .A1(net179),
    .A2(net492));
 sg13g2_nand2_1 _18875_ (.Y(_03138_),
    .A(\top_ihp.oisc.regs[55][26] ),
    .B(net493));
 sg13g2_o21ai_1 _18876_ (.B1(_03138_),
    .Y(_01976_),
    .A1(net90),
    .A2(net492));
 sg13g2_nand2_1 _18877_ (.Y(_03139_),
    .A(\top_ihp.oisc.regs[55][27] ),
    .B(_03124_));
 sg13g2_o21ai_1 _18878_ (.B1(_03139_),
    .Y(_01977_),
    .A1(net45),
    .A2(net492));
 sg13g2_buf_1 _18879_ (.A(_03114_),
    .X(_03140_));
 sg13g2_nand2_1 _18880_ (.Y(_03141_),
    .A(\top_ihp.oisc.regs[55][28] ),
    .B(net491));
 sg13g2_o21ai_1 _18881_ (.B1(_03141_),
    .Y(_01978_),
    .A1(_03092_),
    .A2(net492));
 sg13g2_nand2_1 _18882_ (.Y(_03142_),
    .A(\top_ihp.oisc.regs[55][29] ),
    .B(net491));
 sg13g2_o21ai_1 _18883_ (.B1(_03142_),
    .Y(_01979_),
    .A1(net43),
    .A2(net492));
 sg13g2_buf_2 _18884_ (.A(_09753_),
    .X(_03143_));
 sg13g2_nand2_1 _18885_ (.Y(_03144_),
    .A(\top_ihp.oisc.regs[55][2] ),
    .B(net491));
 sg13g2_o21ai_1 _18886_ (.B1(_03144_),
    .Y(_01980_),
    .A1(net175),
    .A2(net492));
 sg13g2_buf_2 _18887_ (.A(_09761_),
    .X(_03145_));
 sg13g2_nand2_1 _18888_ (.Y(_03146_),
    .A(\top_ihp.oisc.regs[55][30] ),
    .B(net491));
 sg13g2_o21ai_1 _18889_ (.B1(_03146_),
    .Y(_01981_),
    .A1(net41),
    .A2(net492));
 sg13g2_nand2_1 _18890_ (.Y(_03147_),
    .A(\top_ihp.oisc.regs[55][31] ),
    .B(net491));
 sg13g2_o21ai_1 _18891_ (.B1(_03147_),
    .Y(_01982_),
    .A1(_02753_),
    .A2(_03135_));
 sg13g2_buf_2 _18892_ (.A(_09807_),
    .X(_03148_));
 sg13g2_nand2_1 _18893_ (.Y(_03149_),
    .A(\top_ihp.oisc.regs[55][3] ),
    .B(net491));
 sg13g2_o21ai_1 _18894_ (.B1(_03149_),
    .Y(_01983_),
    .A1(net174),
    .A2(_03135_));
 sg13g2_buf_1 _18895_ (.A(net220),
    .X(_03150_));
 sg13g2_nand2_1 _18896_ (.Y(_03151_),
    .A(\top_ihp.oisc.regs[55][4] ),
    .B(net491));
 sg13g2_o21ai_1 _18897_ (.B1(_03151_),
    .Y(_01984_),
    .A1(net88),
    .A2(net494));
 sg13g2_nand2_1 _18898_ (.Y(_03152_),
    .A(\top_ihp.oisc.regs[55][5] ),
    .B(net491));
 sg13g2_o21ai_1 _18899_ (.B1(_03152_),
    .Y(_01985_),
    .A1(net178),
    .A2(net494));
 sg13g2_nand2_1 _18900_ (.Y(_03153_),
    .A(\top_ihp.oisc.regs[55][6] ),
    .B(_03140_));
 sg13g2_o21ai_1 _18901_ (.B1(_03153_),
    .Y(_01986_),
    .A1(net177),
    .A2(_03116_));
 sg13g2_nand2_1 _18902_ (.Y(_03154_),
    .A(\top_ihp.oisc.regs[55][7] ),
    .B(_03140_));
 sg13g2_o21ai_1 _18903_ (.B1(_03154_),
    .Y(_01987_),
    .A1(_02666_),
    .A2(_03116_));
 sg13g2_nand2_1 _18904_ (.Y(_03155_),
    .A(\top_ihp.oisc.regs[55][8] ),
    .B(_03114_));
 sg13g2_o21ai_1 _18905_ (.B1(_03155_),
    .Y(_01988_),
    .A1(net42),
    .A2(net494));
 sg13g2_nand2_1 _18906_ (.Y(_03156_),
    .A(\top_ihp.oisc.regs[55][9] ),
    .B(_03114_));
 sg13g2_o21ai_1 _18907_ (.B1(_03156_),
    .Y(_01989_),
    .A1(net25),
    .A2(net494));
 sg13g2_nand2b_1 _18908_ (.Y(_03157_),
    .B(_02968_),
    .A_N(_09956_));
 sg13g2_buf_1 _18909_ (.A(_03157_),
    .X(_03158_));
 sg13g2_buf_2 _18910_ (.A(net490),
    .X(_03159_));
 sg13g2_mux2_1 _18911_ (.A0(_09946_),
    .A1(\top_ihp.oisc.regs[56][0] ),
    .S(_03159_),
    .X(_01990_));
 sg13g2_nand2_1 _18912_ (.Y(_03160_),
    .A(net545),
    .B(_02968_));
 sg13g2_buf_2 _18913_ (.A(_03160_),
    .X(_03161_));
 sg13g2_nand2_1 _18914_ (.Y(_03162_),
    .A(\top_ihp.oisc.regs[56][10] ),
    .B(net312));
 sg13g2_o21ai_1 _18915_ (.B1(_03162_),
    .Y(_01991_),
    .A1(net26),
    .A2(_03161_));
 sg13g2_buf_1 _18916_ (.A(net490),
    .X(_03163_));
 sg13g2_nand2_1 _18917_ (.Y(_03164_),
    .A(\top_ihp.oisc.regs[56][11] ),
    .B(net311));
 sg13g2_o21ai_1 _18918_ (.B1(_03164_),
    .Y(_01992_),
    .A1(net89),
    .A2(_03161_));
 sg13g2_buf_1 _18919_ (.A(net490),
    .X(_03165_));
 sg13g2_nand2_1 _18920_ (.Y(_03166_),
    .A(\top_ihp.oisc.regs[56][12] ),
    .B(net311));
 sg13g2_o21ai_1 _18921_ (.B1(_03166_),
    .Y(_01993_),
    .A1(net180),
    .A2(net310));
 sg13g2_and2_1 _18922_ (.A(_10029_),
    .B(_02968_),
    .X(_03167_));
 sg13g2_buf_1 _18923_ (.A(_03167_),
    .X(_03168_));
 sg13g2_nor2_1 _18924_ (.A(\top_ihp.oisc.regs[56][13] ),
    .B(net173),
    .Y(_03169_));
 sg13g2_a21oi_1 _18925_ (.A1(net73),
    .A2(net173),
    .Y(_01994_),
    .B1(_03169_));
 sg13g2_nand2_1 _18926_ (.Y(_03170_),
    .A(\top_ihp.oisc.regs[56][14] ),
    .B(net311));
 sg13g2_o21ai_1 _18927_ (.B1(_03170_),
    .Y(_01995_),
    .A1(net95),
    .A2(net310));
 sg13g2_nand2_1 _18928_ (.Y(_03171_),
    .A(\top_ihp.oisc.regs[56][15] ),
    .B(net311));
 sg13g2_o21ai_1 _18929_ (.B1(_03171_),
    .Y(_01996_),
    .A1(net176),
    .A2(net310));
 sg13g2_nor2_1 _18930_ (.A(\top_ihp.oisc.regs[56][16] ),
    .B(net173),
    .Y(_03172_));
 sg13g2_a21oi_1 _18931_ (.A1(net146),
    .A2(net173),
    .Y(_01997_),
    .B1(_03172_));
 sg13g2_nand2_1 _18932_ (.Y(_03173_),
    .A(\top_ihp.oisc.regs[56][17] ),
    .B(net311));
 sg13g2_o21ai_1 _18933_ (.B1(_03173_),
    .Y(_01998_),
    .A1(net94),
    .A2(net310));
 sg13g2_nand2_1 _18934_ (.Y(_03174_),
    .A(\top_ihp.oisc.regs[56][18] ),
    .B(net311));
 sg13g2_o21ai_1 _18935_ (.B1(_03174_),
    .Y(_01999_),
    .A1(net93),
    .A2(net310));
 sg13g2_nand2_1 _18936_ (.Y(_03175_),
    .A(\top_ihp.oisc.regs[56][19] ),
    .B(net311));
 sg13g2_o21ai_1 _18937_ (.B1(_03175_),
    .Y(_02000_),
    .A1(net92),
    .A2(net310));
 sg13g2_nand2_1 _18938_ (.Y(_03176_),
    .A(\top_ihp.oisc.regs[56][1] ),
    .B(_03163_));
 sg13g2_o21ai_1 _18939_ (.B1(_03176_),
    .Y(_02001_),
    .A1(net496),
    .A2(_03165_));
 sg13g2_nor2_1 _18940_ (.A(\top_ihp.oisc.regs[56][20] ),
    .B(net173),
    .Y(_03177_));
 sg13g2_a21oi_1 _18941_ (.A1(net28),
    .A2(net173),
    .Y(_02002_),
    .B1(_03177_));
 sg13g2_nand2_1 _18942_ (.Y(_03178_),
    .A(\top_ihp.oisc.regs[56][21] ),
    .B(net311));
 sg13g2_o21ai_1 _18943_ (.B1(_03178_),
    .Y(_02003_),
    .A1(net46),
    .A2(net310));
 sg13g2_nor2_1 _18944_ (.A(\top_ihp.oisc.regs[56][22] ),
    .B(_03168_),
    .Y(_03179_));
 sg13g2_a21oi_1 _18945_ (.A1(net143),
    .A2(_03168_),
    .Y(_02004_),
    .B1(_03179_));
 sg13g2_nor2_1 _18946_ (.A(\top_ihp.oisc.regs[56][23] ),
    .B(net173),
    .Y(_03180_));
 sg13g2_a21oi_1 _18947_ (.A1(_02697_),
    .A2(net173),
    .Y(_02005_),
    .B1(_03180_));
 sg13g2_nand2_1 _18948_ (.Y(_03181_),
    .A(\top_ihp.oisc.regs[56][24] ),
    .B(_03163_));
 sg13g2_o21ai_1 _18949_ (.B1(_03181_),
    .Y(_02006_),
    .A1(net91),
    .A2(_03161_));
 sg13g2_buf_1 _18950_ (.A(net490),
    .X(_03182_));
 sg13g2_nand2_1 _18951_ (.Y(_03183_),
    .A(\top_ihp.oisc.regs[56][25] ),
    .B(net309));
 sg13g2_o21ai_1 _18952_ (.B1(_03183_),
    .Y(_02007_),
    .A1(net179),
    .A2(_03165_));
 sg13g2_nand2_1 _18953_ (.Y(_03184_),
    .A(\top_ihp.oisc.regs[56][26] ),
    .B(net309));
 sg13g2_o21ai_1 _18954_ (.B1(_03184_),
    .Y(_02008_),
    .A1(net90),
    .A2(net310));
 sg13g2_nand2_1 _18955_ (.Y(_03185_),
    .A(\top_ihp.oisc.regs[56][27] ),
    .B(net309));
 sg13g2_o21ai_1 _18956_ (.B1(_03185_),
    .Y(_02009_),
    .A1(_03090_),
    .A2(_03161_));
 sg13g2_nand2_1 _18957_ (.Y(_03186_),
    .A(\top_ihp.oisc.regs[56][28] ),
    .B(net309));
 sg13g2_o21ai_1 _18958_ (.B1(_03186_),
    .Y(_02010_),
    .A1(net44),
    .A2(net312));
 sg13g2_nand2_1 _18959_ (.Y(_03187_),
    .A(\top_ihp.oisc.regs[56][29] ),
    .B(net309));
 sg13g2_o21ai_1 _18960_ (.B1(_03187_),
    .Y(_02011_),
    .A1(net43),
    .A2(_03159_));
 sg13g2_nand2_1 _18961_ (.Y(_03188_),
    .A(\top_ihp.oisc.regs[56][2] ),
    .B(_03182_));
 sg13g2_o21ai_1 _18962_ (.B1(_03188_),
    .Y(_02012_),
    .A1(net175),
    .A2(net312));
 sg13g2_nand2_1 _18963_ (.Y(_03189_),
    .A(\top_ihp.oisc.regs[56][30] ),
    .B(_03182_));
 sg13g2_o21ai_1 _18964_ (.B1(_03189_),
    .Y(_02013_),
    .A1(net41),
    .A2(net312));
 sg13g2_buf_8 _18965_ (.A(_09781_),
    .X(_03190_));
 sg13g2_nand2_1 _18966_ (.Y(_03191_),
    .A(\top_ihp.oisc.regs[56][31] ),
    .B(net309));
 sg13g2_o21ai_1 _18967_ (.B1(_03191_),
    .Y(_02014_),
    .A1(net87),
    .A2(_03161_));
 sg13g2_nand2_1 _18968_ (.Y(_03192_),
    .A(\top_ihp.oisc.regs[56][3] ),
    .B(net309));
 sg13g2_o21ai_1 _18969_ (.B1(_03192_),
    .Y(_02015_),
    .A1(net174),
    .A2(net312));
 sg13g2_nand2_1 _18970_ (.Y(_03193_),
    .A(\top_ihp.oisc.regs[56][4] ),
    .B(net309));
 sg13g2_o21ai_1 _18971_ (.B1(_03193_),
    .Y(_02016_),
    .A1(_03150_),
    .A2(_03161_));
 sg13g2_nand2_1 _18972_ (.Y(_03194_),
    .A(\top_ihp.oisc.regs[56][5] ),
    .B(net490));
 sg13g2_o21ai_1 _18973_ (.B1(_03194_),
    .Y(_02017_),
    .A1(net178),
    .A2(net312));
 sg13g2_nand2_1 _18974_ (.Y(_03195_),
    .A(\top_ihp.oisc.regs[56][6] ),
    .B(net490));
 sg13g2_o21ai_1 _18975_ (.B1(_03195_),
    .Y(_02018_),
    .A1(net177),
    .A2(net312));
 sg13g2_nand2_1 _18976_ (.Y(_03196_),
    .A(\top_ihp.oisc.regs[56][7] ),
    .B(_03158_));
 sg13g2_o21ai_1 _18977_ (.B1(_03196_),
    .Y(_02019_),
    .A1(net187),
    .A2(net312));
 sg13g2_nand2_1 _18978_ (.Y(_03197_),
    .A(\top_ihp.oisc.regs[56][8] ),
    .B(net490));
 sg13g2_o21ai_1 _18979_ (.B1(_03197_),
    .Y(_02020_),
    .A1(net42),
    .A2(_03161_));
 sg13g2_nand2_1 _18980_ (.Y(_03198_),
    .A(\top_ihp.oisc.regs[56][9] ),
    .B(net490));
 sg13g2_o21ai_1 _18981_ (.B1(_03198_),
    .Y(_02021_),
    .A1(net25),
    .A2(_03161_));
 sg13g2_nor2_2 _18982_ (.A(_09958_),
    .B(_03009_),
    .Y(_03199_));
 sg13g2_mux2_1 _18983_ (.A0(\top_ihp.oisc.regs[57][0] ),
    .A1(_02845_),
    .S(_03199_),
    .X(_02022_));
 sg13g2_or2_1 _18984_ (.X(_03200_),
    .B(_03009_),
    .A(_09958_));
 sg13g2_buf_1 _18985_ (.A(_03200_),
    .X(_03201_));
 sg13g2_buf_8 _18986_ (.A(_03201_),
    .X(_03202_));
 sg13g2_buf_1 _18987_ (.A(net172),
    .X(_03203_));
 sg13g2_buf_2 _18988_ (.A(_03201_),
    .X(_03204_));
 sg13g2_nand2_1 _18989_ (.Y(_03205_),
    .A(\top_ihp.oisc.regs[57][10] ),
    .B(net171));
 sg13g2_o21ai_1 _18990_ (.B1(_03205_),
    .Y(_02023_),
    .A1(net26),
    .A2(_03203_));
 sg13g2_buf_1 _18991_ (.A(_03201_),
    .X(_03206_));
 sg13g2_nand2_1 _18992_ (.Y(_03207_),
    .A(\top_ihp.oisc.regs[57][11] ),
    .B(net170));
 sg13g2_o21ai_1 _18993_ (.B1(_03207_),
    .Y(_02024_),
    .A1(net89),
    .A2(net86));
 sg13g2_nand2_1 _18994_ (.Y(_03208_),
    .A(\top_ihp.oisc.regs[57][12] ),
    .B(_03206_));
 sg13g2_o21ai_1 _18995_ (.B1(_03208_),
    .Y(_02025_),
    .A1(_03061_),
    .A2(_03203_));
 sg13g2_nand2_1 _18996_ (.Y(_03209_),
    .A(\top_ihp.oisc.regs[57][13] ),
    .B(net170));
 sg13g2_o21ai_1 _18997_ (.B1(_03209_),
    .Y(_02026_),
    .A1(net111),
    .A2(net86));
 sg13g2_nand2_1 _18998_ (.Y(_03210_),
    .A(\top_ihp.oisc.regs[57][14] ),
    .B(_03206_));
 sg13g2_o21ai_1 _18999_ (.B1(_03210_),
    .Y(_02027_),
    .A1(_03065_),
    .A2(net86));
 sg13g2_nand2_1 _19000_ (.Y(_03211_),
    .A(\top_ihp.oisc.regs[57][15] ),
    .B(net170));
 sg13g2_o21ai_1 _19001_ (.B1(_03211_),
    .Y(_02028_),
    .A1(_03123_),
    .A2(net86));
 sg13g2_nand2_1 _19002_ (.Y(_03212_),
    .A(\top_ihp.oisc.regs[57][16] ),
    .B(net170));
 sg13g2_o21ai_1 _19003_ (.B1(_03212_),
    .Y(_02029_),
    .A1(_10762_),
    .A2(net86));
 sg13g2_nand2_1 _19004_ (.Y(_03213_),
    .A(\top_ihp.oisc.regs[57][17] ),
    .B(net170));
 sg13g2_o21ai_1 _19005_ (.B1(_03213_),
    .Y(_02030_),
    .A1(_03069_),
    .A2(net86));
 sg13g2_nand2_1 _19006_ (.Y(_03214_),
    .A(\top_ihp.oisc.regs[57][18] ),
    .B(net170));
 sg13g2_o21ai_1 _19007_ (.B1(_03214_),
    .Y(_02031_),
    .A1(net93),
    .A2(net86));
 sg13g2_nand2_1 _19008_ (.Y(_03215_),
    .A(\top_ihp.oisc.regs[57][19] ),
    .B(net170));
 sg13g2_o21ai_1 _19009_ (.B1(_03215_),
    .Y(_02032_),
    .A1(_03073_),
    .A2(net86));
 sg13g2_buf_1 _19010_ (.A(net172),
    .X(_03216_));
 sg13g2_nand2_1 _19011_ (.Y(_03217_),
    .A(\top_ihp.oisc.regs[57][1] ),
    .B(net170));
 sg13g2_o21ai_1 _19012_ (.B1(_03217_),
    .Y(_02033_),
    .A1(net496),
    .A2(net85));
 sg13g2_mux2_1 _19013_ (.A0(\top_ihp.oisc.regs[57][20] ),
    .A1(net245),
    .S(_03199_),
    .X(_02034_));
 sg13g2_buf_1 _19014_ (.A(_03201_),
    .X(_03218_));
 sg13g2_nand2_1 _19015_ (.Y(_03219_),
    .A(\top_ihp.oisc.regs[57][21] ),
    .B(net169));
 sg13g2_o21ai_1 _19016_ (.B1(_03219_),
    .Y(_02035_),
    .A1(net46),
    .A2(net85));
 sg13g2_nand2_1 _19017_ (.Y(_03220_),
    .A(\top_ihp.oisc.regs[57][22] ),
    .B(net169));
 sg13g2_o21ai_1 _19018_ (.B1(_03220_),
    .Y(_02036_),
    .A1(net110),
    .A2(net85));
 sg13g2_mux2_1 _19019_ (.A0(\top_ihp.oisc.regs[57][23] ),
    .A1(_10035_),
    .S(_03199_),
    .X(_02037_));
 sg13g2_nand2_1 _19020_ (.Y(_03221_),
    .A(\top_ihp.oisc.regs[57][24] ),
    .B(net169));
 sg13g2_o21ai_1 _19021_ (.B1(_03221_),
    .Y(_02038_),
    .A1(net91),
    .A2(net85));
 sg13g2_nand2_1 _19022_ (.Y(_03222_),
    .A(\top_ihp.oisc.regs[57][25] ),
    .B(net169));
 sg13g2_o21ai_1 _19023_ (.B1(_03222_),
    .Y(_02039_),
    .A1(net179),
    .A2(net85));
 sg13g2_nand2_1 _19024_ (.Y(_03223_),
    .A(\top_ihp.oisc.regs[57][26] ),
    .B(net169));
 sg13g2_o21ai_1 _19025_ (.B1(_03223_),
    .Y(_02040_),
    .A1(net90),
    .A2(net85));
 sg13g2_nand2_1 _19026_ (.Y(_03224_),
    .A(\top_ihp.oisc.regs[57][27] ),
    .B(net169));
 sg13g2_o21ai_1 _19027_ (.B1(_03224_),
    .Y(_02041_),
    .A1(net45),
    .A2(net85));
 sg13g2_nand2_1 _19028_ (.Y(_03225_),
    .A(\top_ihp.oisc.regs[57][28] ),
    .B(net169));
 sg13g2_o21ai_1 _19029_ (.B1(_03225_),
    .Y(_02042_),
    .A1(net44),
    .A2(_03216_));
 sg13g2_nand2_1 _19030_ (.Y(_03226_),
    .A(\top_ihp.oisc.regs[57][29] ),
    .B(net169));
 sg13g2_o21ai_1 _19031_ (.B1(_03226_),
    .Y(_02043_),
    .A1(net43),
    .A2(net85));
 sg13g2_nand2_1 _19032_ (.Y(_03227_),
    .A(\top_ihp.oisc.regs[57][2] ),
    .B(_03218_));
 sg13g2_o21ai_1 _19033_ (.B1(_03227_),
    .Y(_02044_),
    .A1(net175),
    .A2(_03216_));
 sg13g2_nand2_1 _19034_ (.Y(_03228_),
    .A(\top_ihp.oisc.regs[57][30] ),
    .B(_03218_));
 sg13g2_o21ai_1 _19035_ (.B1(_03228_),
    .Y(_02045_),
    .A1(net41),
    .A2(net171));
 sg13g2_nand2_1 _19036_ (.Y(_03229_),
    .A(\top_ihp.oisc.regs[57][31] ),
    .B(net172));
 sg13g2_o21ai_1 _19037_ (.B1(_03229_),
    .Y(_02046_),
    .A1(net87),
    .A2(net171));
 sg13g2_nand2_1 _19038_ (.Y(_03230_),
    .A(\top_ihp.oisc.regs[57][3] ),
    .B(net172));
 sg13g2_o21ai_1 _19039_ (.B1(_03230_),
    .Y(_02047_),
    .A1(net174),
    .A2(net171));
 sg13g2_nand2_1 _19040_ (.Y(_03231_),
    .A(\top_ihp.oisc.regs[57][4] ),
    .B(net172));
 sg13g2_o21ai_1 _19041_ (.B1(_03231_),
    .Y(_02048_),
    .A1(net88),
    .A2(net171));
 sg13g2_nand2_1 _19042_ (.Y(_03232_),
    .A(\top_ihp.oisc.regs[57][5] ),
    .B(net172));
 sg13g2_o21ai_1 _19043_ (.B1(_03232_),
    .Y(_02049_),
    .A1(net178),
    .A2(net171));
 sg13g2_nand2_1 _19044_ (.Y(_03233_),
    .A(\top_ihp.oisc.regs[57][6] ),
    .B(_03202_));
 sg13g2_o21ai_1 _19045_ (.B1(_03233_),
    .Y(_02050_),
    .A1(net177),
    .A2(_03204_));
 sg13g2_nand2_1 _19046_ (.Y(_03234_),
    .A(\top_ihp.oisc.regs[57][7] ),
    .B(_03202_));
 sg13g2_o21ai_1 _19047_ (.B1(_03234_),
    .Y(_02051_),
    .A1(net47),
    .A2(_03204_));
 sg13g2_nand2_1 _19048_ (.Y(_03235_),
    .A(\top_ihp.oisc.regs[57][8] ),
    .B(net172));
 sg13g2_o21ai_1 _19049_ (.B1(_03235_),
    .Y(_02052_),
    .A1(net42),
    .A2(net171));
 sg13g2_nand2_1 _19050_ (.Y(_03236_),
    .A(\top_ihp.oisc.regs[57][9] ),
    .B(net172));
 sg13g2_o21ai_1 _19051_ (.B1(_03236_),
    .Y(_02053_),
    .A1(net25),
    .A2(net171));
 sg13g2_nor2_2 _19052_ (.A(_09956_),
    .B(_03050_),
    .Y(_03237_));
 sg13g2_mux2_1 _19053_ (.A0(\top_ihp.oisc.regs[58][0] ),
    .A1(_02845_),
    .S(_03237_),
    .X(_02054_));
 sg13g2_or2_1 _19054_ (.X(_03238_),
    .B(_03050_),
    .A(_09956_));
 sg13g2_buf_1 _19055_ (.A(_03238_),
    .X(_03239_));
 sg13g2_buf_1 _19056_ (.A(_03239_),
    .X(_03240_));
 sg13g2_buf_1 _19057_ (.A(net489),
    .X(_03241_));
 sg13g2_buf_2 _19058_ (.A(_03239_),
    .X(_03242_));
 sg13g2_nand2_1 _19059_ (.Y(_03243_),
    .A(\top_ihp.oisc.regs[58][10] ),
    .B(net488));
 sg13g2_o21ai_1 _19060_ (.B1(_03243_),
    .Y(_02055_),
    .A1(net26),
    .A2(_03241_));
 sg13g2_buf_1 _19061_ (.A(_03239_),
    .X(_03244_));
 sg13g2_nand2_1 _19062_ (.Y(_03245_),
    .A(\top_ihp.oisc.regs[58][11] ),
    .B(_03244_));
 sg13g2_o21ai_1 _19063_ (.B1(_03245_),
    .Y(_02056_),
    .A1(net89),
    .A2(_03241_));
 sg13g2_nand2_1 _19064_ (.Y(_03246_),
    .A(\top_ihp.oisc.regs[58][12] ),
    .B(net487));
 sg13g2_o21ai_1 _19065_ (.B1(_03246_),
    .Y(_02057_),
    .A1(net180),
    .A2(net308));
 sg13g2_nand2_1 _19066_ (.Y(_03247_),
    .A(\top_ihp.oisc.regs[58][13] ),
    .B(net487));
 sg13g2_o21ai_1 _19067_ (.B1(_03247_),
    .Y(_02058_),
    .A1(_10799_),
    .A2(net308));
 sg13g2_nand2_1 _19068_ (.Y(_03248_),
    .A(\top_ihp.oisc.regs[58][14] ),
    .B(net487));
 sg13g2_o21ai_1 _19069_ (.B1(_03248_),
    .Y(_02059_),
    .A1(net95),
    .A2(net308));
 sg13g2_nand2_1 _19070_ (.Y(_03249_),
    .A(\top_ihp.oisc.regs[58][15] ),
    .B(net487));
 sg13g2_o21ai_1 _19071_ (.B1(_03249_),
    .Y(_02060_),
    .A1(net176),
    .A2(net308));
 sg13g2_nand2_1 _19072_ (.Y(_03250_),
    .A(\top_ihp.oisc.regs[58][16] ),
    .B(net487));
 sg13g2_o21ai_1 _19073_ (.B1(_03250_),
    .Y(_02061_),
    .A1(net191),
    .A2(net308));
 sg13g2_nand2_1 _19074_ (.Y(_03251_),
    .A(\top_ihp.oisc.regs[58][17] ),
    .B(net487));
 sg13g2_o21ai_1 _19075_ (.B1(_03251_),
    .Y(_02062_),
    .A1(net94),
    .A2(net308));
 sg13g2_nand2_1 _19076_ (.Y(_03252_),
    .A(\top_ihp.oisc.regs[58][18] ),
    .B(net487));
 sg13g2_o21ai_1 _19077_ (.B1(_03252_),
    .Y(_02063_),
    .A1(net93),
    .A2(net308));
 sg13g2_nand2_1 _19078_ (.Y(_03253_),
    .A(\top_ihp.oisc.regs[58][19] ),
    .B(net487));
 sg13g2_o21ai_1 _19079_ (.B1(_03253_),
    .Y(_02064_),
    .A1(net92),
    .A2(net308));
 sg13g2_buf_1 _19080_ (.A(net489),
    .X(_03254_));
 sg13g2_nand2_1 _19081_ (.Y(_03255_),
    .A(\top_ihp.oisc.regs[58][1] ),
    .B(_03244_));
 sg13g2_o21ai_1 _19082_ (.B1(_03255_),
    .Y(_02065_),
    .A1(net496),
    .A2(net307));
 sg13g2_nor2_1 _19083_ (.A(\top_ihp.oisc.regs[58][20] ),
    .B(_03237_),
    .Y(_03256_));
 sg13g2_a21oi_1 _19084_ (.A1(net28),
    .A2(_03237_),
    .Y(_02066_),
    .B1(_03256_));
 sg13g2_buf_1 _19085_ (.A(_03239_),
    .X(_03257_));
 sg13g2_nand2_1 _19086_ (.Y(_03258_),
    .A(\top_ihp.oisc.regs[58][21] ),
    .B(net486));
 sg13g2_o21ai_1 _19087_ (.B1(_03258_),
    .Y(_02067_),
    .A1(net46),
    .A2(net307));
 sg13g2_nand2_1 _19088_ (.Y(_03259_),
    .A(\top_ihp.oisc.regs[58][22] ),
    .B(net486));
 sg13g2_o21ai_1 _19089_ (.B1(_03259_),
    .Y(_02068_),
    .A1(_10811_),
    .A2(net307));
 sg13g2_nor2_1 _19090_ (.A(\top_ihp.oisc.regs[58][23] ),
    .B(_03237_),
    .Y(_03260_));
 sg13g2_a21oi_1 _19091_ (.A1(_02697_),
    .A2(_03237_),
    .Y(_02069_),
    .B1(_03260_));
 sg13g2_nand2_1 _19092_ (.Y(_03261_),
    .A(\top_ihp.oisc.regs[58][24] ),
    .B(net486));
 sg13g2_o21ai_1 _19093_ (.B1(_03261_),
    .Y(_02070_),
    .A1(net91),
    .A2(net307));
 sg13g2_nand2_1 _19094_ (.Y(_03262_),
    .A(\top_ihp.oisc.regs[58][25] ),
    .B(net486));
 sg13g2_o21ai_1 _19095_ (.B1(_03262_),
    .Y(_02071_),
    .A1(net179),
    .A2(net307));
 sg13g2_nand2_1 _19096_ (.Y(_03263_),
    .A(\top_ihp.oisc.regs[58][26] ),
    .B(net486));
 sg13g2_o21ai_1 _19097_ (.B1(_03263_),
    .Y(_02072_),
    .A1(net90),
    .A2(net307));
 sg13g2_nand2_1 _19098_ (.Y(_03264_),
    .A(\top_ihp.oisc.regs[58][27] ),
    .B(net486));
 sg13g2_o21ai_1 _19099_ (.B1(_03264_),
    .Y(_02073_),
    .A1(net45),
    .A2(net307));
 sg13g2_nand2_1 _19100_ (.Y(_03265_),
    .A(\top_ihp.oisc.regs[58][28] ),
    .B(net486));
 sg13g2_o21ai_1 _19101_ (.B1(_03265_),
    .Y(_02074_),
    .A1(net44),
    .A2(net307));
 sg13g2_nand2_1 _19102_ (.Y(_03266_),
    .A(\top_ihp.oisc.regs[58][29] ),
    .B(_03257_));
 sg13g2_o21ai_1 _19103_ (.B1(_03266_),
    .Y(_02075_),
    .A1(net43),
    .A2(_03254_));
 sg13g2_nand2_1 _19104_ (.Y(_03267_),
    .A(\top_ihp.oisc.regs[58][2] ),
    .B(_03257_));
 sg13g2_o21ai_1 _19105_ (.B1(_03267_),
    .Y(_02076_),
    .A1(net175),
    .A2(_03254_));
 sg13g2_nand2_1 _19106_ (.Y(_03268_),
    .A(\top_ihp.oisc.regs[58][30] ),
    .B(net486));
 sg13g2_o21ai_1 _19107_ (.B1(_03268_),
    .Y(_02077_),
    .A1(_03145_),
    .A2(net488));
 sg13g2_nand2_1 _19108_ (.Y(_03269_),
    .A(\top_ihp.oisc.regs[58][31] ),
    .B(net489));
 sg13g2_o21ai_1 _19109_ (.B1(_03269_),
    .Y(_02078_),
    .A1(net87),
    .A2(_03242_));
 sg13g2_nand2_1 _19110_ (.Y(_03270_),
    .A(\top_ihp.oisc.regs[58][3] ),
    .B(net489));
 sg13g2_o21ai_1 _19111_ (.B1(_03270_),
    .Y(_02079_),
    .A1(net174),
    .A2(net488));
 sg13g2_nand2_1 _19112_ (.Y(_03271_),
    .A(\top_ihp.oisc.regs[58][4] ),
    .B(net489));
 sg13g2_o21ai_1 _19113_ (.B1(_03271_),
    .Y(_02080_),
    .A1(net88),
    .A2(net488));
 sg13g2_nand2_1 _19114_ (.Y(_03272_),
    .A(\top_ihp.oisc.regs[58][5] ),
    .B(_03240_));
 sg13g2_o21ai_1 _19115_ (.B1(_03272_),
    .Y(_02081_),
    .A1(net178),
    .A2(net488));
 sg13g2_nand2_1 _19116_ (.Y(_03273_),
    .A(\top_ihp.oisc.regs[58][6] ),
    .B(_03240_));
 sg13g2_o21ai_1 _19117_ (.B1(_03273_),
    .Y(_02082_),
    .A1(net177),
    .A2(net488));
 sg13g2_nand2_1 _19118_ (.Y(_03274_),
    .A(\top_ihp.oisc.regs[58][7] ),
    .B(net489));
 sg13g2_o21ai_1 _19119_ (.B1(_03274_),
    .Y(_02083_),
    .A1(net47),
    .A2(_03242_));
 sg13g2_nand2_1 _19120_ (.Y(_03275_),
    .A(\top_ihp.oisc.regs[58][8] ),
    .B(net489));
 sg13g2_o21ai_1 _19121_ (.B1(_03275_),
    .Y(_02084_),
    .A1(net42),
    .A2(net488));
 sg13g2_nand2_1 _19122_ (.Y(_03276_),
    .A(\top_ihp.oisc.regs[58][9] ),
    .B(net489));
 sg13g2_o21ai_1 _19123_ (.B1(_03276_),
    .Y(_02085_),
    .A1(net25),
    .A2(net488));
 sg13g2_or2_1 _19124_ (.X(_03277_),
    .B(_03110_),
    .A(_09958_));
 sg13g2_buf_2 _19125_ (.A(_03277_),
    .X(_03278_));
 sg13g2_buf_1 _19126_ (.A(_03278_),
    .X(_03279_));
 sg13g2_mux2_1 _19127_ (.A0(_09946_),
    .A1(\top_ihp.oisc.regs[59][0] ),
    .S(_03279_),
    .X(_02086_));
 sg13g2_buf_1 _19128_ (.A(_03278_),
    .X(_03280_));
 sg13g2_nand2_1 _19129_ (.Y(_03281_),
    .A(\top_ihp.oisc.regs[59][10] ),
    .B(net168));
 sg13g2_o21ai_1 _19130_ (.B1(_03281_),
    .Y(_02087_),
    .A1(net26),
    .A2(_03280_));
 sg13g2_nand2_1 _19131_ (.Y(_03282_),
    .A(\top_ihp.oisc.regs[59][11] ),
    .B(net168));
 sg13g2_o21ai_1 _19132_ (.B1(_03282_),
    .Y(_02088_),
    .A1(net89),
    .A2(net167));
 sg13g2_nand2_1 _19133_ (.Y(_03283_),
    .A(\top_ihp.oisc.regs[59][12] ),
    .B(net168));
 sg13g2_o21ai_1 _19134_ (.B1(_03283_),
    .Y(_02089_),
    .A1(net180),
    .A2(net167));
 sg13g2_nand2_1 _19135_ (.Y(_03284_),
    .A(\top_ihp.oisc.regs[59][13] ),
    .B(net168));
 sg13g2_o21ai_1 _19136_ (.B1(_03284_),
    .Y(_02090_),
    .A1(net147),
    .A2(net167));
 sg13g2_nand2_1 _19137_ (.Y(_03285_),
    .A(\top_ihp.oisc.regs[59][14] ),
    .B(net168));
 sg13g2_o21ai_1 _19138_ (.B1(_03285_),
    .Y(_02091_),
    .A1(_03065_),
    .A2(_03280_));
 sg13g2_nand2_1 _19139_ (.Y(_03286_),
    .A(\top_ihp.oisc.regs[59][15] ),
    .B(net168));
 sg13g2_o21ai_1 _19140_ (.B1(_03286_),
    .Y(_02092_),
    .A1(_03123_),
    .A2(net167));
 sg13g2_nand2_1 _19141_ (.Y(_03287_),
    .A(\top_ihp.oisc.regs[59][16] ),
    .B(_03279_));
 sg13g2_o21ai_1 _19142_ (.B1(_03287_),
    .Y(_02093_),
    .A1(net247),
    .A2(net167));
 sg13g2_nand2_1 _19143_ (.Y(_03288_),
    .A(\top_ihp.oisc.regs[59][17] ),
    .B(net168));
 sg13g2_o21ai_1 _19144_ (.B1(_03288_),
    .Y(_02094_),
    .A1(net94),
    .A2(net167));
 sg13g2_buf_1 _19145_ (.A(_03278_),
    .X(_03289_));
 sg13g2_nand2_1 _19146_ (.Y(_03290_),
    .A(\top_ihp.oisc.regs[59][18] ),
    .B(net166));
 sg13g2_o21ai_1 _19147_ (.B1(_03290_),
    .Y(_02095_),
    .A1(net93),
    .A2(net167));
 sg13g2_nand2_1 _19148_ (.Y(_03291_),
    .A(\top_ihp.oisc.regs[59][19] ),
    .B(net166));
 sg13g2_o21ai_1 _19149_ (.B1(_03291_),
    .Y(_02096_),
    .A1(net92),
    .A2(net167));
 sg13g2_buf_1 _19150_ (.A(_03278_),
    .X(_03292_));
 sg13g2_nand2_1 _19151_ (.Y(_03293_),
    .A(\top_ihp.oisc.regs[59][1] ),
    .B(net166));
 sg13g2_o21ai_1 _19152_ (.B1(_03293_),
    .Y(_02097_),
    .A1(net496),
    .A2(net165));
 sg13g2_nand2_1 _19153_ (.Y(_03294_),
    .A(\top_ihp.oisc.regs[59][20] ),
    .B(net166));
 sg13g2_o21ai_1 _19154_ (.B1(_03294_),
    .Y(_02098_),
    .A1(_09581_),
    .A2(net165));
 sg13g2_nand2_1 _19155_ (.Y(_03295_),
    .A(\top_ihp.oisc.regs[59][21] ),
    .B(net166));
 sg13g2_o21ai_1 _19156_ (.B1(_03295_),
    .Y(_02099_),
    .A1(net46),
    .A2(net165));
 sg13g2_nand2_1 _19157_ (.Y(_03296_),
    .A(\top_ihp.oisc.regs[59][22] ),
    .B(net166));
 sg13g2_o21ai_1 _19158_ (.B1(_03296_),
    .Y(_02100_),
    .A1(net244),
    .A2(net165));
 sg13g2_mux2_1 _19159_ (.A0(net224),
    .A1(\top_ihp.oisc.regs[59][23] ),
    .S(net168),
    .X(_02101_));
 sg13g2_nand2_1 _19160_ (.Y(_03297_),
    .A(\top_ihp.oisc.regs[59][24] ),
    .B(net166));
 sg13g2_o21ai_1 _19161_ (.B1(_03297_),
    .Y(_02102_),
    .A1(net91),
    .A2(net165));
 sg13g2_nand2_1 _19162_ (.Y(_03298_),
    .A(\top_ihp.oisc.regs[59][25] ),
    .B(net166));
 sg13g2_o21ai_1 _19163_ (.B1(_03298_),
    .Y(_02103_),
    .A1(net179),
    .A2(net165));
 sg13g2_nand2_1 _19164_ (.Y(_03299_),
    .A(\top_ihp.oisc.regs[59][26] ),
    .B(_03289_));
 sg13g2_o21ai_1 _19165_ (.B1(_03299_),
    .Y(_02104_),
    .A1(_03088_),
    .A2(net165));
 sg13g2_nand2_1 _19166_ (.Y(_03300_),
    .A(\top_ihp.oisc.regs[59][27] ),
    .B(_03289_));
 sg13g2_o21ai_1 _19167_ (.B1(_03300_),
    .Y(_02105_),
    .A1(net45),
    .A2(_03292_));
 sg13g2_buf_1 _19168_ (.A(_03278_),
    .X(_03301_));
 sg13g2_nand2_1 _19169_ (.Y(_03302_),
    .A(\top_ihp.oisc.regs[59][28] ),
    .B(net164));
 sg13g2_o21ai_1 _19170_ (.B1(_03302_),
    .Y(_02106_),
    .A1(net44),
    .A2(_03292_));
 sg13g2_nand2_1 _19171_ (.Y(_03303_),
    .A(\top_ihp.oisc.regs[59][29] ),
    .B(_03301_));
 sg13g2_o21ai_1 _19172_ (.B1(_03303_),
    .Y(_02107_),
    .A1(net43),
    .A2(net165));
 sg13g2_buf_1 _19173_ (.A(_03278_),
    .X(_03304_));
 sg13g2_nand2_1 _19174_ (.Y(_03305_),
    .A(\top_ihp.oisc.regs[59][2] ),
    .B(net164));
 sg13g2_o21ai_1 _19175_ (.B1(_03305_),
    .Y(_02108_),
    .A1(net175),
    .A2(net163));
 sg13g2_nand2_1 _19176_ (.Y(_03306_),
    .A(\top_ihp.oisc.regs[59][30] ),
    .B(net164));
 sg13g2_o21ai_1 _19177_ (.B1(_03306_),
    .Y(_02109_),
    .A1(net41),
    .A2(net163));
 sg13g2_nand2_1 _19178_ (.Y(_03307_),
    .A(\top_ihp.oisc.regs[59][31] ),
    .B(net164));
 sg13g2_o21ai_1 _19179_ (.B1(_03307_),
    .Y(_02110_),
    .A1(net87),
    .A2(_03304_));
 sg13g2_nand2_1 _19180_ (.Y(_03308_),
    .A(\top_ihp.oisc.regs[59][3] ),
    .B(_03301_));
 sg13g2_o21ai_1 _19181_ (.B1(_03308_),
    .Y(_02111_),
    .A1(net174),
    .A2(net163));
 sg13g2_nand2_1 _19182_ (.Y(_03309_),
    .A(\top_ihp.oisc.regs[59][4] ),
    .B(net164));
 sg13g2_o21ai_1 _19183_ (.B1(_03309_),
    .Y(_02112_),
    .A1(net88),
    .A2(net163));
 sg13g2_nand2_1 _19184_ (.Y(_03310_),
    .A(\top_ihp.oisc.regs[59][5] ),
    .B(net164));
 sg13g2_o21ai_1 _19185_ (.B1(_03310_),
    .Y(_02113_),
    .A1(net178),
    .A2(net163));
 sg13g2_nand2_1 _19186_ (.Y(_03311_),
    .A(\top_ihp.oisc.regs[59][6] ),
    .B(net164));
 sg13g2_o21ai_1 _19187_ (.B1(_03311_),
    .Y(_02114_),
    .A1(net177),
    .A2(net163));
 sg13g2_nand2_1 _19188_ (.Y(_03312_),
    .A(\top_ihp.oisc.regs[59][7] ),
    .B(net164));
 sg13g2_o21ai_1 _19189_ (.B1(_03312_),
    .Y(_02115_),
    .A1(_02718_),
    .A2(_03304_));
 sg13g2_nand2_1 _19190_ (.Y(_03313_),
    .A(\top_ihp.oisc.regs[59][8] ),
    .B(_03278_));
 sg13g2_o21ai_1 _19191_ (.B1(_03313_),
    .Y(_02116_),
    .A1(net42),
    .A2(net163));
 sg13g2_nand2_1 _19192_ (.Y(_03314_),
    .A(\top_ihp.oisc.regs[59][9] ),
    .B(_03278_));
 sg13g2_o21ai_1 _19193_ (.B1(_03314_),
    .Y(_02117_),
    .A1(net25),
    .A2(net163));
 sg13g2_nor2_1 _19194_ (.A(_10093_),
    .B(net682),
    .Y(_03315_));
 sg13g2_buf_1 _19195_ (.A(_03315_),
    .X(_03316_));
 sg13g2_mux2_1 _19196_ (.A0(\top_ihp.oisc.regs[5][0] ),
    .A1(net334),
    .S(net630),
    .X(_02118_));
 sg13g2_inv_1 _19197_ (.Y(_03317_),
    .A(_10093_));
 sg13g2_nand2_1 _19198_ (.Y(_03318_),
    .A(_03317_),
    .B(net663));
 sg13g2_buf_1 _19199_ (.A(_03318_),
    .X(_03319_));
 sg13g2_buf_1 _19200_ (.A(net485),
    .X(_03320_));
 sg13g2_buf_1 _19201_ (.A(net485),
    .X(_03321_));
 sg13g2_nand2_1 _19202_ (.Y(_03322_),
    .A(\top_ihp.oisc.regs[5][10] ),
    .B(net305));
 sg13g2_o21ai_1 _19203_ (.B1(_03322_),
    .Y(_02119_),
    .A1(_03053_),
    .A2(net306));
 sg13g2_nand2_1 _19204_ (.Y(_03323_),
    .A(\top_ihp.oisc.regs[5][11] ),
    .B(net305));
 sg13g2_o21ai_1 _19205_ (.B1(_03323_),
    .Y(_02120_),
    .A1(net89),
    .A2(net306));
 sg13g2_nand2_1 _19206_ (.Y(_03324_),
    .A(\top_ihp.oisc.regs[5][12] ),
    .B(_03321_));
 sg13g2_o21ai_1 _19207_ (.B1(_03324_),
    .Y(_02121_),
    .A1(_03061_),
    .A2(net306));
 sg13g2_nor2_1 _19208_ (.A(\top_ihp.oisc.regs[5][13] ),
    .B(net630),
    .Y(_03325_));
 sg13g2_a21oi_1 _19209_ (.A1(net73),
    .A2(net630),
    .Y(_02122_),
    .B1(_03325_));
 sg13g2_buf_1 _19210_ (.A(net485),
    .X(_03326_));
 sg13g2_nand2_1 _19211_ (.Y(_03327_),
    .A(\top_ihp.oisc.regs[5][14] ),
    .B(net304));
 sg13g2_o21ai_1 _19212_ (.B1(_03327_),
    .Y(_02123_),
    .A1(net95),
    .A2(net306));
 sg13g2_nand2_1 _19213_ (.Y(_03328_),
    .A(\top_ihp.oisc.regs[5][15] ),
    .B(net304));
 sg13g2_o21ai_1 _19214_ (.B1(_03328_),
    .Y(_02124_),
    .A1(net176),
    .A2(net306));
 sg13g2_nor2_1 _19215_ (.A(\top_ihp.oisc.regs[5][16] ),
    .B(net630),
    .Y(_03329_));
 sg13g2_a21oi_1 _19216_ (.A1(net146),
    .A2(net630),
    .Y(_02125_),
    .B1(_03329_));
 sg13g2_nand2_1 _19217_ (.Y(_03330_),
    .A(\top_ihp.oisc.regs[5][17] ),
    .B(net304));
 sg13g2_o21ai_1 _19218_ (.B1(_03330_),
    .Y(_02126_),
    .A1(net94),
    .A2(net306));
 sg13g2_nand2_1 _19219_ (.Y(_03331_),
    .A(\top_ihp.oisc.regs[5][18] ),
    .B(net304));
 sg13g2_o21ai_1 _19220_ (.B1(_03331_),
    .Y(_02127_),
    .A1(_03071_),
    .A2(_03320_));
 sg13g2_nand2_1 _19221_ (.Y(_03332_),
    .A(\top_ihp.oisc.regs[5][19] ),
    .B(net304));
 sg13g2_o21ai_1 _19222_ (.B1(_03332_),
    .Y(_02128_),
    .A1(net92),
    .A2(net306));
 sg13g2_nand2_1 _19223_ (.Y(_03333_),
    .A(\top_ihp.oisc.regs[5][1] ),
    .B(_03326_));
 sg13g2_o21ai_1 _19224_ (.B1(_03333_),
    .Y(_02129_),
    .A1(_03075_),
    .A2(_03320_));
 sg13g2_nand2_1 _19225_ (.Y(_03334_),
    .A(\top_ihp.oisc.regs[5][20] ),
    .B(net304));
 sg13g2_o21ai_1 _19226_ (.B1(_03334_),
    .Y(_02130_),
    .A1(_09563_),
    .A2(net306));
 sg13g2_buf_1 _19227_ (.A(net485),
    .X(_03335_));
 sg13g2_nand2_1 _19228_ (.Y(_03336_),
    .A(\top_ihp.oisc.regs[5][21] ),
    .B(net304));
 sg13g2_o21ai_1 _19229_ (.B1(_03336_),
    .Y(_02131_),
    .A1(_03078_),
    .A2(net303));
 sg13g2_nor2_1 _19230_ (.A(\top_ihp.oisc.regs[5][22] ),
    .B(_03316_),
    .Y(_03337_));
 sg13g2_a21oi_1 _19231_ (.A1(net143),
    .A2(net630),
    .Y(_02132_),
    .B1(_03337_));
 sg13g2_nor2_1 _19232_ (.A(\top_ihp.oisc.regs[5][23] ),
    .B(net630),
    .Y(_03338_));
 sg13g2_a21oi_1 _19233_ (.A1(net100),
    .A2(net630),
    .Y(_02133_),
    .B1(_03338_));
 sg13g2_nand2_1 _19234_ (.Y(_03339_),
    .A(\top_ihp.oisc.regs[5][24] ),
    .B(_03326_));
 sg13g2_o21ai_1 _19235_ (.B1(_03339_),
    .Y(_02134_),
    .A1(net91),
    .A2(_03335_));
 sg13g2_nand2_1 _19236_ (.Y(_03340_),
    .A(\top_ihp.oisc.regs[5][25] ),
    .B(net304));
 sg13g2_o21ai_1 _19237_ (.B1(_03340_),
    .Y(_02135_),
    .A1(_03086_),
    .A2(net303));
 sg13g2_buf_1 _19238_ (.A(_03319_),
    .X(_03341_));
 sg13g2_nand2_1 _19239_ (.Y(_03342_),
    .A(\top_ihp.oisc.regs[5][26] ),
    .B(net302));
 sg13g2_o21ai_1 _19240_ (.B1(_03342_),
    .Y(_02136_),
    .A1(_03088_),
    .A2(_03335_));
 sg13g2_nand2_1 _19241_ (.Y(_03343_),
    .A(\top_ihp.oisc.regs[5][27] ),
    .B(net302));
 sg13g2_o21ai_1 _19242_ (.B1(_03343_),
    .Y(_02137_),
    .A1(_03090_),
    .A2(net303));
 sg13g2_nand2_1 _19243_ (.Y(_03344_),
    .A(\top_ihp.oisc.regs[5][28] ),
    .B(net302));
 sg13g2_o21ai_1 _19244_ (.B1(_03344_),
    .Y(_02138_),
    .A1(_03092_),
    .A2(net303));
 sg13g2_nand2_1 _19245_ (.Y(_03345_),
    .A(\top_ihp.oisc.regs[5][29] ),
    .B(_03341_));
 sg13g2_o21ai_1 _19246_ (.B1(_03345_),
    .Y(_02139_),
    .A1(_03094_),
    .A2(net303));
 sg13g2_nand2_1 _19247_ (.Y(_03346_),
    .A(\top_ihp.oisc.regs[5][2] ),
    .B(net302));
 sg13g2_o21ai_1 _19248_ (.B1(_03346_),
    .Y(_02140_),
    .A1(_03143_),
    .A2(net303));
 sg13g2_nand2_1 _19249_ (.Y(_03347_),
    .A(\top_ihp.oisc.regs[5][30] ),
    .B(_03341_));
 sg13g2_o21ai_1 _19250_ (.B1(_03347_),
    .Y(_02141_),
    .A1(net41),
    .A2(net303));
 sg13g2_nand2_1 _19251_ (.Y(_03348_),
    .A(\top_ihp.oisc.regs[5][31] ),
    .B(net302));
 sg13g2_o21ai_1 _19252_ (.B1(_03348_),
    .Y(_02142_),
    .A1(net87),
    .A2(net303));
 sg13g2_nand2_1 _19253_ (.Y(_03349_),
    .A(\top_ihp.oisc.regs[5][3] ),
    .B(net302));
 sg13g2_o21ai_1 _19254_ (.B1(_03349_),
    .Y(_02143_),
    .A1(_03148_),
    .A2(net305));
 sg13g2_nand2_1 _19255_ (.Y(_03350_),
    .A(\top_ihp.oisc.regs[5][4] ),
    .B(net302));
 sg13g2_o21ai_1 _19256_ (.B1(_03350_),
    .Y(_02144_),
    .A1(_03150_),
    .A2(net305));
 sg13g2_nand2_1 _19257_ (.Y(_03351_),
    .A(\top_ihp.oisc.regs[5][5] ),
    .B(net302));
 sg13g2_o21ai_1 _19258_ (.B1(_03351_),
    .Y(_02145_),
    .A1(net178),
    .A2(net305));
 sg13g2_nand2_1 _19259_ (.Y(_03352_),
    .A(\top_ihp.oisc.regs[5][6] ),
    .B(net485));
 sg13g2_o21ai_1 _19260_ (.B1(_03352_),
    .Y(_02146_),
    .A1(_03103_),
    .A2(net305));
 sg13g2_nand2_1 _19261_ (.Y(_03353_),
    .A(\top_ihp.oisc.regs[5][7] ),
    .B(net485));
 sg13g2_o21ai_1 _19262_ (.B1(_03353_),
    .Y(_02147_),
    .A1(_02666_),
    .A2(net305));
 sg13g2_nand2_1 _19263_ (.Y(_03354_),
    .A(\top_ihp.oisc.regs[5][8] ),
    .B(net485));
 sg13g2_o21ai_1 _19264_ (.B1(_03354_),
    .Y(_02148_),
    .A1(_03106_),
    .A2(_03321_));
 sg13g2_nand2_1 _19265_ (.Y(_03355_),
    .A(\top_ihp.oisc.regs[5][9] ),
    .B(net485));
 sg13g2_o21ai_1 _19266_ (.B1(_03355_),
    .Y(_02149_),
    .A1(_03108_),
    .A2(net305));
 sg13g2_and2_1 _19267_ (.A(net665),
    .B(_02968_),
    .X(_03356_));
 sg13g2_buf_1 _19268_ (.A(_03356_),
    .X(_03357_));
 sg13g2_mux2_1 _19269_ (.A0(\top_ihp.oisc.regs[60][0] ),
    .A1(net412),
    .S(_03357_),
    .X(_02150_));
 sg13g2_nand2_1 _19270_ (.Y(_03358_),
    .A(_10055_),
    .B(_02968_));
 sg13g2_buf_1 _19271_ (.A(_03358_),
    .X(_03359_));
 sg13g2_buf_1 _19272_ (.A(_03359_),
    .X(_03360_));
 sg13g2_buf_1 _19273_ (.A(net301),
    .X(_03361_));
 sg13g2_buf_1 _19274_ (.A(_03359_),
    .X(_03362_));
 sg13g2_nand2_1 _19275_ (.Y(_03363_),
    .A(\top_ihp.oisc.regs[60][10] ),
    .B(net300));
 sg13g2_o21ai_1 _19276_ (.B1(_03363_),
    .Y(_02151_),
    .A1(net26),
    .A2(_03361_));
 sg13g2_buf_1 _19277_ (.A(_03359_),
    .X(_03364_));
 sg13g2_nand2_1 _19278_ (.Y(_03365_),
    .A(\top_ihp.oisc.regs[60][11] ),
    .B(net299));
 sg13g2_o21ai_1 _19279_ (.B1(_03365_),
    .Y(_02152_),
    .A1(_03118_),
    .A2(net162));
 sg13g2_nand2_1 _19280_ (.Y(_03366_),
    .A(\top_ihp.oisc.regs[60][12] ),
    .B(_03364_));
 sg13g2_o21ai_1 _19281_ (.B1(_03366_),
    .Y(_02153_),
    .A1(net180),
    .A2(_03361_));
 sg13g2_nand2_1 _19282_ (.Y(_03367_),
    .A(\top_ihp.oisc.regs[60][13] ),
    .B(net299));
 sg13g2_o21ai_1 _19283_ (.B1(_03367_),
    .Y(_02154_),
    .A1(net147),
    .A2(net162));
 sg13g2_nand2_1 _19284_ (.Y(_03368_),
    .A(\top_ihp.oisc.regs[60][14] ),
    .B(net299));
 sg13g2_o21ai_1 _19285_ (.B1(_03368_),
    .Y(_02155_),
    .A1(net95),
    .A2(net162));
 sg13g2_nand2_1 _19286_ (.Y(_03369_),
    .A(\top_ihp.oisc.regs[60][15] ),
    .B(net299));
 sg13g2_o21ai_1 _19287_ (.B1(_03369_),
    .Y(_02156_),
    .A1(net176),
    .A2(net162));
 sg13g2_nand2_1 _19288_ (.Y(_03370_),
    .A(\top_ihp.oisc.regs[60][16] ),
    .B(net299));
 sg13g2_o21ai_1 _19289_ (.B1(_03370_),
    .Y(_02157_),
    .A1(net247),
    .A2(net162));
 sg13g2_nand2_1 _19290_ (.Y(_03371_),
    .A(\top_ihp.oisc.regs[60][17] ),
    .B(net299));
 sg13g2_o21ai_1 _19291_ (.B1(_03371_),
    .Y(_02158_),
    .A1(net94),
    .A2(net162));
 sg13g2_nand2_1 _19292_ (.Y(_03372_),
    .A(\top_ihp.oisc.regs[60][18] ),
    .B(net299));
 sg13g2_o21ai_1 _19293_ (.B1(_03372_),
    .Y(_02159_),
    .A1(net93),
    .A2(net162));
 sg13g2_nand2_1 _19294_ (.Y(_03373_),
    .A(\top_ihp.oisc.regs[60][19] ),
    .B(net299));
 sg13g2_o21ai_1 _19295_ (.B1(_03373_),
    .Y(_02160_),
    .A1(net92),
    .A2(net162));
 sg13g2_buf_1 _19296_ (.A(_03360_),
    .X(_03374_));
 sg13g2_nand2_1 _19297_ (.Y(_03375_),
    .A(\top_ihp.oisc.regs[60][1] ),
    .B(_03364_));
 sg13g2_o21ai_1 _19298_ (.B1(_03375_),
    .Y(_02161_),
    .A1(net496),
    .A2(net161));
 sg13g2_mux2_1 _19299_ (.A0(\top_ihp.oisc.regs[60][20] ),
    .A1(net245),
    .S(_03357_),
    .X(_02162_));
 sg13g2_buf_1 _19300_ (.A(_03359_),
    .X(_03376_));
 sg13g2_nand2_1 _19301_ (.Y(_03377_),
    .A(\top_ihp.oisc.regs[60][21] ),
    .B(net298));
 sg13g2_o21ai_1 _19302_ (.B1(_03377_),
    .Y(_02163_),
    .A1(net46),
    .A2(net161));
 sg13g2_nand2_1 _19303_ (.Y(_03378_),
    .A(\top_ihp.oisc.regs[60][22] ),
    .B(net298));
 sg13g2_o21ai_1 _19304_ (.B1(_03378_),
    .Y(_02164_),
    .A1(_09622_),
    .A2(net161));
 sg13g2_mux2_1 _19305_ (.A0(\top_ihp.oisc.regs[60][23] ),
    .A1(_10035_),
    .S(_03357_),
    .X(_02165_));
 sg13g2_nand2_1 _19306_ (.Y(_03379_),
    .A(\top_ihp.oisc.regs[60][24] ),
    .B(net298));
 sg13g2_o21ai_1 _19307_ (.B1(_03379_),
    .Y(_02166_),
    .A1(net91),
    .A2(net161));
 sg13g2_nand2_1 _19308_ (.Y(_03380_),
    .A(\top_ihp.oisc.regs[60][25] ),
    .B(net298));
 sg13g2_o21ai_1 _19309_ (.B1(_03380_),
    .Y(_02167_),
    .A1(net179),
    .A2(net161));
 sg13g2_nand2_1 _19310_ (.Y(_03381_),
    .A(\top_ihp.oisc.regs[60][26] ),
    .B(net298));
 sg13g2_o21ai_1 _19311_ (.B1(_03381_),
    .Y(_02168_),
    .A1(net90),
    .A2(net161));
 sg13g2_nand2_1 _19312_ (.Y(_03382_),
    .A(\top_ihp.oisc.regs[60][27] ),
    .B(_03376_));
 sg13g2_o21ai_1 _19313_ (.B1(_03382_),
    .Y(_02169_),
    .A1(net45),
    .A2(net161));
 sg13g2_nand2_1 _19314_ (.Y(_03383_),
    .A(\top_ihp.oisc.regs[60][28] ),
    .B(net298));
 sg13g2_o21ai_1 _19315_ (.B1(_03383_),
    .Y(_02170_),
    .A1(net44),
    .A2(net161));
 sg13g2_nand2_1 _19316_ (.Y(_03384_),
    .A(\top_ihp.oisc.regs[60][29] ),
    .B(net298));
 sg13g2_o21ai_1 _19317_ (.B1(_03384_),
    .Y(_02171_),
    .A1(net43),
    .A2(_03374_));
 sg13g2_nand2_1 _19318_ (.Y(_03385_),
    .A(\top_ihp.oisc.regs[60][2] ),
    .B(_03376_));
 sg13g2_o21ai_1 _19319_ (.B1(_03385_),
    .Y(_02172_),
    .A1(_03143_),
    .A2(_03374_));
 sg13g2_nand2_1 _19320_ (.Y(_03386_),
    .A(\top_ihp.oisc.regs[60][30] ),
    .B(net298));
 sg13g2_o21ai_1 _19321_ (.B1(_03386_),
    .Y(_02173_),
    .A1(net41),
    .A2(_03362_));
 sg13g2_nand2_1 _19322_ (.Y(_03387_),
    .A(\top_ihp.oisc.regs[60][31] ),
    .B(net301));
 sg13g2_o21ai_1 _19323_ (.B1(_03387_),
    .Y(_02174_),
    .A1(net87),
    .A2(net300));
 sg13g2_nand2_1 _19324_ (.Y(_03388_),
    .A(\top_ihp.oisc.regs[60][3] ),
    .B(_03360_));
 sg13g2_o21ai_1 _19325_ (.B1(_03388_),
    .Y(_02175_),
    .A1(net174),
    .A2(_03362_));
 sg13g2_nand2_1 _19326_ (.Y(_03389_),
    .A(\top_ihp.oisc.regs[60][4] ),
    .B(net301));
 sg13g2_o21ai_1 _19327_ (.B1(_03389_),
    .Y(_02176_),
    .A1(net88),
    .A2(net300));
 sg13g2_nand2_1 _19328_ (.Y(_03390_),
    .A(\top_ihp.oisc.regs[60][5] ),
    .B(net301));
 sg13g2_o21ai_1 _19329_ (.B1(_03390_),
    .Y(_02177_),
    .A1(net178),
    .A2(net300));
 sg13g2_nand2_1 _19330_ (.Y(_03391_),
    .A(\top_ihp.oisc.regs[60][6] ),
    .B(net301));
 sg13g2_o21ai_1 _19331_ (.B1(_03391_),
    .Y(_02178_),
    .A1(_03103_),
    .A2(net300));
 sg13g2_nand2_1 _19332_ (.Y(_03392_),
    .A(\top_ihp.oisc.regs[60][7] ),
    .B(net301));
 sg13g2_o21ai_1 _19333_ (.B1(_03392_),
    .Y(_02179_),
    .A1(net408),
    .A2(net300));
 sg13g2_nand2_1 _19334_ (.Y(_03393_),
    .A(\top_ihp.oisc.regs[60][8] ),
    .B(net301));
 sg13g2_o21ai_1 _19335_ (.B1(_03393_),
    .Y(_02180_),
    .A1(net42),
    .A2(net300));
 sg13g2_nand2_1 _19336_ (.Y(_03394_),
    .A(\top_ihp.oisc.regs[60][9] ),
    .B(net301));
 sg13g2_o21ai_1 _19337_ (.B1(_03394_),
    .Y(_02181_),
    .A1(net25),
    .A2(net300));
 sg13g2_nor2_1 _19338_ (.A(_10090_),
    .B(_03009_),
    .Y(_03395_));
 sg13g2_buf_1 _19339_ (.A(_03395_),
    .X(_03396_));
 sg13g2_mux2_1 _19340_ (.A0(\top_ihp.oisc.regs[61][0] ),
    .A1(net412),
    .S(net484),
    .X(_02182_));
 sg13g2_nand3_1 _19341_ (.B(_10092_),
    .C(_02763_),
    .A(_10151_),
    .Y(_03397_));
 sg13g2_buf_2 _19342_ (.A(_03397_),
    .X(_03398_));
 sg13g2_buf_1 _19343_ (.A(_03398_),
    .X(_03399_));
 sg13g2_buf_1 _19344_ (.A(_03398_),
    .X(_03400_));
 sg13g2_nand2_1 _19345_ (.Y(_03401_),
    .A(\top_ihp.oisc.regs[61][10] ),
    .B(net296));
 sg13g2_o21ai_1 _19346_ (.B1(_03401_),
    .Y(_02183_),
    .A1(_03053_),
    .A2(_03399_));
 sg13g2_nand2_1 _19347_ (.Y(_03402_),
    .A(\top_ihp.oisc.regs[61][11] ),
    .B(net296));
 sg13g2_o21ai_1 _19348_ (.B1(_03402_),
    .Y(_02184_),
    .A1(_03118_),
    .A2(net297));
 sg13g2_nand2_1 _19349_ (.Y(_03403_),
    .A(\top_ihp.oisc.regs[61][12] ),
    .B(net296));
 sg13g2_o21ai_1 _19350_ (.B1(_03403_),
    .Y(_02185_),
    .A1(net180),
    .A2(_03399_));
 sg13g2_nor2_1 _19351_ (.A(\top_ihp.oisc.regs[61][13] ),
    .B(net484),
    .Y(_03404_));
 sg13g2_a21oi_1 _19352_ (.A1(_09375_),
    .A2(net484),
    .Y(_02186_),
    .B1(_03404_));
 sg13g2_nand2_1 _19353_ (.Y(_03405_),
    .A(\top_ihp.oisc.regs[61][14] ),
    .B(net296));
 sg13g2_o21ai_1 _19354_ (.B1(_03405_),
    .Y(_02187_),
    .A1(net95),
    .A2(net297));
 sg13g2_buf_1 _19355_ (.A(_03398_),
    .X(_03406_));
 sg13g2_nand2_1 _19356_ (.Y(_03407_),
    .A(\top_ihp.oisc.regs[61][15] ),
    .B(net295));
 sg13g2_o21ai_1 _19357_ (.B1(_03407_),
    .Y(_02188_),
    .A1(net176),
    .A2(net297));
 sg13g2_nor2_1 _19358_ (.A(\top_ihp.oisc.regs[61][16] ),
    .B(net484),
    .Y(_03408_));
 sg13g2_a21oi_1 _19359_ (.A1(_09437_),
    .A2(net484),
    .Y(_02189_),
    .B1(_03408_));
 sg13g2_nand2_1 _19360_ (.Y(_03409_),
    .A(\top_ihp.oisc.regs[61][17] ),
    .B(net295));
 sg13g2_o21ai_1 _19361_ (.B1(_03409_),
    .Y(_02190_),
    .A1(_03069_),
    .A2(net297));
 sg13g2_nand2_1 _19362_ (.Y(_03410_),
    .A(\top_ihp.oisc.regs[61][18] ),
    .B(net295));
 sg13g2_o21ai_1 _19363_ (.B1(_03410_),
    .Y(_02191_),
    .A1(net93),
    .A2(net297));
 sg13g2_nand2_1 _19364_ (.Y(_03411_),
    .A(\top_ihp.oisc.regs[61][19] ),
    .B(net295));
 sg13g2_o21ai_1 _19365_ (.B1(_03411_),
    .Y(_02192_),
    .A1(net92),
    .A2(net297));
 sg13g2_nand2_1 _19366_ (.Y(_03412_),
    .A(\top_ihp.oisc.regs[61][1] ),
    .B(net295));
 sg13g2_o21ai_1 _19367_ (.B1(_03412_),
    .Y(_02193_),
    .A1(net496),
    .A2(net297));
 sg13g2_nor2_1 _19368_ (.A(\top_ihp.oisc.regs[61][20] ),
    .B(_03396_),
    .Y(_03413_));
 sg13g2_a21oi_1 _19369_ (.A1(net28),
    .A2(_03396_),
    .Y(_02194_),
    .B1(_03413_));
 sg13g2_nand2_1 _19370_ (.Y(_03414_),
    .A(\top_ihp.oisc.regs[61][21] ),
    .B(net295));
 sg13g2_o21ai_1 _19371_ (.B1(_03414_),
    .Y(_02195_),
    .A1(net46),
    .A2(net297));
 sg13g2_nor2_1 _19372_ (.A(\top_ihp.oisc.regs[61][22] ),
    .B(net484),
    .Y(_03415_));
 sg13g2_a21oi_1 _19373_ (.A1(_09623_),
    .A2(net484),
    .Y(_02196_),
    .B1(_03415_));
 sg13g2_nor2_1 _19374_ (.A(\top_ihp.oisc.regs[61][23] ),
    .B(_03395_),
    .Y(_03416_));
 sg13g2_a21oi_1 _19375_ (.A1(_09643_),
    .A2(net484),
    .Y(_02197_),
    .B1(_03416_));
 sg13g2_buf_1 _19376_ (.A(_03398_),
    .X(_03417_));
 sg13g2_nand2_1 _19377_ (.Y(_03418_),
    .A(\top_ihp.oisc.regs[61][24] ),
    .B(net295));
 sg13g2_o21ai_1 _19378_ (.B1(_03418_),
    .Y(_02198_),
    .A1(net91),
    .A2(net294));
 sg13g2_nand2_1 _19379_ (.Y(_03419_),
    .A(\top_ihp.oisc.regs[61][25] ),
    .B(net295));
 sg13g2_o21ai_1 _19380_ (.B1(_03419_),
    .Y(_02199_),
    .A1(net179),
    .A2(net294));
 sg13g2_nand2_1 _19381_ (.Y(_03420_),
    .A(\top_ihp.oisc.regs[61][26] ),
    .B(_03406_));
 sg13g2_o21ai_1 _19382_ (.B1(_03420_),
    .Y(_02200_),
    .A1(net90),
    .A2(_03417_));
 sg13g2_nand2_1 _19383_ (.Y(_03421_),
    .A(\top_ihp.oisc.regs[61][27] ),
    .B(_03406_));
 sg13g2_o21ai_1 _19384_ (.B1(_03421_),
    .Y(_02201_),
    .A1(net45),
    .A2(net294));
 sg13g2_buf_1 _19385_ (.A(_03398_),
    .X(_03422_));
 sg13g2_nand2_1 _19386_ (.Y(_03423_),
    .A(\top_ihp.oisc.regs[61][28] ),
    .B(_03422_));
 sg13g2_o21ai_1 _19387_ (.B1(_03423_),
    .Y(_02202_),
    .A1(net44),
    .A2(net294));
 sg13g2_nand2_1 _19388_ (.Y(_03424_),
    .A(\top_ihp.oisc.regs[61][29] ),
    .B(net293));
 sg13g2_o21ai_1 _19389_ (.B1(_03424_),
    .Y(_02203_),
    .A1(net43),
    .A2(net294));
 sg13g2_nand2_1 _19390_ (.Y(_03425_),
    .A(\top_ihp.oisc.regs[61][2] ),
    .B(_03422_));
 sg13g2_o21ai_1 _19391_ (.B1(_03425_),
    .Y(_02204_),
    .A1(net175),
    .A2(net294));
 sg13g2_nand2_1 _19392_ (.Y(_03426_),
    .A(\top_ihp.oisc.regs[61][30] ),
    .B(net293));
 sg13g2_o21ai_1 _19393_ (.B1(_03426_),
    .Y(_02205_),
    .A1(net41),
    .A2(_03417_));
 sg13g2_nand2_1 _19394_ (.Y(_03427_),
    .A(\top_ihp.oisc.regs[61][31] ),
    .B(net293));
 sg13g2_o21ai_1 _19395_ (.B1(_03427_),
    .Y(_02206_),
    .A1(net87),
    .A2(net294));
 sg13g2_nand2_1 _19396_ (.Y(_03428_),
    .A(\top_ihp.oisc.regs[61][3] ),
    .B(net293));
 sg13g2_o21ai_1 _19397_ (.B1(_03428_),
    .Y(_02207_),
    .A1(net174),
    .A2(net294));
 sg13g2_nand2_1 _19398_ (.Y(_03429_),
    .A(\top_ihp.oisc.regs[61][4] ),
    .B(net293));
 sg13g2_o21ai_1 _19399_ (.B1(_03429_),
    .Y(_02208_),
    .A1(net88),
    .A2(net296));
 sg13g2_nand2_1 _19400_ (.Y(_03430_),
    .A(\top_ihp.oisc.regs[61][5] ),
    .B(net293));
 sg13g2_o21ai_1 _19401_ (.B1(_03430_),
    .Y(_02209_),
    .A1(_03101_),
    .A2(net296));
 sg13g2_nand2_1 _19402_ (.Y(_03431_),
    .A(\top_ihp.oisc.regs[61][6] ),
    .B(net293));
 sg13g2_o21ai_1 _19403_ (.B1(_03431_),
    .Y(_02210_),
    .A1(net177),
    .A2(net296));
 sg13g2_nand2_1 _19404_ (.Y(_03432_),
    .A(\top_ihp.oisc.regs[61][7] ),
    .B(net293));
 sg13g2_o21ai_1 _19405_ (.B1(_03432_),
    .Y(_02211_),
    .A1(_09910_),
    .A2(_03400_));
 sg13g2_nand2_1 _19406_ (.Y(_03433_),
    .A(\top_ihp.oisc.regs[61][8] ),
    .B(_03398_));
 sg13g2_o21ai_1 _19407_ (.B1(_03433_),
    .Y(_02212_),
    .A1(net42),
    .A2(_03400_));
 sg13g2_nand2_1 _19408_ (.Y(_03434_),
    .A(\top_ihp.oisc.regs[61][9] ),
    .B(_03398_));
 sg13g2_o21ai_1 _19409_ (.B1(_03434_),
    .Y(_02213_),
    .A1(_03108_),
    .A2(net296));
 sg13g2_nor2_1 _19410_ (.A(_10090_),
    .B(_03050_),
    .Y(_03435_));
 sg13g2_buf_1 _19411_ (.A(_03435_),
    .X(_03436_));
 sg13g2_mux2_1 _19412_ (.A0(\top_ihp.oisc.regs[62][0] ),
    .A1(_09199_),
    .S(net629),
    .X(_02214_));
 sg13g2_nand3_1 _19413_ (.B(net665),
    .C(_02763_),
    .A(net711),
    .Y(_03437_));
 sg13g2_buf_2 _19414_ (.A(_03437_),
    .X(_03438_));
 sg13g2_buf_1 _19415_ (.A(_03438_),
    .X(_03439_));
 sg13g2_buf_1 _19416_ (.A(_03438_),
    .X(_03440_));
 sg13g2_nand2_1 _19417_ (.Y(_03441_),
    .A(\top_ihp.oisc.regs[62][10] ),
    .B(net291));
 sg13g2_o21ai_1 _19418_ (.B1(_03441_),
    .Y(_02215_),
    .A1(net26),
    .A2(net292));
 sg13g2_nand2_1 _19419_ (.Y(_03442_),
    .A(\top_ihp.oisc.regs[62][11] ),
    .B(net291));
 sg13g2_o21ai_1 _19420_ (.B1(_03442_),
    .Y(_02216_),
    .A1(net89),
    .A2(net292));
 sg13g2_nand2_1 _19421_ (.Y(_03443_),
    .A(\top_ihp.oisc.regs[62][12] ),
    .B(net291));
 sg13g2_o21ai_1 _19422_ (.B1(_03443_),
    .Y(_02217_),
    .A1(net180),
    .A2(net292));
 sg13g2_nor2_1 _19423_ (.A(\top_ihp.oisc.regs[62][13] ),
    .B(net629),
    .Y(_03444_));
 sg13g2_a21oi_1 _19424_ (.A1(_09375_),
    .A2(net629),
    .Y(_02218_),
    .B1(_03444_));
 sg13g2_nand2_1 _19425_ (.Y(_03445_),
    .A(\top_ihp.oisc.regs[62][14] ),
    .B(net291));
 sg13g2_o21ai_1 _19426_ (.B1(_03445_),
    .Y(_02219_),
    .A1(net95),
    .A2(net292));
 sg13g2_buf_1 _19427_ (.A(_03438_),
    .X(_03446_));
 sg13g2_nand2_1 _19428_ (.Y(_03447_),
    .A(\top_ihp.oisc.regs[62][15] ),
    .B(net290));
 sg13g2_o21ai_1 _19429_ (.B1(_03447_),
    .Y(_02220_),
    .A1(net176),
    .A2(net292));
 sg13g2_nor2_1 _19430_ (.A(\top_ihp.oisc.regs[62][16] ),
    .B(net629),
    .Y(_03448_));
 sg13g2_a21oi_1 _19431_ (.A1(_09437_),
    .A2(net629),
    .Y(_02221_),
    .B1(_03448_));
 sg13g2_nand2_1 _19432_ (.Y(_03449_),
    .A(\top_ihp.oisc.regs[62][17] ),
    .B(net290));
 sg13g2_o21ai_1 _19433_ (.B1(_03449_),
    .Y(_02222_),
    .A1(net94),
    .A2(net292));
 sg13g2_nand2_1 _19434_ (.Y(_03450_),
    .A(\top_ihp.oisc.regs[62][18] ),
    .B(net290));
 sg13g2_o21ai_1 _19435_ (.B1(_03450_),
    .Y(_02223_),
    .A1(net93),
    .A2(net292));
 sg13g2_nand2_1 _19436_ (.Y(_03451_),
    .A(\top_ihp.oisc.regs[62][19] ),
    .B(net290));
 sg13g2_o21ai_1 _19437_ (.B1(_03451_),
    .Y(_02224_),
    .A1(net92),
    .A2(net292));
 sg13g2_nand2_1 _19438_ (.Y(_03452_),
    .A(\top_ihp.oisc.regs[62][1] ),
    .B(_03446_));
 sg13g2_o21ai_1 _19439_ (.B1(_03452_),
    .Y(_02225_),
    .A1(net496),
    .A2(_03439_));
 sg13g2_nor2_1 _19440_ (.A(\top_ihp.oisc.regs[62][20] ),
    .B(net629),
    .Y(_03453_));
 sg13g2_a21oi_1 _19441_ (.A1(_09581_),
    .A2(net629),
    .Y(_02226_),
    .B1(_03453_));
 sg13g2_nand2_1 _19442_ (.Y(_03454_),
    .A(\top_ihp.oisc.regs[62][21] ),
    .B(net290));
 sg13g2_o21ai_1 _19443_ (.B1(_03454_),
    .Y(_02227_),
    .A1(_03078_),
    .A2(_03439_));
 sg13g2_nor2_1 _19444_ (.A(\top_ihp.oisc.regs[62][22] ),
    .B(_03436_),
    .Y(_03455_));
 sg13g2_a21oi_1 _19445_ (.A1(_09623_),
    .A2(_03436_),
    .Y(_02228_),
    .B1(_03455_));
 sg13g2_nor2_1 _19446_ (.A(\top_ihp.oisc.regs[62][23] ),
    .B(_03435_),
    .Y(_03456_));
 sg13g2_a21oi_1 _19447_ (.A1(_09643_),
    .A2(net629),
    .Y(_02229_),
    .B1(_03456_));
 sg13g2_buf_1 _19448_ (.A(_03438_),
    .X(_03457_));
 sg13g2_nand2_1 _19449_ (.Y(_03458_),
    .A(\top_ihp.oisc.regs[62][24] ),
    .B(net290));
 sg13g2_o21ai_1 _19450_ (.B1(_03458_),
    .Y(_02230_),
    .A1(_03083_),
    .A2(net289));
 sg13g2_nand2_1 _19451_ (.Y(_03459_),
    .A(\top_ihp.oisc.regs[62][25] ),
    .B(net290));
 sg13g2_o21ai_1 _19452_ (.B1(_03459_),
    .Y(_02231_),
    .A1(_03086_),
    .A2(net289));
 sg13g2_nand2_1 _19453_ (.Y(_03460_),
    .A(\top_ihp.oisc.regs[62][26] ),
    .B(_03446_));
 sg13g2_o21ai_1 _19454_ (.B1(_03460_),
    .Y(_02232_),
    .A1(net90),
    .A2(net289));
 sg13g2_nand2_1 _19455_ (.Y(_03461_),
    .A(\top_ihp.oisc.regs[62][27] ),
    .B(net290));
 sg13g2_o21ai_1 _19456_ (.B1(_03461_),
    .Y(_02233_),
    .A1(net45),
    .A2(net289));
 sg13g2_buf_1 _19457_ (.A(_03438_),
    .X(_03462_));
 sg13g2_nand2_1 _19458_ (.Y(_03463_),
    .A(\top_ihp.oisc.regs[62][28] ),
    .B(net288));
 sg13g2_o21ai_1 _19459_ (.B1(_03463_),
    .Y(_02234_),
    .A1(net44),
    .A2(net289));
 sg13g2_nand2_1 _19460_ (.Y(_03464_),
    .A(\top_ihp.oisc.regs[62][29] ),
    .B(net288));
 sg13g2_o21ai_1 _19461_ (.B1(_03464_),
    .Y(_02235_),
    .A1(_03094_),
    .A2(net289));
 sg13g2_nand2_1 _19462_ (.Y(_03465_),
    .A(\top_ihp.oisc.regs[62][2] ),
    .B(net288));
 sg13g2_o21ai_1 _19463_ (.B1(_03465_),
    .Y(_02236_),
    .A1(net175),
    .A2(_03457_));
 sg13g2_nand2_1 _19464_ (.Y(_03466_),
    .A(\top_ihp.oisc.regs[62][30] ),
    .B(_03462_));
 sg13g2_o21ai_1 _19465_ (.B1(_03466_),
    .Y(_02237_),
    .A1(_03145_),
    .A2(net289));
 sg13g2_nand2_1 _19466_ (.Y(_03467_),
    .A(\top_ihp.oisc.regs[62][31] ),
    .B(net288));
 sg13g2_o21ai_1 _19467_ (.B1(_03467_),
    .Y(_02238_),
    .A1(_03190_),
    .A2(net289));
 sg13g2_nand2_1 _19468_ (.Y(_03468_),
    .A(\top_ihp.oisc.regs[62][3] ),
    .B(_03462_));
 sg13g2_o21ai_1 _19469_ (.B1(_03468_),
    .Y(_02239_),
    .A1(_03148_),
    .A2(_03457_));
 sg13g2_nand2_1 _19470_ (.Y(_03469_),
    .A(\top_ihp.oisc.regs[62][4] ),
    .B(net288));
 sg13g2_o21ai_1 _19471_ (.B1(_03469_),
    .Y(_02240_),
    .A1(net88),
    .A2(net291));
 sg13g2_nand2_1 _19472_ (.Y(_03470_),
    .A(\top_ihp.oisc.regs[62][5] ),
    .B(net288));
 sg13g2_o21ai_1 _19473_ (.B1(_03470_),
    .Y(_02241_),
    .A1(_03101_),
    .A2(_03440_));
 sg13g2_nand2_1 _19474_ (.Y(_03471_),
    .A(\top_ihp.oisc.regs[62][6] ),
    .B(net288));
 sg13g2_o21ai_1 _19475_ (.B1(_03471_),
    .Y(_02242_),
    .A1(net177),
    .A2(_03440_));
 sg13g2_nand2_1 _19476_ (.Y(_03472_),
    .A(\top_ihp.oisc.regs[62][7] ),
    .B(net288));
 sg13g2_o21ai_1 _19477_ (.B1(_03472_),
    .Y(_02243_),
    .A1(_02718_),
    .A2(net291));
 sg13g2_nand2_1 _19478_ (.Y(_03473_),
    .A(\top_ihp.oisc.regs[62][8] ),
    .B(_03438_));
 sg13g2_o21ai_1 _19479_ (.B1(_03473_),
    .Y(_02244_),
    .A1(_03106_),
    .A2(net291));
 sg13g2_nand2_1 _19480_ (.Y(_03474_),
    .A(\top_ihp.oisc.regs[62][9] ),
    .B(_03438_));
 sg13g2_o21ai_1 _19481_ (.B1(_03474_),
    .Y(_02245_),
    .A1(net25),
    .A2(net291));
 sg13g2_nor2_2 _19482_ (.A(_10090_),
    .B(_03110_),
    .Y(_03475_));
 sg13g2_mux2_1 _19483_ (.A0(\top_ihp.oisc.regs[63][0] ),
    .A1(_09199_),
    .S(_03475_),
    .X(_02246_));
 sg13g2_nand3_1 _19484_ (.B(_10055_),
    .C(_02763_),
    .A(_10009_),
    .Y(_03476_));
 sg13g2_buf_1 _19485_ (.A(_03476_),
    .X(_03477_));
 sg13g2_buf_2 _19486_ (.A(_03477_),
    .X(_03478_));
 sg13g2_buf_1 _19487_ (.A(net483),
    .X(_03479_));
 sg13g2_buf_1 _19488_ (.A(_03477_),
    .X(_03480_));
 sg13g2_nand2_1 _19489_ (.Y(_03481_),
    .A(\top_ihp.oisc.regs[63][10] ),
    .B(net482));
 sg13g2_o21ai_1 _19490_ (.B1(_03481_),
    .Y(_02247_),
    .A1(_10063_),
    .A2(net287));
 sg13g2_buf_1 _19491_ (.A(_03477_),
    .X(_03482_));
 sg13g2_nand2_1 _19492_ (.Y(_03483_),
    .A(\top_ihp.oisc.regs[63][11] ),
    .B(net481));
 sg13g2_o21ai_1 _19493_ (.B1(_03483_),
    .Y(_02248_),
    .A1(net89),
    .A2(net287));
 sg13g2_nand2_1 _19494_ (.Y(_03484_),
    .A(\top_ihp.oisc.regs[63][12] ),
    .B(net481));
 sg13g2_o21ai_1 _19495_ (.B1(_03484_),
    .Y(_02249_),
    .A1(net218),
    .A2(net287));
 sg13g2_nand2_1 _19496_ (.Y(_03485_),
    .A(\top_ihp.oisc.regs[63][13] ),
    .B(net481));
 sg13g2_o21ai_1 _19497_ (.B1(_03485_),
    .Y(_02250_),
    .A1(_09374_),
    .A2(_03479_));
 sg13g2_nand2_1 _19498_ (.Y(_03486_),
    .A(\top_ihp.oisc.regs[63][14] ),
    .B(net481));
 sg13g2_o21ai_1 _19499_ (.B1(_03486_),
    .Y(_02251_),
    .A1(_10066_),
    .A2(net287));
 sg13g2_nand2_1 _19500_ (.Y(_03487_),
    .A(\top_ihp.oisc.regs[63][15] ),
    .B(net481));
 sg13g2_o21ai_1 _19501_ (.B1(_03487_),
    .Y(_02252_),
    .A1(net176),
    .A2(net287));
 sg13g2_nand2_1 _19502_ (.Y(_03488_),
    .A(\top_ihp.oisc.regs[63][16] ),
    .B(_03482_));
 sg13g2_o21ai_1 _19503_ (.B1(_03488_),
    .Y(_02253_),
    .A1(net247),
    .A2(_03479_));
 sg13g2_nand2_1 _19504_ (.Y(_03489_),
    .A(\top_ihp.oisc.regs[63][17] ),
    .B(net481));
 sg13g2_o21ai_1 _19505_ (.B1(_03489_),
    .Y(_02254_),
    .A1(_10070_),
    .A2(net287));
 sg13g2_nand2_1 _19506_ (.Y(_03490_),
    .A(\top_ihp.oisc.regs[63][18] ),
    .B(_03482_));
 sg13g2_o21ai_1 _19507_ (.B1(_03490_),
    .Y(_02255_),
    .A1(net135),
    .A2(net287));
 sg13g2_nand2_1 _19508_ (.Y(_03491_),
    .A(\top_ihp.oisc.regs[63][19] ),
    .B(net481));
 sg13g2_o21ai_1 _19509_ (.B1(_03491_),
    .Y(_02256_),
    .A1(_10072_),
    .A2(net287));
 sg13g2_buf_2 _19510_ (.A(net483),
    .X(_03492_));
 sg13g2_nand2_1 _19511_ (.Y(_03493_),
    .A(\top_ihp.oisc.regs[63][1] ),
    .B(net481));
 sg13g2_o21ai_1 _19512_ (.B1(_03493_),
    .Y(_02257_),
    .A1(_09553_),
    .A2(net286));
 sg13g2_mux2_1 _19513_ (.A0(\top_ihp.oisc.regs[63][20] ),
    .A1(_09573_),
    .S(_03475_),
    .X(_02258_));
 sg13g2_buf_1 _19514_ (.A(_03477_),
    .X(_03494_));
 sg13g2_nand2_1 _19515_ (.Y(_03495_),
    .A(\top_ihp.oisc.regs[63][21] ),
    .B(net480));
 sg13g2_o21ai_1 _19516_ (.B1(_03495_),
    .Y(_02259_),
    .A1(net64),
    .A2(net286));
 sg13g2_nand2_1 _19517_ (.Y(_03496_),
    .A(\top_ihp.oisc.regs[63][22] ),
    .B(net480));
 sg13g2_o21ai_1 _19518_ (.B1(_03496_),
    .Y(_02260_),
    .A1(_09622_),
    .A2(net286));
 sg13g2_mux2_1 _19519_ (.A0(\top_ihp.oisc.regs[63][23] ),
    .A1(net406),
    .S(_03475_),
    .X(_02261_));
 sg13g2_nand2_1 _19520_ (.Y(_03497_),
    .A(\top_ihp.oisc.regs[63][24] ),
    .B(net480));
 sg13g2_o21ai_1 _19521_ (.B1(_03497_),
    .Y(_02262_),
    .A1(_10077_),
    .A2(net286));
 sg13g2_nand2_1 _19522_ (.Y(_03498_),
    .A(\top_ihp.oisc.regs[63][25] ),
    .B(net480));
 sg13g2_o21ai_1 _19523_ (.B1(_03498_),
    .Y(_02263_),
    .A1(_10078_),
    .A2(net286));
 sg13g2_nand2_1 _19524_ (.Y(_03499_),
    .A(\top_ihp.oisc.regs[63][26] ),
    .B(net480));
 sg13g2_o21ai_1 _19525_ (.B1(_03499_),
    .Y(_02264_),
    .A1(net134),
    .A2(net286));
 sg13g2_nand2_1 _19526_ (.Y(_03500_),
    .A(\top_ihp.oisc.regs[63][27] ),
    .B(net480));
 sg13g2_o21ai_1 _19527_ (.B1(_03500_),
    .Y(_02265_),
    .A1(_09702_),
    .A2(net286));
 sg13g2_nand2_1 _19528_ (.Y(_03501_),
    .A(\top_ihp.oisc.regs[63][28] ),
    .B(_03494_));
 sg13g2_o21ai_1 _19529_ (.B1(_03501_),
    .Y(_02266_),
    .A1(_10081_),
    .A2(_03492_));
 sg13g2_nand2_1 _19530_ (.Y(_03502_),
    .A(\top_ihp.oisc.regs[63][29] ),
    .B(net480));
 sg13g2_o21ai_1 _19531_ (.B1(_03502_),
    .Y(_02267_),
    .A1(_10083_),
    .A2(net286));
 sg13g2_nand2_1 _19532_ (.Y(_03503_),
    .A(\top_ihp.oisc.regs[63][2] ),
    .B(_03494_));
 sg13g2_o21ai_1 _19533_ (.B1(_03503_),
    .Y(_02268_),
    .A1(net175),
    .A2(_03492_));
 sg13g2_nand2_1 _19534_ (.Y(_03504_),
    .A(\top_ihp.oisc.regs[63][30] ),
    .B(net480));
 sg13g2_o21ai_1 _19535_ (.B1(_03504_),
    .Y(_02269_),
    .A1(net41),
    .A2(net482));
 sg13g2_nand2_1 _19536_ (.Y(_03505_),
    .A(\top_ihp.oisc.regs[63][31] ),
    .B(net483));
 sg13g2_o21ai_1 _19537_ (.B1(_03505_),
    .Y(_02270_),
    .A1(_03190_),
    .A2(_03480_));
 sg13g2_nand2_1 _19538_ (.Y(_03506_),
    .A(\top_ihp.oisc.regs[63][3] ),
    .B(net483));
 sg13g2_o21ai_1 _19539_ (.B1(_03506_),
    .Y(_02271_),
    .A1(net174),
    .A2(net482));
 sg13g2_nand2_1 _19540_ (.Y(_03507_),
    .A(\top_ihp.oisc.regs[63][4] ),
    .B(_03478_));
 sg13g2_o21ai_1 _19541_ (.B1(_03507_),
    .Y(_02272_),
    .A1(net88),
    .A2(net482));
 sg13g2_nand2_1 _19542_ (.Y(_03508_),
    .A(\top_ihp.oisc.regs[63][5] ),
    .B(net483));
 sg13g2_o21ai_1 _19543_ (.B1(_03508_),
    .Y(_02273_),
    .A1(_10085_),
    .A2(net482));
 sg13g2_nand2_1 _19544_ (.Y(_03509_),
    .A(\top_ihp.oisc.regs[63][6] ),
    .B(net483));
 sg13g2_o21ai_1 _19545_ (.B1(_03509_),
    .Y(_02274_),
    .A1(_10086_),
    .A2(net482));
 sg13g2_nand2_1 _19546_ (.Y(_03510_),
    .A(\top_ihp.oisc.regs[63][7] ),
    .B(_03478_));
 sg13g2_o21ai_1 _19547_ (.B1(_03510_),
    .Y(_02275_),
    .A1(_09910_),
    .A2(_03480_));
 sg13g2_nand2_1 _19548_ (.Y(_03511_),
    .A(\top_ihp.oisc.regs[63][8] ),
    .B(net483));
 sg13g2_o21ai_1 _19549_ (.B1(_03511_),
    .Y(_02276_),
    .A1(_10087_),
    .A2(net482));
 sg13g2_nand2_1 _19550_ (.Y(_03512_),
    .A(\top_ihp.oisc.regs[63][9] ),
    .B(net483));
 sg13g2_o21ai_1 _19551_ (.B1(_03512_),
    .Y(_02277_),
    .A1(_10088_),
    .A2(net482));
 sg13g2_nor2_2 _19552_ (.A(_09962_),
    .B(net682),
    .Y(_03513_));
 sg13g2_mux2_1 _19553_ (.A0(\top_ihp.oisc.regs[6][0] ),
    .A1(net412),
    .S(_03513_),
    .X(_02278_));
 sg13g2_nand2b_1 _19554_ (.Y(_03514_),
    .B(_10397_),
    .A_N(_09962_));
 sg13g2_buf_1 _19555_ (.A(_03514_),
    .X(_03515_));
 sg13g2_buf_1 _19556_ (.A(_03515_),
    .X(_03516_));
 sg13g2_buf_1 _19557_ (.A(net285),
    .X(_03517_));
 sg13g2_buf_1 _19558_ (.A(_03515_),
    .X(_03518_));
 sg13g2_nand2_1 _19559_ (.Y(_03519_),
    .A(\top_ihp.oisc.regs[6][10] ),
    .B(net284));
 sg13g2_o21ai_1 _19560_ (.B1(_03519_),
    .Y(_02279_),
    .A1(net65),
    .A2(net160));
 sg13g2_buf_1 _19561_ (.A(_03515_),
    .X(_03520_));
 sg13g2_nand2_1 _19562_ (.Y(_03521_),
    .A(\top_ihp.oisc.regs[6][11] ),
    .B(net283));
 sg13g2_o21ai_1 _19563_ (.B1(_03521_),
    .Y(_02280_),
    .A1(net251),
    .A2(net160));
 sg13g2_nand2_1 _19564_ (.Y(_03522_),
    .A(\top_ihp.oisc.regs[6][12] ),
    .B(net283));
 sg13g2_o21ai_1 _19565_ (.B1(_03522_),
    .Y(_02281_),
    .A1(net218),
    .A2(net160));
 sg13g2_nand2_1 _19566_ (.Y(_03523_),
    .A(\top_ihp.oisc.regs[6][13] ),
    .B(_03520_));
 sg13g2_o21ai_1 _19567_ (.B1(_03523_),
    .Y(_02282_),
    .A1(net147),
    .A2(_03517_));
 sg13g2_nand2_1 _19568_ (.Y(_03524_),
    .A(\top_ihp.oisc.regs[6][14] ),
    .B(net283));
 sg13g2_o21ai_1 _19569_ (.B1(_03524_),
    .Y(_02283_),
    .A1(net217),
    .A2(net160));
 sg13g2_nand2_1 _19570_ (.Y(_03525_),
    .A(\top_ihp.oisc.regs[6][15] ),
    .B(net283));
 sg13g2_o21ai_1 _19571_ (.B1(_03525_),
    .Y(_02284_),
    .A1(net216),
    .A2(net160));
 sg13g2_nand2_1 _19572_ (.Y(_03526_),
    .A(\top_ihp.oisc.regs[6][16] ),
    .B(_03520_));
 sg13g2_o21ai_1 _19573_ (.B1(_03526_),
    .Y(_02285_),
    .A1(net247),
    .A2(net160));
 sg13g2_nand2_1 _19574_ (.Y(_03527_),
    .A(\top_ihp.oisc.regs[6][17] ),
    .B(net283));
 sg13g2_o21ai_1 _19575_ (.B1(_03527_),
    .Y(_02286_),
    .A1(net136),
    .A2(net160));
 sg13g2_nand2_1 _19576_ (.Y(_03528_),
    .A(\top_ihp.oisc.regs[6][18] ),
    .B(net283));
 sg13g2_o21ai_1 _19577_ (.B1(_03528_),
    .Y(_02287_),
    .A1(net135),
    .A2(net160));
 sg13g2_nand2_1 _19578_ (.Y(_03529_),
    .A(\top_ihp.oisc.regs[6][19] ),
    .B(net283));
 sg13g2_o21ai_1 _19579_ (.B1(_03529_),
    .Y(_02288_),
    .A1(net215),
    .A2(_03517_));
 sg13g2_buf_1 _19580_ (.A(net285),
    .X(_03530_));
 sg13g2_nand2_1 _19581_ (.Y(_03531_),
    .A(\top_ihp.oisc.regs[6][1] ),
    .B(net283));
 sg13g2_o21ai_1 _19582_ (.B1(_03531_),
    .Y(_02289_),
    .A1(net547),
    .A2(net159));
 sg13g2_nor2_1 _19583_ (.A(\top_ihp.oisc.regs[6][20] ),
    .B(_03513_),
    .Y(_03532_));
 sg13g2_a21oi_1 _19584_ (.A1(_09581_),
    .A2(_03513_),
    .Y(_02290_),
    .B1(_03532_));
 sg13g2_buf_1 _19585_ (.A(_03515_),
    .X(_03533_));
 sg13g2_nand2_1 _19586_ (.Y(_03534_),
    .A(\top_ihp.oisc.regs[6][21] ),
    .B(_03533_));
 sg13g2_o21ai_1 _19587_ (.B1(_03534_),
    .Y(_02291_),
    .A1(net64),
    .A2(net159));
 sg13g2_nand2_1 _19588_ (.Y(_03535_),
    .A(\top_ihp.oisc.regs[6][22] ),
    .B(net282));
 sg13g2_o21ai_1 _19589_ (.B1(_03535_),
    .Y(_02292_),
    .A1(net244),
    .A2(net159));
 sg13g2_nor2_1 _19590_ (.A(\top_ihp.oisc.regs[6][23] ),
    .B(_03513_),
    .Y(_03536_));
 sg13g2_a21oi_1 _19591_ (.A1(net243),
    .A2(_03513_),
    .Y(_02293_),
    .B1(_03536_));
 sg13g2_nand2_1 _19592_ (.Y(_03537_),
    .A(\top_ihp.oisc.regs[6][24] ),
    .B(net282));
 sg13g2_o21ai_1 _19593_ (.B1(_03537_),
    .Y(_02294_),
    .A1(net214),
    .A2(net159));
 sg13g2_nand2_1 _19594_ (.Y(_03538_),
    .A(\top_ihp.oisc.regs[6][25] ),
    .B(net282));
 sg13g2_o21ai_1 _19595_ (.B1(_03538_),
    .Y(_02295_),
    .A1(_10078_),
    .A2(net159));
 sg13g2_nand2_1 _19596_ (.Y(_03539_),
    .A(\top_ihp.oisc.regs[6][26] ),
    .B(net282));
 sg13g2_o21ai_1 _19597_ (.B1(_03539_),
    .Y(_02296_),
    .A1(_10079_),
    .A2(net159));
 sg13g2_nand2_1 _19598_ (.Y(_03540_),
    .A(\top_ihp.oisc.regs[6][27] ),
    .B(net282));
 sg13g2_o21ai_1 _19599_ (.B1(_03540_),
    .Y(_02297_),
    .A1(net141),
    .A2(net159));
 sg13g2_nand2_1 _19600_ (.Y(_03541_),
    .A(\top_ihp.oisc.regs[6][28] ),
    .B(_03533_));
 sg13g2_o21ai_1 _19601_ (.B1(_03541_),
    .Y(_02298_),
    .A1(net63),
    .A2(_03530_));
 sg13g2_nand2_1 _19602_ (.Y(_03542_),
    .A(\top_ihp.oisc.regs[6][29] ),
    .B(net282));
 sg13g2_o21ai_1 _19603_ (.B1(_03542_),
    .Y(_02299_),
    .A1(net133),
    .A2(net159));
 sg13g2_nand2_1 _19604_ (.Y(_03543_),
    .A(\top_ihp.oisc.regs[6][2] ),
    .B(net282));
 sg13g2_o21ai_1 _19605_ (.B1(_03543_),
    .Y(_02300_),
    .A1(_10044_),
    .A2(_03530_));
 sg13g2_nand2_1 _19606_ (.Y(_03544_),
    .A(\top_ihp.oisc.regs[6][30] ),
    .B(net282));
 sg13g2_o21ai_1 _19607_ (.B1(_03544_),
    .Y(_02301_),
    .A1(_10084_),
    .A2(_03518_));
 sg13g2_nand2_1 _19608_ (.Y(_03545_),
    .A(\top_ihp.oisc.regs[6][31] ),
    .B(_03516_));
 sg13g2_o21ai_1 _19609_ (.B1(_03545_),
    .Y(_02302_),
    .A1(net87),
    .A2(net284));
 sg13g2_nand2_1 _19610_ (.Y(_03546_),
    .A(\top_ihp.oisc.regs[6][3] ),
    .B(_03516_));
 sg13g2_o21ai_1 _19611_ (.B1(_03546_),
    .Y(_02303_),
    .A1(_10047_),
    .A2(net284));
 sg13g2_nand2_1 _19612_ (.Y(_03547_),
    .A(\top_ihp.oisc.regs[6][4] ),
    .B(net285));
 sg13g2_o21ai_1 _19613_ (.B1(_03547_),
    .Y(_02304_),
    .A1(_10048_),
    .A2(_03518_));
 sg13g2_nand2_1 _19614_ (.Y(_03548_),
    .A(\top_ihp.oisc.regs[6][5] ),
    .B(net285));
 sg13g2_o21ai_1 _19615_ (.B1(_03548_),
    .Y(_02305_),
    .A1(net212),
    .A2(net284));
 sg13g2_nand2_1 _19616_ (.Y(_03549_),
    .A(\top_ihp.oisc.regs[6][6] ),
    .B(net285));
 sg13g2_o21ai_1 _19617_ (.B1(_03549_),
    .Y(_02306_),
    .A1(_10086_),
    .A2(net284));
 sg13g2_nand2_1 _19618_ (.Y(_03550_),
    .A(\top_ihp.oisc.regs[6][7] ),
    .B(net285));
 sg13g2_o21ai_1 _19619_ (.B1(_03550_),
    .Y(_02307_),
    .A1(net47),
    .A2(net284));
 sg13g2_nand2_1 _19620_ (.Y(_03551_),
    .A(\top_ihp.oisc.regs[6][8] ),
    .B(net285));
 sg13g2_o21ai_1 _19621_ (.B1(_03551_),
    .Y(_02308_),
    .A1(_10087_),
    .A2(net284));
 sg13g2_nand2_1 _19622_ (.Y(_03552_),
    .A(\top_ihp.oisc.regs[6][9] ),
    .B(net285));
 sg13g2_o21ai_1 _19623_ (.B1(_03552_),
    .Y(_02309_),
    .A1(_10088_),
    .A2(net284));
 sg13g2_and2_1 _19624_ (.A(_10011_),
    .B(net663),
    .X(_03553_));
 sg13g2_buf_1 _19625_ (.A(_03553_),
    .X(_03554_));
 sg13g2_mux2_1 _19626_ (.A0(\top_ihp.oisc.regs[7][0] ),
    .A1(net412),
    .S(_03554_),
    .X(_02310_));
 sg13g2_nand2_1 _19627_ (.Y(_03555_),
    .A(_10011_),
    .B(net663));
 sg13g2_buf_1 _19628_ (.A(_03555_),
    .X(_03556_));
 sg13g2_buf_1 _19629_ (.A(net478),
    .X(_03557_));
 sg13g2_buf_1 _19630_ (.A(net478),
    .X(_03558_));
 sg13g2_nand2_1 _19631_ (.Y(_03559_),
    .A(\top_ihp.oisc.regs[7][10] ),
    .B(net280));
 sg13g2_o21ai_1 _19632_ (.B1(_03559_),
    .Y(_02311_),
    .A1(net65),
    .A2(net281));
 sg13g2_nand2_1 _19633_ (.Y(_03560_),
    .A(\top_ihp.oisc.regs[7][11] ),
    .B(net280));
 sg13g2_o21ai_1 _19634_ (.B1(_03560_),
    .Y(_02312_),
    .A1(net251),
    .A2(net281));
 sg13g2_nand2_1 _19635_ (.Y(_03561_),
    .A(\top_ihp.oisc.regs[7][12] ),
    .B(net280));
 sg13g2_o21ai_1 _19636_ (.B1(_03561_),
    .Y(_02313_),
    .A1(net218),
    .A2(net281));
 sg13g2_nor2_1 _19637_ (.A(\top_ihp.oisc.regs[7][13] ),
    .B(net479),
    .Y(_03562_));
 sg13g2_a21oi_1 _19638_ (.A1(net73),
    .A2(net479),
    .Y(_02314_),
    .B1(_03562_));
 sg13g2_buf_1 _19639_ (.A(net478),
    .X(_03563_));
 sg13g2_nand2_1 _19640_ (.Y(_03564_),
    .A(\top_ihp.oisc.regs[7][14] ),
    .B(net279));
 sg13g2_o21ai_1 _19641_ (.B1(_03564_),
    .Y(_02315_),
    .A1(net217),
    .A2(net281));
 sg13g2_nand2_1 _19642_ (.Y(_03565_),
    .A(\top_ihp.oisc.regs[7][15] ),
    .B(net279));
 sg13g2_o21ai_1 _19643_ (.B1(_03565_),
    .Y(_02316_),
    .A1(net216),
    .A2(net281));
 sg13g2_nor2_1 _19644_ (.A(\top_ihp.oisc.regs[7][16] ),
    .B(net479),
    .Y(_03566_));
 sg13g2_a21oi_1 _19645_ (.A1(net146),
    .A2(net479),
    .Y(_02317_),
    .B1(_03566_));
 sg13g2_nand2_1 _19646_ (.Y(_03567_),
    .A(\top_ihp.oisc.regs[7][17] ),
    .B(net279));
 sg13g2_o21ai_1 _19647_ (.B1(_03567_),
    .Y(_02318_),
    .A1(net136),
    .A2(net281));
 sg13g2_nand2_1 _19648_ (.Y(_03568_),
    .A(\top_ihp.oisc.regs[7][18] ),
    .B(net279));
 sg13g2_o21ai_1 _19649_ (.B1(_03568_),
    .Y(_02319_),
    .A1(net135),
    .A2(net281));
 sg13g2_nand2_1 _19650_ (.Y(_03569_),
    .A(\top_ihp.oisc.regs[7][19] ),
    .B(_03563_));
 sg13g2_o21ai_1 _19651_ (.B1(_03569_),
    .Y(_02320_),
    .A1(net215),
    .A2(_03557_));
 sg13g2_nand2_1 _19652_ (.Y(_03570_),
    .A(\top_ihp.oisc.regs[7][1] ),
    .B(net279));
 sg13g2_o21ai_1 _19653_ (.B1(_03570_),
    .Y(_02321_),
    .A1(net547),
    .A2(net281));
 sg13g2_nand2_1 _19654_ (.Y(_03571_),
    .A(\top_ihp.oisc.regs[7][20] ),
    .B(net279));
 sg13g2_o21ai_1 _19655_ (.B1(_03571_),
    .Y(_02322_),
    .A1(_09563_),
    .A2(_03557_));
 sg13g2_buf_1 _19656_ (.A(net478),
    .X(_03572_));
 sg13g2_nand2_1 _19657_ (.Y(_03573_),
    .A(\top_ihp.oisc.regs[7][21] ),
    .B(_03563_));
 sg13g2_o21ai_1 _19658_ (.B1(_03573_),
    .Y(_02323_),
    .A1(net64),
    .A2(_03572_));
 sg13g2_nor2_1 _19659_ (.A(\top_ihp.oisc.regs[7][22] ),
    .B(net479),
    .Y(_03574_));
 sg13g2_a21oi_1 _19660_ (.A1(net143),
    .A2(net479),
    .Y(_02324_),
    .B1(_03574_));
 sg13g2_nor2_1 _19661_ (.A(\top_ihp.oisc.regs[7][23] ),
    .B(net479),
    .Y(_03575_));
 sg13g2_a21oi_1 _19662_ (.A1(net243),
    .A2(net479),
    .Y(_02325_),
    .B1(_03575_));
 sg13g2_nand2_1 _19663_ (.Y(_03576_),
    .A(\top_ihp.oisc.regs[7][24] ),
    .B(net279));
 sg13g2_o21ai_1 _19664_ (.B1(_03576_),
    .Y(_02326_),
    .A1(net214),
    .A2(net278));
 sg13g2_nand2_1 _19665_ (.Y(_03577_),
    .A(\top_ihp.oisc.regs[7][25] ),
    .B(net279));
 sg13g2_o21ai_1 _19666_ (.B1(_03577_),
    .Y(_02327_),
    .A1(net213),
    .A2(net278));
 sg13g2_buf_1 _19667_ (.A(_03556_),
    .X(_03578_));
 sg13g2_nand2_1 _19668_ (.Y(_03579_),
    .A(\top_ihp.oisc.regs[7][26] ),
    .B(net277));
 sg13g2_o21ai_1 _19669_ (.B1(_03579_),
    .Y(_02328_),
    .A1(_10079_),
    .A2(net278));
 sg13g2_nand2_1 _19670_ (.Y(_03580_),
    .A(\top_ihp.oisc.regs[7][27] ),
    .B(net277));
 sg13g2_o21ai_1 _19671_ (.B1(_03580_),
    .Y(_02329_),
    .A1(net141),
    .A2(net278));
 sg13g2_nand2_1 _19672_ (.Y(_03581_),
    .A(\top_ihp.oisc.regs[7][28] ),
    .B(net277));
 sg13g2_o21ai_1 _19673_ (.B1(_03581_),
    .Y(_02330_),
    .A1(net63),
    .A2(net278));
 sg13g2_nand2_1 _19674_ (.Y(_03582_),
    .A(\top_ihp.oisc.regs[7][29] ),
    .B(net277));
 sg13g2_o21ai_1 _19675_ (.B1(_03582_),
    .Y(_02331_),
    .A1(net133),
    .A2(net278));
 sg13g2_nand2_1 _19676_ (.Y(_03583_),
    .A(\top_ihp.oisc.regs[7][2] ),
    .B(net277));
 sg13g2_o21ai_1 _19677_ (.B1(_03583_),
    .Y(_02332_),
    .A1(net222),
    .A2(net278));
 sg13g2_nand2_1 _19678_ (.Y(_03584_),
    .A(\top_ihp.oisc.regs[7][30] ),
    .B(_03578_));
 sg13g2_o21ai_1 _19679_ (.B1(_03584_),
    .Y(_02333_),
    .A1(_10084_),
    .A2(net278));
 sg13g2_nand2_1 _19680_ (.Y(_03585_),
    .A(\top_ihp.oisc.regs[7][31] ),
    .B(_03578_));
 sg13g2_o21ai_1 _19681_ (.B1(_03585_),
    .Y(_02334_),
    .A1(net239),
    .A2(_03572_));
 sg13g2_nand2_1 _19682_ (.Y(_03586_),
    .A(\top_ihp.oisc.regs[7][3] ),
    .B(net277));
 sg13g2_o21ai_1 _19683_ (.B1(_03586_),
    .Y(_02335_),
    .A1(net221),
    .A2(_03558_));
 sg13g2_nand2_1 _19684_ (.Y(_03587_),
    .A(\top_ihp.oisc.regs[7][4] ),
    .B(net277));
 sg13g2_o21ai_1 _19685_ (.B1(_03587_),
    .Y(_02336_),
    .A1(net220),
    .A2(_03558_));
 sg13g2_nand2_1 _19686_ (.Y(_03588_),
    .A(\top_ihp.oisc.regs[7][5] ),
    .B(net277));
 sg13g2_o21ai_1 _19687_ (.B1(_03588_),
    .Y(_02337_),
    .A1(net212),
    .A2(net280));
 sg13g2_nand2_1 _19688_ (.Y(_03589_),
    .A(\top_ihp.oisc.regs[7][6] ),
    .B(net478));
 sg13g2_o21ai_1 _19689_ (.B1(_03589_),
    .Y(_02338_),
    .A1(net211),
    .A2(net280));
 sg13g2_nand2_1 _19690_ (.Y(_03590_),
    .A(\top_ihp.oisc.regs[7][7] ),
    .B(net478));
 sg13g2_o21ai_1 _19691_ (.B1(_03590_),
    .Y(_02339_),
    .A1(net408),
    .A2(net280));
 sg13g2_nand2_1 _19692_ (.Y(_03591_),
    .A(\top_ihp.oisc.regs[7][8] ),
    .B(net478));
 sg13g2_o21ai_1 _19693_ (.B1(_03591_),
    .Y(_02340_),
    .A1(net61),
    .A2(net280));
 sg13g2_nand2_1 _19694_ (.Y(_03592_),
    .A(\top_ihp.oisc.regs[7][9] ),
    .B(net478));
 sg13g2_o21ai_1 _19695_ (.B1(_03592_),
    .Y(_02341_),
    .A1(net60),
    .A2(net280));
 sg13g2_and2_1 _19696_ (.A(net545),
    .B(_10057_),
    .X(_03593_));
 sg13g2_buf_2 _19697_ (.A(_03593_),
    .X(_03594_));
 sg13g2_mux2_1 _19698_ (.A0(\top_ihp.oisc.regs[8][0] ),
    .A1(net412),
    .S(_03594_),
    .X(_02342_));
 sg13g2_nand2_1 _19699_ (.Y(_03595_),
    .A(_10007_),
    .B(_10057_));
 sg13g2_buf_1 _19700_ (.A(_03595_),
    .X(_03596_));
 sg13g2_buf_1 _19701_ (.A(_03596_),
    .X(_03597_));
 sg13g2_buf_1 _19702_ (.A(net158),
    .X(_03598_));
 sg13g2_buf_1 _19703_ (.A(_03596_),
    .X(_03599_));
 sg13g2_nand2_1 _19704_ (.Y(_03600_),
    .A(\top_ihp.oisc.regs[8][10] ),
    .B(net157));
 sg13g2_o21ai_1 _19705_ (.B1(_03600_),
    .Y(_02343_),
    .A1(net65),
    .A2(net84));
 sg13g2_buf_1 _19706_ (.A(_03596_),
    .X(_03601_));
 sg13g2_nand2_1 _19707_ (.Y(_03602_),
    .A(\top_ihp.oisc.regs[8][11] ),
    .B(net156));
 sg13g2_o21ai_1 _19708_ (.B1(_03602_),
    .Y(_02344_),
    .A1(_09303_),
    .A2(net84));
 sg13g2_nand2_1 _19709_ (.Y(_03603_),
    .A(\top_ihp.oisc.regs[8][12] ),
    .B(net156));
 sg13g2_o21ai_1 _19710_ (.B1(_03603_),
    .Y(_02345_),
    .A1(net218),
    .A2(net84));
 sg13g2_nand2_1 _19711_ (.Y(_03604_),
    .A(\top_ihp.oisc.regs[8][13] ),
    .B(_03601_));
 sg13g2_o21ai_1 _19712_ (.B1(_03604_),
    .Y(_02346_),
    .A1(_09374_),
    .A2(net84));
 sg13g2_nand2_1 _19713_ (.Y(_03605_),
    .A(\top_ihp.oisc.regs[8][14] ),
    .B(net156));
 sg13g2_o21ai_1 _19714_ (.B1(_03605_),
    .Y(_02347_),
    .A1(net217),
    .A2(net84));
 sg13g2_nand2_1 _19715_ (.Y(_03606_),
    .A(\top_ihp.oisc.regs[8][15] ),
    .B(net156));
 sg13g2_o21ai_1 _19716_ (.B1(_03606_),
    .Y(_02348_),
    .A1(net216),
    .A2(net84));
 sg13g2_nand2_1 _19717_ (.Y(_03607_),
    .A(\top_ihp.oisc.regs[8][16] ),
    .B(net156));
 sg13g2_o21ai_1 _19718_ (.B1(_03607_),
    .Y(_02349_),
    .A1(net247),
    .A2(_03598_));
 sg13g2_nand2_1 _19719_ (.Y(_03608_),
    .A(\top_ihp.oisc.regs[8][17] ),
    .B(net156));
 sg13g2_o21ai_1 _19720_ (.B1(_03608_),
    .Y(_02350_),
    .A1(net136),
    .A2(net84));
 sg13g2_nand2_1 _19721_ (.Y(_03609_),
    .A(\top_ihp.oisc.regs[8][18] ),
    .B(net156));
 sg13g2_o21ai_1 _19722_ (.B1(_03609_),
    .Y(_02351_),
    .A1(net135),
    .A2(_03598_));
 sg13g2_nand2_1 _19723_ (.Y(_03610_),
    .A(\top_ihp.oisc.regs[8][19] ),
    .B(net156));
 sg13g2_o21ai_1 _19724_ (.B1(_03610_),
    .Y(_02352_),
    .A1(net215),
    .A2(net84));
 sg13g2_buf_1 _19725_ (.A(net158),
    .X(_03611_));
 sg13g2_nand2_1 _19726_ (.Y(_03612_),
    .A(\top_ihp.oisc.regs[8][1] ),
    .B(_03601_));
 sg13g2_o21ai_1 _19727_ (.B1(_03612_),
    .Y(_02353_),
    .A1(net547),
    .A2(net83));
 sg13g2_nor2_1 _19728_ (.A(\top_ihp.oisc.regs[8][20] ),
    .B(_03594_),
    .Y(_03613_));
 sg13g2_a21oi_1 _19729_ (.A1(_09581_),
    .A2(_03594_),
    .Y(_02354_),
    .B1(_03613_));
 sg13g2_buf_1 _19730_ (.A(_03596_),
    .X(_03614_));
 sg13g2_nand2_1 _19731_ (.Y(_03615_),
    .A(\top_ihp.oisc.regs[8][21] ),
    .B(net155));
 sg13g2_o21ai_1 _19732_ (.B1(_03615_),
    .Y(_02355_),
    .A1(net64),
    .A2(net83));
 sg13g2_nand2_1 _19733_ (.Y(_03616_),
    .A(\top_ihp.oisc.regs[8][22] ),
    .B(net155));
 sg13g2_o21ai_1 _19734_ (.B1(_03616_),
    .Y(_02356_),
    .A1(net244),
    .A2(net83));
 sg13g2_nor2_1 _19735_ (.A(\top_ihp.oisc.regs[8][23] ),
    .B(_03594_),
    .Y(_03617_));
 sg13g2_a21oi_1 _19736_ (.A1(net243),
    .A2(_03594_),
    .Y(_02357_),
    .B1(_03617_));
 sg13g2_nand2_1 _19737_ (.Y(_03618_),
    .A(\top_ihp.oisc.regs[8][24] ),
    .B(_03614_));
 sg13g2_o21ai_1 _19738_ (.B1(_03618_),
    .Y(_02358_),
    .A1(net214),
    .A2(_03611_));
 sg13g2_nand2_1 _19739_ (.Y(_03619_),
    .A(\top_ihp.oisc.regs[8][25] ),
    .B(net155));
 sg13g2_o21ai_1 _19740_ (.B1(_03619_),
    .Y(_02359_),
    .A1(net213),
    .A2(net83));
 sg13g2_nand2_1 _19741_ (.Y(_03620_),
    .A(\top_ihp.oisc.regs[8][26] ),
    .B(net155));
 sg13g2_o21ai_1 _19742_ (.B1(_03620_),
    .Y(_02360_),
    .A1(net134),
    .A2(net83));
 sg13g2_nand2_1 _19743_ (.Y(_03621_),
    .A(\top_ihp.oisc.regs[8][27] ),
    .B(net155));
 sg13g2_o21ai_1 _19744_ (.B1(_03621_),
    .Y(_02361_),
    .A1(net141),
    .A2(net83));
 sg13g2_nand2_1 _19745_ (.Y(_03622_),
    .A(\top_ihp.oisc.regs[8][28] ),
    .B(_03614_));
 sg13g2_o21ai_1 _19746_ (.B1(_03622_),
    .Y(_02362_),
    .A1(net63),
    .A2(net83));
 sg13g2_nand2_1 _19747_ (.Y(_03623_),
    .A(\top_ihp.oisc.regs[8][29] ),
    .B(net155));
 sg13g2_o21ai_1 _19748_ (.B1(_03623_),
    .Y(_02363_),
    .A1(net133),
    .A2(_03611_));
 sg13g2_nand2_1 _19749_ (.Y(_03624_),
    .A(\top_ihp.oisc.regs[8][2] ),
    .B(net155));
 sg13g2_o21ai_1 _19750_ (.B1(_03624_),
    .Y(_02364_),
    .A1(net222),
    .A2(net83));
 sg13g2_nand2_1 _19751_ (.Y(_03625_),
    .A(\top_ihp.oisc.regs[8][30] ),
    .B(net155));
 sg13g2_o21ai_1 _19752_ (.B1(_03625_),
    .Y(_02365_),
    .A1(net62),
    .A2(_03599_));
 sg13g2_nand2_1 _19753_ (.Y(_03626_),
    .A(\top_ihp.oisc.regs[8][31] ),
    .B(net158));
 sg13g2_o21ai_1 _19754_ (.B1(_03626_),
    .Y(_02366_),
    .A1(net239),
    .A2(net157));
 sg13g2_nand2_1 _19755_ (.Y(_03627_),
    .A(\top_ihp.oisc.regs[8][3] ),
    .B(_03597_));
 sg13g2_o21ai_1 _19756_ (.B1(_03627_),
    .Y(_02367_),
    .A1(_10047_),
    .A2(net157));
 sg13g2_nand2_1 _19757_ (.Y(_03628_),
    .A(\top_ihp.oisc.regs[8][4] ),
    .B(_03597_));
 sg13g2_o21ai_1 _19758_ (.B1(_03628_),
    .Y(_02368_),
    .A1(_10048_),
    .A2(_03599_));
 sg13g2_nand2_1 _19759_ (.Y(_03629_),
    .A(\top_ihp.oisc.regs[8][5] ),
    .B(net158));
 sg13g2_o21ai_1 _19760_ (.B1(_03629_),
    .Y(_02369_),
    .A1(net212),
    .A2(net157));
 sg13g2_nand2_1 _19761_ (.Y(_03630_),
    .A(\top_ihp.oisc.regs[8][6] ),
    .B(net158));
 sg13g2_o21ai_1 _19762_ (.B1(_03630_),
    .Y(_02370_),
    .A1(net211),
    .A2(net157));
 sg13g2_nand2_1 _19763_ (.Y(_03631_),
    .A(\top_ihp.oisc.regs[8][7] ),
    .B(net158));
 sg13g2_o21ai_1 _19764_ (.B1(_03631_),
    .Y(_02371_),
    .A1(net47),
    .A2(net157));
 sg13g2_nand2_1 _19765_ (.Y(_03632_),
    .A(\top_ihp.oisc.regs[8][8] ),
    .B(net158));
 sg13g2_o21ai_1 _19766_ (.B1(_03632_),
    .Y(_02372_),
    .A1(net61),
    .A2(net157));
 sg13g2_nand2_1 _19767_ (.Y(_03633_),
    .A(\top_ihp.oisc.regs[8][9] ),
    .B(net158));
 sg13g2_o21ai_1 _19768_ (.B1(_03633_),
    .Y(_02373_),
    .A1(net60),
    .A2(net157));
 sg13g2_nand3b_1 _19769_ (.B(_03317_),
    .C(_09083_),
    .Y(_03634_),
    .A_N(_09956_));
 sg13g2_buf_1 _19770_ (.A(_03634_),
    .X(_03635_));
 sg13g2_buf_2 _19771_ (.A(_03635_),
    .X(_03636_));
 sg13g2_mux2_1 _19772_ (.A0(net407),
    .A1(\top_ihp.oisc.regs[9][0] ),
    .S(_03636_),
    .X(_02374_));
 sg13g2_nand2_1 _19773_ (.Y(_03637_),
    .A(net545),
    .B(_03317_));
 sg13g2_buf_2 _19774_ (.A(_03637_),
    .X(_03638_));
 sg13g2_buf_8 _19775_ (.A(_03638_),
    .X(_03639_));
 sg13g2_nand2_1 _19776_ (.Y(_03640_),
    .A(\top_ihp.oisc.regs[9][10] ),
    .B(net276));
 sg13g2_o21ai_1 _19777_ (.B1(_03640_),
    .Y(_02375_),
    .A1(net65),
    .A2(net82));
 sg13g2_nand2_1 _19778_ (.Y(_03641_),
    .A(\top_ihp.oisc.regs[9][11] ),
    .B(net276));
 sg13g2_o21ai_1 _19779_ (.B1(_03641_),
    .Y(_02376_),
    .A1(_09303_),
    .A2(net82));
 sg13g2_nand2_1 _19780_ (.Y(_03642_),
    .A(\top_ihp.oisc.regs[9][12] ),
    .B(net276));
 sg13g2_o21ai_1 _19781_ (.B1(_03642_),
    .Y(_02377_),
    .A1(net218),
    .A2(net82));
 sg13g2_nor2_1 _19782_ (.A(_09958_),
    .B(_10093_),
    .Y(_03643_));
 sg13g2_buf_2 _19783_ (.A(_03643_),
    .X(_03644_));
 sg13g2_nor2_1 _19784_ (.A(\top_ihp.oisc.regs[9][13] ),
    .B(_03644_),
    .Y(_03645_));
 sg13g2_a21oi_1 _19785_ (.A1(net73),
    .A2(_03644_),
    .Y(_02378_),
    .B1(_03645_));
 sg13g2_nand2_1 _19786_ (.Y(_03646_),
    .A(\top_ihp.oisc.regs[9][14] ),
    .B(net276));
 sg13g2_o21ai_1 _19787_ (.B1(_03646_),
    .Y(_02379_),
    .A1(net217),
    .A2(net82));
 sg13g2_nand2_1 _19788_ (.Y(_03647_),
    .A(\top_ihp.oisc.regs[9][15] ),
    .B(net276));
 sg13g2_o21ai_1 _19789_ (.B1(_03647_),
    .Y(_02380_),
    .A1(net216),
    .A2(net82));
 sg13g2_nor2_1 _19790_ (.A(\top_ihp.oisc.regs[9][16] ),
    .B(_03644_),
    .Y(_03648_));
 sg13g2_a21oi_1 _19791_ (.A1(net146),
    .A2(_03644_),
    .Y(_02381_),
    .B1(_03648_));
 sg13g2_nand2_1 _19792_ (.Y(_03649_),
    .A(\top_ihp.oisc.regs[9][17] ),
    .B(net276));
 sg13g2_o21ai_1 _19793_ (.B1(_03649_),
    .Y(_02382_),
    .A1(net136),
    .A2(net82));
 sg13g2_nand2_1 _19794_ (.Y(_03650_),
    .A(\top_ihp.oisc.regs[9][18] ),
    .B(_03636_));
 sg13g2_o21ai_1 _19795_ (.B1(_03650_),
    .Y(_02383_),
    .A1(net135),
    .A2(net82));
 sg13g2_buf_1 _19796_ (.A(_03635_),
    .X(_03651_));
 sg13g2_nand2_1 _19797_ (.Y(_03652_),
    .A(\top_ihp.oisc.regs[9][19] ),
    .B(net275));
 sg13g2_o21ai_1 _19798_ (.B1(_03652_),
    .Y(_02384_),
    .A1(net215),
    .A2(_03639_));
 sg13g2_nand2_1 _19799_ (.Y(_03653_),
    .A(\top_ihp.oisc.regs[9][1] ),
    .B(net275));
 sg13g2_o21ai_1 _19800_ (.B1(_03653_),
    .Y(_02385_),
    .A1(net547),
    .A2(net82));
 sg13g2_nand2_1 _19801_ (.Y(_03654_),
    .A(\top_ihp.oisc.regs[9][20] ),
    .B(net275));
 sg13g2_o21ai_1 _19802_ (.B1(_03654_),
    .Y(_02386_),
    .A1(_09563_),
    .A2(net276));
 sg13g2_nand2_1 _19803_ (.Y(_03655_),
    .A(\top_ihp.oisc.regs[9][21] ),
    .B(net275));
 sg13g2_o21ai_1 _19804_ (.B1(_03655_),
    .Y(_02387_),
    .A1(net64),
    .A2(_03639_));
 sg13g2_nor2_1 _19805_ (.A(\top_ihp.oisc.regs[9][22] ),
    .B(_03644_),
    .Y(_03656_));
 sg13g2_a21oi_1 _19806_ (.A1(net143),
    .A2(_03644_),
    .Y(_02388_),
    .B1(_03656_));
 sg13g2_nor2_1 _19807_ (.A(\top_ihp.oisc.regs[9][23] ),
    .B(_03644_),
    .Y(_03657_));
 sg13g2_a21oi_1 _19808_ (.A1(net243),
    .A2(_03644_),
    .Y(_02389_),
    .B1(_03657_));
 sg13g2_buf_1 _19809_ (.A(_03638_),
    .X(_03658_));
 sg13g2_nand2_1 _19810_ (.Y(_03659_),
    .A(\top_ihp.oisc.regs[9][24] ),
    .B(net275));
 sg13g2_o21ai_1 _19811_ (.B1(_03659_),
    .Y(_02390_),
    .A1(net214),
    .A2(net81));
 sg13g2_nand2_1 _19812_ (.Y(_03660_),
    .A(\top_ihp.oisc.regs[9][25] ),
    .B(net275));
 sg13g2_o21ai_1 _19813_ (.B1(_03660_),
    .Y(_02391_),
    .A1(net213),
    .A2(net81));
 sg13g2_nand2_1 _19814_ (.Y(_03661_),
    .A(\top_ihp.oisc.regs[9][26] ),
    .B(_03651_));
 sg13g2_o21ai_1 _19815_ (.B1(_03661_),
    .Y(_02392_),
    .A1(net134),
    .A2(net81));
 sg13g2_nand2_1 _19816_ (.Y(_03662_),
    .A(\top_ihp.oisc.regs[9][27] ),
    .B(net275));
 sg13g2_o21ai_1 _19817_ (.B1(_03662_),
    .Y(_02393_),
    .A1(net141),
    .A2(net81));
 sg13g2_nand2_1 _19818_ (.Y(_03663_),
    .A(\top_ihp.oisc.regs[9][28] ),
    .B(net275));
 sg13g2_o21ai_1 _19819_ (.B1(_03663_),
    .Y(_02394_),
    .A1(net63),
    .A2(net81));
 sg13g2_nand2_1 _19820_ (.Y(_03664_),
    .A(\top_ihp.oisc.regs[9][29] ),
    .B(_03651_));
 sg13g2_o21ai_1 _19821_ (.B1(_03664_),
    .Y(_02395_),
    .A1(net133),
    .A2(_03658_));
 sg13g2_buf_1 _19822_ (.A(_03635_),
    .X(_03665_));
 sg13g2_nand2_1 _19823_ (.Y(_03666_),
    .A(\top_ihp.oisc.regs[9][2] ),
    .B(net274));
 sg13g2_o21ai_1 _19824_ (.B1(_03666_),
    .Y(_02396_),
    .A1(net222),
    .A2(_03658_));
 sg13g2_nand2_1 _19825_ (.Y(_03667_),
    .A(\top_ihp.oisc.regs[9][30] ),
    .B(net274));
 sg13g2_o21ai_1 _19826_ (.B1(_03667_),
    .Y(_02397_),
    .A1(net62),
    .A2(net81));
 sg13g2_nand2_1 _19827_ (.Y(_03668_),
    .A(\top_ihp.oisc.regs[9][31] ),
    .B(_03665_));
 sg13g2_o21ai_1 _19828_ (.B1(_03668_),
    .Y(_02398_),
    .A1(net239),
    .A2(net81));
 sg13g2_nand2_1 _19829_ (.Y(_03669_),
    .A(\top_ihp.oisc.regs[9][3] ),
    .B(_03665_));
 sg13g2_o21ai_1 _19830_ (.B1(_03669_),
    .Y(_02399_),
    .A1(net221),
    .A2(net81));
 sg13g2_nand2_1 _19831_ (.Y(_03670_),
    .A(\top_ihp.oisc.regs[9][4] ),
    .B(net274));
 sg13g2_o21ai_1 _19832_ (.B1(_03670_),
    .Y(_02400_),
    .A1(net220),
    .A2(_03638_));
 sg13g2_nand2_1 _19833_ (.Y(_03671_),
    .A(\top_ihp.oisc.regs[9][5] ),
    .B(net274));
 sg13g2_o21ai_1 _19834_ (.B1(_03671_),
    .Y(_02401_),
    .A1(net212),
    .A2(_03638_));
 sg13g2_nand2_1 _19835_ (.Y(_03672_),
    .A(\top_ihp.oisc.regs[9][6] ),
    .B(net274));
 sg13g2_o21ai_1 _19836_ (.B1(_03672_),
    .Y(_02402_),
    .A1(net211),
    .A2(_03638_));
 sg13g2_nand2_1 _19837_ (.Y(_03673_),
    .A(\top_ihp.oisc.regs[9][7] ),
    .B(net274));
 sg13g2_o21ai_1 _19838_ (.B1(_03673_),
    .Y(_02403_),
    .A1(net408),
    .A2(net276));
 sg13g2_nand2_1 _19839_ (.Y(_03674_),
    .A(\top_ihp.oisc.regs[9][8] ),
    .B(net274));
 sg13g2_o21ai_1 _19840_ (.B1(_03674_),
    .Y(_02404_),
    .A1(net61),
    .A2(_03638_));
 sg13g2_nand2_1 _19841_ (.Y(_03675_),
    .A(\top_ihp.oisc.regs[9][9] ),
    .B(net274));
 sg13g2_o21ai_1 _19842_ (.B1(_03675_),
    .Y(_02405_),
    .A1(net60),
    .A2(_03638_));
 sg13g2_a21oi_1 _19843_ (.A1(_07419_),
    .A2(net823),
    .Y(_03676_),
    .B1(_07420_));
 sg13g2_nand2_1 _19844_ (.Y(_03677_),
    .A(net879),
    .B(_03676_));
 sg13g2_o21ai_1 _19845_ (.B1(_03677_),
    .Y(_03678_),
    .A1(_13205_),
    .A2(_07436_));
 sg13g2_nand2_1 _19846_ (.Y(_03679_),
    .A(net1017),
    .B(net823));
 sg13g2_buf_1 _19847_ (.A(_03679_),
    .X(_03680_));
 sg13g2_inv_1 _19848_ (.Y(_03681_),
    .A(_08241_));
 sg13g2_a221oi_1 _19849_ (.B2(_03681_),
    .C1(net979),
    .B1(_03680_),
    .A1(_13205_),
    .Y(_03682_),
    .A2(net823));
 sg13g2_a21oi_1 _19850_ (.A1(net979),
    .A2(_03678_),
    .Y(_02406_),
    .B1(_03682_));
 sg13g2_buf_1 _19851_ (.A(_07678_),
    .X(_03683_));
 sg13g2_buf_1 _19852_ (.A(_00069_),
    .X(_03684_));
 sg13g2_nand3_1 _19853_ (.B(_03684_),
    .C(net774),
    .A(_09090_),
    .Y(_03685_));
 sg13g2_nor2_1 _19854_ (.A(_08237_),
    .B(_03685_),
    .Y(_03686_));
 sg13g2_a21oi_1 _19855_ (.A1(_03683_),
    .A2(_08237_),
    .Y(_03687_),
    .B1(_03686_));
 sg13g2_nor2_1 _19856_ (.A(net940),
    .B(net845),
    .Y(_03688_));
 sg13g2_buf_1 _19857_ (.A(_03688_),
    .X(_03689_));
 sg13g2_buf_2 _19858_ (.A(_03689_),
    .X(_03690_));
 sg13g2_buf_1 _19859_ (.A(net772),
    .X(_03691_));
 sg13g2_buf_1 _19860_ (.A(net735),
    .X(_03692_));
 sg13g2_nor2_1 _19861_ (.A(net979),
    .B(_03692_),
    .Y(_03693_));
 sg13g2_a22oi_1 _19862_ (.Y(_02407_),
    .B1(_03693_),
    .B2(_03685_),
    .A2(_03687_),
    .A1(net979));
 sg13g2_nand2_1 _19863_ (.Y(_03694_),
    .A(net1016),
    .B(_08237_));
 sg13g2_o21ai_1 _19864_ (.B1(_03694_),
    .Y(_03695_),
    .A1(_07423_),
    .A2(net774));
 sg13g2_nor2_1 _19865_ (.A(_07648_),
    .B(_08244_),
    .Y(_03696_));
 sg13g2_buf_1 _19866_ (.A(_03696_),
    .X(_03697_));
 sg13g2_nand2_1 _19867_ (.Y(_03698_),
    .A(_03684_),
    .B(_03697_));
 sg13g2_nand2_1 _19868_ (.Y(_03699_),
    .A(net998),
    .B(_03695_));
 sg13g2_o21ai_1 _19869_ (.B1(_03699_),
    .Y(_02408_),
    .A1(_03695_),
    .A2(_03698_));
 sg13g2_nand2_1 _19870_ (.Y(_03700_),
    .A(net999),
    .B(_08250_));
 sg13g2_nand3_1 _19871_ (.B(_03684_),
    .C(net774),
    .A(net998),
    .Y(_03701_));
 sg13g2_o21ai_1 _19872_ (.B1(_03701_),
    .Y(_03702_),
    .A1(_08992_),
    .A2(net774));
 sg13g2_nand2b_1 _19873_ (.Y(_03703_),
    .B(_03702_),
    .A_N(_08247_));
 sg13g2_nand4_1 _19874_ (.B(_03684_),
    .C(net879),
    .A(net998),
    .Y(_03704_),
    .D(net774));
 sg13g2_nand3_1 _19875_ (.B(_03703_),
    .C(_03704_),
    .A(_03700_),
    .Y(_02409_));
 sg13g2_nand2_1 _19876_ (.Y(_03705_),
    .A(_09294_),
    .B(_08250_));
 sg13g2_nand3_1 _19877_ (.B(_03684_),
    .C(net774),
    .A(_08944_),
    .Y(_03706_));
 sg13g2_o21ai_1 _19878_ (.B1(_03706_),
    .Y(_03707_),
    .A1(_09122_),
    .A2(net774));
 sg13g2_nand2b_1 _19879_ (.Y(_03708_),
    .B(_03707_),
    .A_N(_08247_));
 sg13g2_nand4_1 _19880_ (.B(_03684_),
    .C(net879),
    .A(_08944_),
    .Y(_03709_),
    .D(_08246_));
 sg13g2_nand3_1 _19881_ (.B(_03708_),
    .C(_03709_),
    .A(_03705_),
    .Y(_02410_));
 sg13g2_o21ai_1 _19882_ (.B1(_03694_),
    .Y(_03710_),
    .A1(net1016),
    .A2(net845));
 sg13g2_nand2_1 _19883_ (.Y(_03711_),
    .A(_08241_),
    .B(_03710_));
 sg13g2_o21ai_1 _19884_ (.B1(_03711_),
    .Y(_02411_),
    .A1(_07654_),
    .A2(_03676_));
 sg13g2_buf_2 _19885_ (.A(\top_ihp.oisc.wb_dat_o[0] ),
    .X(_03712_));
 sg13g2_nand2_1 _19886_ (.Y(_03713_),
    .A(_07419_),
    .B(_08943_));
 sg13g2_buf_1 _19887_ (.A(_03713_),
    .X(_03714_));
 sg13g2_buf_1 _19888_ (.A(_03714_),
    .X(_03715_));
 sg13g2_mux2_1 _19889_ (.A0(net407),
    .A1(_03712_),
    .S(_03715_),
    .X(_02412_));
 sg13g2_buf_1 _19890_ (.A(_03714_),
    .X(_03716_));
 sg13g2_buf_1 _19891_ (.A(net910),
    .X(_03717_));
 sg13g2_buf_1 _19892_ (.A(\top_ihp.oisc.wb_dat_o[10] ),
    .X(_03718_));
 sg13g2_buf_1 _19893_ (.A(_03714_),
    .X(_03719_));
 sg13g2_nand2_1 _19894_ (.Y(_03720_),
    .A(_03718_),
    .B(net909));
 sg13g2_o21ai_1 _19895_ (.B1(_03720_),
    .Y(_02413_),
    .A1(net65),
    .A2(net881));
 sg13g2_buf_1 _19896_ (.A(\top_ihp.oisc.wb_dat_o[11] ),
    .X(_03721_));
 sg13g2_nand2_1 _19897_ (.Y(_03722_),
    .A(_03721_),
    .B(net909));
 sg13g2_o21ai_1 _19898_ (.B1(_03722_),
    .Y(_02414_),
    .A1(net251),
    .A2(net881));
 sg13g2_buf_1 _19899_ (.A(\top_ihp.oisc.wb_dat_o[12] ),
    .X(_03723_));
 sg13g2_nand2_1 _19900_ (.Y(_03724_),
    .A(_03723_),
    .B(net909));
 sg13g2_o21ai_1 _19901_ (.B1(_03724_),
    .Y(_02415_),
    .A1(net218),
    .A2(net881));
 sg13g2_buf_1 _19902_ (.A(\top_ihp.oisc.wb_dat_o[13] ),
    .X(_03725_));
 sg13g2_nand2_1 _19903_ (.Y(_03726_),
    .A(_03725_),
    .B(net909));
 sg13g2_o21ai_1 _19904_ (.B1(_03726_),
    .Y(_02416_),
    .A1(net147),
    .A2(net881));
 sg13g2_buf_1 _19905_ (.A(\top_ihp.oisc.wb_dat_o[14] ),
    .X(_03727_));
 sg13g2_mux2_1 _19906_ (.A0(_07521_),
    .A1(_03727_),
    .S(net911),
    .X(_02417_));
 sg13g2_buf_1 _19907_ (.A(\top_ihp.oisc.wb_dat_o[15] ),
    .X(_03728_));
 sg13g2_nand2_1 _19908_ (.Y(_03729_),
    .A(_03728_),
    .B(net909));
 sg13g2_o21ai_1 _19909_ (.B1(_03729_),
    .Y(_02418_),
    .A1(_10068_),
    .A2(net881));
 sg13g2_nand2_1 _19910_ (.Y(_03730_),
    .A(\top_ihp.oisc.wb_dat_o[16] ),
    .B(_03719_));
 sg13g2_o21ai_1 _19911_ (.B1(_03730_),
    .Y(_02419_),
    .A1(_09436_),
    .A2(net881));
 sg13g2_nand2_1 _19912_ (.Y(_03731_),
    .A(\top_ihp.oisc.wb_dat_o[17] ),
    .B(_03719_));
 sg13g2_o21ai_1 _19913_ (.B1(_03731_),
    .Y(_02420_),
    .A1(net136),
    .A2(net881));
 sg13g2_nand2_1 _19914_ (.Y(_03732_),
    .A(\top_ihp.oisc.wb_dat_o[18] ),
    .B(net909));
 sg13g2_o21ai_1 _19915_ (.B1(_03732_),
    .Y(_02421_),
    .A1(_10071_),
    .A2(net881));
 sg13g2_buf_1 _19916_ (.A(_03714_),
    .X(_03733_));
 sg13g2_nand2_1 _19917_ (.Y(_03734_),
    .A(\top_ihp.oisc.wb_dat_o[19] ),
    .B(net908));
 sg13g2_o21ai_1 _19918_ (.B1(_03734_),
    .Y(_02422_),
    .A1(_09557_),
    .A2(_03717_));
 sg13g2_buf_1 _19919_ (.A(\top_ihp.oisc.wb_dat_o[1] ),
    .X(_03735_));
 sg13g2_nand2_1 _19920_ (.Y(_03736_),
    .A(_03735_),
    .B(_03733_));
 sg13g2_o21ai_1 _19921_ (.B1(_03736_),
    .Y(_02423_),
    .A1(net547),
    .A2(_03717_));
 sg13g2_buf_1 _19922_ (.A(net910),
    .X(_03737_));
 sg13g2_nand2_1 _19923_ (.Y(_03738_),
    .A(\top_ihp.oisc.wb_dat_o[20] ),
    .B(net908));
 sg13g2_o21ai_1 _19924_ (.B1(_03738_),
    .Y(_02424_),
    .A1(_09556_),
    .A2(_03737_));
 sg13g2_nand2_1 _19925_ (.Y(_03739_),
    .A(\top_ihp.oisc.wb_dat_o[21] ),
    .B(net908));
 sg13g2_o21ai_1 _19926_ (.B1(_03739_),
    .Y(_02425_),
    .A1(net64),
    .A2(net880));
 sg13g2_nand2_1 _19927_ (.Y(_03740_),
    .A(\top_ihp.oisc.wb_dat_o[22] ),
    .B(net908));
 sg13g2_o21ai_1 _19928_ (.B1(_03740_),
    .Y(_02426_),
    .A1(_07801_),
    .A2(net880));
 sg13g2_mux2_1 _19929_ (.A0(_07442_),
    .A1(\top_ihp.oisc.wb_dat_o[23] ),
    .S(_03715_),
    .X(_02427_));
 sg13g2_nand2_1 _19930_ (.Y(_03741_),
    .A(\top_ihp.oisc.wb_dat_o[24] ),
    .B(net908));
 sg13g2_o21ai_1 _19931_ (.B1(_03741_),
    .Y(_02428_),
    .A1(net214),
    .A2(net880));
 sg13g2_nand2_1 _19932_ (.Y(_03742_),
    .A(\top_ihp.oisc.wb_dat_o[25] ),
    .B(net908));
 sg13g2_o21ai_1 _19933_ (.B1(_03742_),
    .Y(_02429_),
    .A1(net213),
    .A2(net880));
 sg13g2_nand2_1 _19934_ (.Y(_03743_),
    .A(\top_ihp.oisc.wb_dat_o[26] ),
    .B(net908));
 sg13g2_o21ai_1 _19935_ (.B1(_03743_),
    .Y(_02430_),
    .A1(net134),
    .A2(net880));
 sg13g2_mux2_1 _19936_ (.A0(_07681_),
    .A1(\top_ihp.oisc.wb_dat_o[27] ),
    .S(net911),
    .X(_02431_));
 sg13g2_nand2_1 _19937_ (.Y(_03744_),
    .A(\top_ihp.oisc.wb_dat_o[28] ),
    .B(net908));
 sg13g2_o21ai_1 _19938_ (.B1(_03744_),
    .Y(_02432_),
    .A1(net63),
    .A2(net880));
 sg13g2_mux2_1 _19939_ (.A0(_07721_),
    .A1(\top_ihp.oisc.wb_dat_o[29] ),
    .S(net909),
    .X(_02433_));
 sg13g2_buf_1 _19940_ (.A(\top_ihp.oisc.wb_dat_o[2] ),
    .X(_03745_));
 sg13g2_nand2_1 _19941_ (.Y(_03746_),
    .A(_03745_),
    .B(_03733_));
 sg13g2_o21ai_1 _19942_ (.B1(_03746_),
    .Y(_02434_),
    .A1(net222),
    .A2(_03737_));
 sg13g2_nand2_1 _19943_ (.Y(_03747_),
    .A(\top_ihp.oisc.wb_dat_o[30] ),
    .B(net910));
 sg13g2_o21ai_1 _19944_ (.B1(_03747_),
    .Y(_02435_),
    .A1(net62),
    .A2(net880));
 sg13g2_mux2_1 _19945_ (.A0(_08946_),
    .A1(\top_ihp.oisc.wb_dat_o[31] ),
    .S(net909),
    .X(_02436_));
 sg13g2_buf_1 _19946_ (.A(\top_ihp.oisc.wb_dat_o[3] ),
    .X(_03748_));
 sg13g2_nand2_1 _19947_ (.Y(_03749_),
    .A(_03748_),
    .B(net910));
 sg13g2_o21ai_1 _19948_ (.B1(_03749_),
    .Y(_02437_),
    .A1(net221),
    .A2(net880));
 sg13g2_buf_1 _19949_ (.A(\top_ihp.oisc.wb_dat_o[4] ),
    .X(_03750_));
 sg13g2_nand2_1 _19950_ (.Y(_03751_),
    .A(_03750_),
    .B(_03716_));
 sg13g2_o21ai_1 _19951_ (.B1(_03751_),
    .Y(_02438_),
    .A1(net220),
    .A2(net911));
 sg13g2_buf_1 _19952_ (.A(\top_ihp.oisc.wb_dat_o[5] ),
    .X(_03752_));
 sg13g2_nand2_1 _19953_ (.Y(_03753_),
    .A(_03752_),
    .B(_03716_));
 sg13g2_o21ai_1 _19954_ (.B1(_03753_),
    .Y(_02439_),
    .A1(net212),
    .A2(net911));
 sg13g2_buf_1 _19955_ (.A(\top_ihp.oisc.wb_dat_o[6] ),
    .X(_03754_));
 sg13g2_nand2_1 _19956_ (.Y(_03755_),
    .A(_03754_),
    .B(net910));
 sg13g2_o21ai_1 _19957_ (.B1(_03755_),
    .Y(_02440_),
    .A1(net211),
    .A2(net911));
 sg13g2_buf_1 _19958_ (.A(\top_ihp.oisc.wb_dat_o[7] ),
    .X(_03756_));
 sg13g2_nand2_1 _19959_ (.Y(_03757_),
    .A(_03756_),
    .B(net910));
 sg13g2_o21ai_1 _19960_ (.B1(_03757_),
    .Y(_02441_),
    .A1(_09911_),
    .A2(net911));
 sg13g2_buf_1 _19961_ (.A(\top_ihp.oisc.wb_dat_o[8] ),
    .X(_03758_));
 sg13g2_nand2_1 _19962_ (.Y(_03759_),
    .A(_03758_),
    .B(net910));
 sg13g2_o21ai_1 _19963_ (.B1(_03759_),
    .Y(_02442_),
    .A1(net61),
    .A2(net911));
 sg13g2_buf_1 _19964_ (.A(\top_ihp.oisc.wb_dat_o[9] ),
    .X(_03760_));
 sg13g2_nand2_1 _19965_ (.Y(_03761_),
    .A(_03760_),
    .B(net910));
 sg13g2_o21ai_1 _19966_ (.B1(_03761_),
    .Y(_02443_),
    .A1(net60),
    .A2(net911));
 sg13g2_inv_1 _19967_ (.Y(_03762_),
    .A(_00138_));
 sg13g2_nand2_2 _19968_ (.Y(_03763_),
    .A(_08181_),
    .B(_08182_));
 sg13g2_nand2b_1 _19969_ (.Y(_03764_),
    .B(net869),
    .A_N(_03763_));
 sg13g2_buf_2 _19970_ (.A(_03764_),
    .X(_03765_));
 sg13g2_buf_1 _19971_ (.A(\top_ihp.wb_emem.bit_counter[0] ),
    .X(_03766_));
 sg13g2_nand3_1 _19972_ (.B(net868),
    .C(_03765_),
    .A(_03766_),
    .Y(_03767_));
 sg13g2_o21ai_1 _19973_ (.B1(_03767_),
    .Y(_02444_),
    .A1(_03762_),
    .A2(_03765_));
 sg13g2_buf_1 _19974_ (.A(\top_ihp.wb_emem.bit_counter[1] ),
    .X(_03768_));
 sg13g2_nor2_2 _19975_ (.A(_08188_),
    .B(_03763_),
    .Y(_03769_));
 sg13g2_nand2_1 _19976_ (.Y(_03770_),
    .A(_03766_),
    .B(_03769_));
 sg13g2_nor2_2 _19977_ (.A(_08184_),
    .B(_03769_),
    .Y(_03771_));
 sg13g2_nor2_1 _19978_ (.A(_03766_),
    .B(_03765_),
    .Y(_03772_));
 sg13g2_o21ai_1 _19979_ (.B1(_03768_),
    .Y(_03773_),
    .A1(_03771_),
    .A2(_03772_));
 sg13g2_o21ai_1 _19980_ (.B1(_03773_),
    .Y(_02445_),
    .A1(_03768_),
    .A2(_03770_));
 sg13g2_nand2_1 _19981_ (.Y(_03774_),
    .A(_03768_),
    .B(_03766_));
 sg13g2_xor2_1 _19982_ (.B(_03774_),
    .A(\top_ihp.wb_emem.bit_counter[2] ),
    .X(_03775_));
 sg13g2_nand3_1 _19983_ (.B(net868),
    .C(_03765_),
    .A(\top_ihp.wb_emem.bit_counter[2] ),
    .Y(_03776_));
 sg13g2_o21ai_1 _19984_ (.B1(_03776_),
    .Y(_02446_),
    .A1(_03765_),
    .A2(_03775_));
 sg13g2_buf_2 _19985_ (.A(\top_ihp.wb_emem.bit_counter[3] ),
    .X(_03777_));
 sg13g2_and3_1 _19986_ (.X(_03778_),
    .A(_03768_),
    .B(_03766_),
    .C(\top_ihp.wb_emem.bit_counter[2] ));
 sg13g2_buf_1 _19987_ (.A(_03778_),
    .X(_03779_));
 sg13g2_nand2_1 _19988_ (.Y(_03780_),
    .A(_03769_),
    .B(_03779_));
 sg13g2_nor2_1 _19989_ (.A(_03765_),
    .B(_03779_),
    .Y(_03781_));
 sg13g2_o21ai_1 _19990_ (.B1(_03777_),
    .Y(_03782_),
    .A1(_03771_),
    .A2(_03781_));
 sg13g2_o21ai_1 _19991_ (.B1(_03782_),
    .Y(_02447_),
    .A1(_03777_),
    .A2(_03780_));
 sg13g2_buf_1 _19992_ (.A(\top_ihp.wb_emem.bit_counter[4] ),
    .X(_03783_));
 sg13g2_nand3_1 _19993_ (.B(_03769_),
    .C(_03779_),
    .A(_03777_),
    .Y(_03784_));
 sg13g2_a21oi_1 _19994_ (.A1(_03777_),
    .A2(_03779_),
    .Y(_03785_),
    .B1(_03765_));
 sg13g2_o21ai_1 _19995_ (.B1(_03783_),
    .Y(_03786_),
    .A1(_03771_),
    .A2(_03785_));
 sg13g2_o21ai_1 _19996_ (.B1(_03786_),
    .Y(_02448_),
    .A1(_03783_),
    .A2(_03784_));
 sg13g2_inv_1 _19997_ (.Y(_03787_),
    .A(_03783_));
 sg13g2_nor2_1 _19998_ (.A(_03787_),
    .B(_03784_),
    .Y(_03788_));
 sg13g2_nand3_1 _19999_ (.B(_03783_),
    .C(_03779_),
    .A(_03777_),
    .Y(_03789_));
 sg13g2_a21o_1 _20000_ (.A2(_03789_),
    .A1(_03769_),
    .B1(_03771_),
    .X(_03790_));
 sg13g2_buf_1 _20001_ (.A(\top_ihp.wb_emem.bit_counter[5] ),
    .X(_03791_));
 sg13g2_mux2_1 _20002_ (.A0(_03788_),
    .A1(_03790_),
    .S(_03791_),
    .X(_02449_));
 sg13g2_buf_1 _20003_ (.A(\top_ihp.wb_emem.bit_counter[6] ),
    .X(_03792_));
 sg13g2_nand2_1 _20004_ (.Y(_03793_),
    .A(_03791_),
    .B(_03788_));
 sg13g2_xor2_1 _20005_ (.B(_03793_),
    .A(_03792_),
    .X(_03794_));
 sg13g2_nor2_1 _20006_ (.A(_08184_),
    .B(_03794_),
    .Y(_02450_));
 sg13g2_nand2_1 _20007_ (.Y(_03795_),
    .A(\top_ihp.wb_emem.bit_counter[7] ),
    .B(net868));
 sg13g2_nand3_1 _20008_ (.B(_03792_),
    .C(_03788_),
    .A(_03791_),
    .Y(_03796_));
 sg13g2_mux2_1 _20009_ (.A0(\top_ihp.wb_emem.bit_counter[7] ),
    .A1(_03795_),
    .S(_03796_),
    .X(_03797_));
 sg13g2_inv_1 _20010_ (.Y(_02451_),
    .A(_03797_));
 sg13g2_inv_1 _20011_ (.Y(_03798_),
    .A(_08182_));
 sg13g2_a21oi_1 _20012_ (.A1(_03798_),
    .A2(_08188_),
    .Y(_03799_),
    .B1(_08181_));
 sg13g2_buf_1 _20013_ (.A(_03799_),
    .X(_03800_));
 sg13g2_buf_1 _20014_ (.A(_03800_),
    .X(_03801_));
 sg13g2_buf_1 _20015_ (.A(_03801_),
    .X(_03802_));
 sg13g2_nand2_1 _20016_ (.Y(_03803_),
    .A(_08184_),
    .B(_08188_));
 sg13g2_buf_1 _20017_ (.A(_03803_),
    .X(_03804_));
 sg13g2_buf_1 _20018_ (.A(net866),
    .X(_03805_));
 sg13g2_nand2_1 _20019_ (.Y(_03806_),
    .A(net3),
    .B(net858));
 sg13g2_buf_1 _20020_ (.A(_07656_),
    .X(_03807_));
 sg13g2_nor2_1 _20021_ (.A(_09337_),
    .B(net869),
    .Y(_03808_));
 sg13g2_buf_1 _20022_ (.A(_03808_),
    .X(_03809_));
 sg13g2_buf_1 _20023_ (.A(net837),
    .X(_03810_));
 sg13g2_nand3_1 _20024_ (.B(net820),
    .C(net819),
    .A(\top_ihp.oisc.wb_dat_o[24] ),
    .Y(_03811_));
 sg13g2_buf_1 _20025_ (.A(_03800_),
    .X(_03812_));
 sg13g2_a21oi_1 _20026_ (.A1(_03806_),
    .A2(_03811_),
    .Y(_03813_),
    .B1(net857));
 sg13g2_a21o_1 _20027_ (.A2(_03802_),
    .A1(\top_ihp.wb_dati_ram[24] ),
    .B1(_03813_),
    .X(_02452_));
 sg13g2_buf_1 _20028_ (.A(_03801_),
    .X(_03814_));
 sg13g2_buf_1 _20029_ (.A(net866),
    .X(_03815_));
 sg13g2_buf_1 _20030_ (.A(net837),
    .X(_03816_));
 sg13g2_and2_1 _20031_ (.A(\top_ihp.oisc.wb_dat_o[18] ),
    .B(net818),
    .X(_03817_));
 sg13g2_buf_1 _20032_ (.A(_03800_),
    .X(_03818_));
 sg13g2_a221oi_1 _20033_ (.B2(net806),
    .C1(_03818_),
    .B1(_03817_),
    .A1(\top_ihp.wb_dati_ram[17] ),
    .Y(_03819_),
    .A2(net856));
 sg13g2_a21oi_1 _20034_ (.A1(_09469_),
    .A2(net836),
    .Y(_02453_),
    .B1(_03819_));
 sg13g2_and2_1 _20035_ (.A(\top_ihp.oisc.wb_dat_o[19] ),
    .B(net818),
    .X(_03820_));
 sg13g2_buf_1 _20036_ (.A(_03800_),
    .X(_03821_));
 sg13g2_a221oi_1 _20037_ (.B2(net806),
    .C1(_03821_),
    .B1(_03820_),
    .A1(\top_ihp.wb_dati_ram[18] ),
    .Y(_03822_),
    .A2(_03815_));
 sg13g2_a21oi_1 _20038_ (.A1(_09496_),
    .A2(net836),
    .Y(_02454_),
    .B1(_03822_));
 sg13g2_and2_1 _20039_ (.A(\top_ihp.oisc.wb_dat_o[20] ),
    .B(net818),
    .X(_03823_));
 sg13g2_a221oi_1 _20040_ (.B2(net806),
    .C1(_03821_),
    .B1(_03823_),
    .A1(\top_ihp.wb_dati_ram[19] ),
    .Y(_03824_),
    .A2(_03815_));
 sg13g2_a21oi_1 _20041_ (.A1(_09566_),
    .A2(_03814_),
    .Y(_02455_),
    .B1(_03824_));
 sg13g2_nand2_1 _20042_ (.Y(_03825_),
    .A(\top_ihp.wb_dati_ram[20] ),
    .B(net858));
 sg13g2_nand3_1 _20043_ (.B(net820),
    .C(net819),
    .A(\top_ihp.oisc.wb_dat_o[21] ),
    .Y(_03826_));
 sg13g2_buf_1 _20044_ (.A(_03800_),
    .X(_03827_));
 sg13g2_a21oi_1 _20045_ (.A1(_03825_),
    .A2(_03826_),
    .Y(_03828_),
    .B1(net853));
 sg13g2_a21o_1 _20046_ (.A2(net838),
    .A1(\top_ihp.wb_dati_ram[21] ),
    .B1(_03828_),
    .X(_02456_));
 sg13g2_nand2_1 _20047_ (.Y(_03829_),
    .A(\top_ihp.wb_dati_ram[21] ),
    .B(net858));
 sg13g2_nand3_1 _20048_ (.B(net820),
    .C(net819),
    .A(\top_ihp.oisc.wb_dat_o[22] ),
    .Y(_03830_));
 sg13g2_a21oi_1 _20049_ (.A1(_03829_),
    .A2(_03830_),
    .Y(_03831_),
    .B1(net853));
 sg13g2_a21o_1 _20050_ (.A2(_03802_),
    .A1(\top_ihp.wb_dati_ram[22] ),
    .B1(_03831_),
    .X(_02457_));
 sg13g2_and2_1 _20051_ (.A(\top_ihp.oisc.wb_dat_o[23] ),
    .B(net818),
    .X(_03832_));
 sg13g2_a221oi_1 _20052_ (.B2(_07658_),
    .C1(net854),
    .B1(_03832_),
    .A1(\top_ihp.wb_dati_ram[22] ),
    .Y(_03833_),
    .A2(net856));
 sg13g2_a21oi_1 _20053_ (.A1(_09213_),
    .A2(_03814_),
    .Y(_02458_),
    .B1(_03833_));
 sg13g2_buf_1 _20054_ (.A(_03801_),
    .X(_03834_));
 sg13g2_nand2_1 _20055_ (.Y(_03835_),
    .A(\top_ihp.wb_dati_ram[23] ),
    .B(net858));
 sg13g2_nand3_1 _20056_ (.B(net824),
    .C(net819),
    .A(_03758_),
    .Y(_03836_));
 sg13g2_a21oi_1 _20057_ (.A1(_03835_),
    .A2(_03836_),
    .Y(_03837_),
    .B1(net853));
 sg13g2_a21o_1 _20058_ (.A2(net835),
    .A1(\top_ihp.wb_dati_ram[8] ),
    .B1(_03837_),
    .X(_02459_));
 sg13g2_nand2_1 _20059_ (.Y(_03838_),
    .A(\top_ihp.wb_dati_ram[8] ),
    .B(net858));
 sg13g2_nand3_1 _20060_ (.B(net824),
    .C(net819),
    .A(_03760_),
    .Y(_03839_));
 sg13g2_a21oi_1 _20061_ (.A1(_03838_),
    .A2(_03839_),
    .Y(_03840_),
    .B1(net853));
 sg13g2_a21o_1 _20062_ (.A2(net835),
    .A1(\top_ihp.wb_dati_ram[9] ),
    .B1(_03840_),
    .X(_02460_));
 sg13g2_buf_1 _20063_ (.A(net837),
    .X(_03841_));
 sg13g2_and2_1 _20064_ (.A(_03718_),
    .B(net817),
    .X(_03842_));
 sg13g2_buf_1 _20065_ (.A(net824),
    .X(_03843_));
 sg13g2_a221oi_1 _20066_ (.B2(net802),
    .C1(net854),
    .B1(_03842_),
    .A1(\top_ihp.wb_dati_ram[9] ),
    .Y(_03844_),
    .A2(net856));
 sg13g2_a21oi_1 _20067_ (.A1(_09249_),
    .A2(net836),
    .Y(_02461_),
    .B1(_03844_));
 sg13g2_inv_1 _20068_ (.Y(_03845_),
    .A(\top_ihp.wb_dati_ram[11] ));
 sg13g2_and2_1 _20069_ (.A(_03721_),
    .B(_03841_),
    .X(_03846_));
 sg13g2_a221oi_1 _20070_ (.B2(net802),
    .C1(net854),
    .B1(_03846_),
    .A1(\top_ihp.wb_dati_ram[10] ),
    .Y(_03847_),
    .A2(net856));
 sg13g2_a21oi_1 _20071_ (.A1(_03845_),
    .A2(net836),
    .Y(_02462_),
    .B1(_03847_));
 sg13g2_and2_1 _20072_ (.A(\top_ihp.oisc.wb_dat_o[25] ),
    .B(net817),
    .X(_03848_));
 sg13g2_a221oi_1 _20073_ (.B2(_03843_),
    .C1(net854),
    .B1(_03848_),
    .A1(\top_ihp.wb_dati_ram[24] ),
    .Y(_03849_),
    .A2(net856));
 sg13g2_a21oi_1 _20074_ (.A1(_09517_),
    .A2(net836),
    .Y(_02463_),
    .B1(_03849_));
 sg13g2_and2_1 _20075_ (.A(_03723_),
    .B(net817),
    .X(_03850_));
 sg13g2_a221oi_1 _20076_ (.B2(net802),
    .C1(net854),
    .B1(_03850_),
    .A1(\top_ihp.wb_dati_ram[11] ),
    .Y(_03851_),
    .A2(net856));
 sg13g2_a21oi_1 _20077_ (.A1(_09328_),
    .A2(net836),
    .Y(_02464_),
    .B1(_03851_));
 sg13g2_buf_1 _20078_ (.A(net866),
    .X(_03852_));
 sg13g2_and2_1 _20079_ (.A(_03725_),
    .B(_03841_),
    .X(_03853_));
 sg13g2_a221oi_1 _20080_ (.B2(_03843_),
    .C1(net854),
    .B1(_03853_),
    .A1(\top_ihp.wb_dati_ram[12] ),
    .Y(_03854_),
    .A2(net852));
 sg13g2_a21oi_1 _20081_ (.A1(_09354_),
    .A2(net836),
    .Y(_02465_),
    .B1(_03854_));
 sg13g2_and2_1 _20082_ (.A(_03727_),
    .B(net817),
    .X(_03855_));
 sg13g2_a221oi_1 _20083_ (.B2(net802),
    .C1(net854),
    .B1(_03855_),
    .A1(\top_ihp.wb_dati_ram[13] ),
    .Y(_03856_),
    .A2(net852));
 sg13g2_a21oi_1 _20084_ (.A1(_09379_),
    .A2(net836),
    .Y(_02466_),
    .B1(_03856_));
 sg13g2_buf_1 _20085_ (.A(_03801_),
    .X(_03857_));
 sg13g2_and2_1 _20086_ (.A(_03728_),
    .B(net817),
    .X(_03858_));
 sg13g2_a221oi_1 _20087_ (.B2(net802),
    .C1(net854),
    .B1(_03858_),
    .A1(\top_ihp.wb_dati_ram[14] ),
    .Y(_03859_),
    .A2(net852));
 sg13g2_a21oi_1 _20088_ (.A1(_08195_),
    .A2(_03857_),
    .Y(_02467_),
    .B1(_03859_));
 sg13g2_and2_1 _20089_ (.A(_03712_),
    .B(_03816_),
    .X(_03860_));
 sg13g2_a22oi_1 _20090_ (.Y(_03861_),
    .B1(_03860_),
    .B2(net806),
    .A2(net856),
    .A1(\top_ihp.wb_dati_ram[15] ));
 sg13g2_buf_1 _20091_ (.A(_03801_),
    .X(_03862_));
 sg13g2_nand2_1 _20092_ (.Y(_03863_),
    .A(\top_ihp.wb_dati_ram[0] ),
    .B(net833));
 sg13g2_o21ai_1 _20093_ (.B1(_03863_),
    .Y(_02468_),
    .A1(net838),
    .A2(_03861_));
 sg13g2_nand2_1 _20094_ (.Y(_03864_),
    .A(\top_ihp.wb_dati_ram[0] ),
    .B(_03805_));
 sg13g2_nand3_1 _20095_ (.B(net824),
    .C(net819),
    .A(_03735_),
    .Y(_03865_));
 sg13g2_a21oi_1 _20096_ (.A1(_03864_),
    .A2(_03865_),
    .Y(_03866_),
    .B1(net853));
 sg13g2_a21o_1 _20097_ (.A2(_03834_),
    .A1(\top_ihp.wb_dati_ram[1] ),
    .B1(_03866_),
    .X(_02469_));
 sg13g2_nand2_1 _20098_ (.Y(_03867_),
    .A(\top_ihp.wb_dati_ram[1] ),
    .B(net858));
 sg13g2_nand3_1 _20099_ (.B(net824),
    .C(net819),
    .A(_03745_),
    .Y(_03868_));
 sg13g2_a21oi_1 _20100_ (.A1(_03867_),
    .A2(_03868_),
    .Y(_03869_),
    .B1(net853));
 sg13g2_a21o_1 _20101_ (.A2(_03834_),
    .A1(\top_ihp.wb_dati_ram[2] ),
    .B1(_03869_),
    .X(_02470_));
 sg13g2_nand2_1 _20102_ (.Y(_03870_),
    .A(\top_ihp.wb_dati_ram[2] ),
    .B(net858));
 sg13g2_nand3_1 _20103_ (.B(net824),
    .C(net818),
    .A(_03748_),
    .Y(_03871_));
 sg13g2_a21oi_1 _20104_ (.A1(_03870_),
    .A2(_03871_),
    .Y(_03872_),
    .B1(net853));
 sg13g2_a21o_1 _20105_ (.A2(net835),
    .A1(\top_ihp.wb_dati_ram[3] ),
    .B1(_03872_),
    .X(_02471_));
 sg13g2_and2_1 _20106_ (.A(_03750_),
    .B(net817),
    .X(_03873_));
 sg13g2_a221oi_1 _20107_ (.B2(net802),
    .C1(net857),
    .B1(_03873_),
    .A1(\top_ihp.wb_dati_ram[3] ),
    .Y(_03874_),
    .A2(net852));
 sg13g2_a21oi_1 _20108_ (.A1(_09820_),
    .A2(net834),
    .Y(_02472_),
    .B1(_03874_));
 sg13g2_and2_1 _20109_ (.A(_03752_),
    .B(net817),
    .X(_03875_));
 sg13g2_a221oi_1 _20110_ (.B2(net802),
    .C1(net857),
    .B1(_03875_),
    .A1(\top_ihp.wb_dati_ram[4] ),
    .Y(_03876_),
    .A2(net852));
 sg13g2_a21oi_1 _20111_ (.A1(_09846_),
    .A2(net834),
    .Y(_02473_),
    .B1(_03876_));
 sg13g2_nand2_1 _20112_ (.Y(_03877_),
    .A(\top_ihp.wb_dati_ram[25] ),
    .B(net858));
 sg13g2_nand3_1 _20113_ (.B(net824),
    .C(net818),
    .A(\top_ihp.oisc.wb_dat_o[26] ),
    .Y(_03878_));
 sg13g2_a21oi_1 _20114_ (.A1(_03877_),
    .A2(_03878_),
    .Y(_03879_),
    .B1(net853));
 sg13g2_a21o_1 _20115_ (.A2(net835),
    .A1(\top_ihp.wb_dati_ram[26] ),
    .B1(_03879_),
    .X(_02474_));
 sg13g2_and2_1 _20116_ (.A(_03754_),
    .B(net817),
    .X(_03880_));
 sg13g2_a221oi_1 _20117_ (.B2(net802),
    .C1(net857),
    .B1(_03880_),
    .A1(\top_ihp.wb_dati_ram[5] ),
    .Y(_03881_),
    .A2(net852));
 sg13g2_a21oi_1 _20118_ (.A1(_09879_),
    .A2(net834),
    .Y(_02475_),
    .B1(_03881_));
 sg13g2_and2_1 _20119_ (.A(_03756_),
    .B(net837),
    .X(_03882_));
 sg13g2_a221oi_1 _20120_ (.B2(net820),
    .C1(net857),
    .B1(_03882_),
    .A1(\top_ihp.wb_dati_ram[6] ),
    .Y(_03883_),
    .A2(net852));
 sg13g2_a21oi_1 _20121_ (.A1(_09220_),
    .A2(net834),
    .Y(_02476_),
    .B1(_03883_));
 sg13g2_buf_1 _20122_ (.A(net866),
    .X(_03884_));
 sg13g2_buf_1 _20123_ (.A(net866),
    .X(_03885_));
 sg13g2_nor2_1 _20124_ (.A(_08173_),
    .B(_03885_),
    .Y(_03886_));
 sg13g2_a21oi_1 _20125_ (.A1(\top_ihp.wb_dati_ram[7] ),
    .A2(net851),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_nand2_1 _20126_ (.Y(_03888_),
    .A(\top_ihp.wb_emem.cmd[32] ),
    .B(net833));
 sg13g2_o21ai_1 _20127_ (.B1(_03888_),
    .Y(_02477_),
    .A1(net838),
    .A2(_03887_));
 sg13g2_nor2_1 _20128_ (.A(_08178_),
    .B(_03885_),
    .Y(_03889_));
 sg13g2_a21oi_1 _20129_ (.A1(\top_ihp.wb_emem.cmd[32] ),
    .A2(net851),
    .Y(_03890_),
    .B1(_03889_));
 sg13g2_nand2_1 _20130_ (.Y(_03891_),
    .A(\top_ihp.wb_emem.cmd[33] ),
    .B(net833));
 sg13g2_o21ai_1 _20131_ (.B1(_03891_),
    .Y(_02478_),
    .A1(net838),
    .A2(_03890_));
 sg13g2_buf_1 _20132_ (.A(net807),
    .X(_03892_));
 sg13g2_a21o_1 _20133_ (.A2(_09740_),
    .A1(net770),
    .B1(net982),
    .X(_03893_));
 sg13g2_nor2_1 _20134_ (.A(net1040),
    .B(_09740_),
    .Y(_03894_));
 sg13g2_a22oi_1 _20135_ (.Y(_03895_),
    .B1(_03894_),
    .B2(net777),
    .A2(_03893_),
    .A1(net1040));
 sg13g2_nor2_1 _20136_ (.A(net850),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_a21oi_1 _20137_ (.A1(\top_ihp.wb_emem.cmd[33] ),
    .A2(net851),
    .Y(_03897_),
    .B1(_03896_));
 sg13g2_nand2_1 _20138_ (.Y(_03898_),
    .A(\top_ihp.wb_emem.cmd[34] ),
    .B(net833));
 sg13g2_o21ai_1 _20139_ (.B1(_03898_),
    .Y(_02479_),
    .A1(net838),
    .A2(_03897_));
 sg13g2_a21o_1 _20140_ (.A2(_09794_),
    .A1(_03892_),
    .B1(net982),
    .X(_03899_));
 sg13g2_buf_1 _20141_ (.A(_07708_),
    .X(_03900_));
 sg13g2_nor3_1 _20142_ (.A(net1037),
    .B(_03900_),
    .C(_09794_),
    .Y(_03901_));
 sg13g2_a21oi_1 _20143_ (.A1(net1037),
    .A2(_03899_),
    .Y(_03902_),
    .B1(_03901_));
 sg13g2_nor2_1 _20144_ (.A(_03805_),
    .B(_03902_),
    .Y(_03903_));
 sg13g2_a21oi_1 _20145_ (.A1(\top_ihp.wb_emem.cmd[34] ),
    .A2(net851),
    .Y(_03904_),
    .B1(_03903_));
 sg13g2_nand2_1 _20146_ (.Y(_03905_),
    .A(\top_ihp.wb_emem.cmd[35] ),
    .B(net833));
 sg13g2_o21ai_1 _20147_ (.B1(_03905_),
    .Y(_02480_),
    .A1(net838),
    .A2(_03904_));
 sg13g2_nand2_1 _20148_ (.Y(_03906_),
    .A(net770),
    .B(_09834_));
 sg13g2_o21ai_1 _20149_ (.B1(net940),
    .Y(_03907_),
    .A1(_07708_),
    .A2(_09834_));
 sg13g2_nand2_1 _20150_ (.Y(_03908_),
    .A(net1039),
    .B(_03907_));
 sg13g2_o21ai_1 _20151_ (.B1(_03908_),
    .Y(_03909_),
    .A1(net1039),
    .A2(_03906_));
 sg13g2_and2_1 _20152_ (.A(_03816_),
    .B(_03909_),
    .X(_03910_));
 sg13g2_a21oi_1 _20153_ (.A1(\top_ihp.wb_emem.cmd[35] ),
    .A2(net851),
    .Y(_03911_),
    .B1(_03910_));
 sg13g2_nand2_1 _20154_ (.Y(_03912_),
    .A(\top_ihp.wb_emem.cmd[36] ),
    .B(net833));
 sg13g2_o21ai_1 _20155_ (.B1(_03912_),
    .Y(_02481_),
    .A1(net838),
    .A2(_03911_));
 sg13g2_nand2_1 _20156_ (.Y(_03913_),
    .A(net770),
    .B(_09862_));
 sg13g2_o21ai_1 _20157_ (.B1(net940),
    .Y(_03914_),
    .A1(_07708_),
    .A2(_09862_));
 sg13g2_nand2_1 _20158_ (.Y(_03915_),
    .A(net1038),
    .B(_03914_));
 sg13g2_o21ai_1 _20159_ (.B1(_03915_),
    .Y(_03916_),
    .A1(net1038),
    .A2(_03913_));
 sg13g2_buf_1 _20160_ (.A(_08181_),
    .X(_03917_));
 sg13g2_inv_1 _20161_ (.Y(_03918_),
    .A(_03917_));
 sg13g2_nand2b_1 _20162_ (.Y(_03919_),
    .B(net907),
    .A_N(_03916_));
 sg13g2_o21ai_1 _20163_ (.B1(_03919_),
    .Y(_03920_),
    .A1(\top_ihp.wb_emem.cmd[36] ),
    .A2(net819));
 sg13g2_buf_1 _20164_ (.A(_03801_),
    .X(_03921_));
 sg13g2_nand2_1 _20165_ (.Y(_03922_),
    .A(\top_ihp.wb_emem.cmd[37] ),
    .B(net832));
 sg13g2_o21ai_1 _20166_ (.B1(_03922_),
    .Y(_02482_),
    .A1(net838),
    .A2(_03920_));
 sg13g2_inv_1 _20167_ (.Y(_03923_),
    .A(\top_ihp.wb_emem.cmd[37] ));
 sg13g2_a21o_1 _20168_ (.A2(_09874_),
    .A1(net770),
    .B1(net912),
    .X(_03924_));
 sg13g2_buf_1 _20169_ (.A(net769),
    .X(_03925_));
 sg13g2_nor3_1 _20170_ (.A(net1031),
    .B(net734),
    .C(_09874_),
    .Y(_03926_));
 sg13g2_a21oi_1 _20171_ (.A1(net1031),
    .A2(_03924_),
    .Y(_03927_),
    .B1(_03926_));
 sg13g2_a221oi_1 _20172_ (.B2(net907),
    .C1(_03801_),
    .B1(_03927_),
    .A1(_03923_),
    .Y(_03928_),
    .A2(net850));
 sg13g2_a21o_1 _20173_ (.A2(net835),
    .A1(\top_ihp.wb_emem.cmd[38] ),
    .B1(_03928_),
    .X(_02483_));
 sg13g2_buf_1 _20174_ (.A(net856),
    .X(_03929_));
 sg13g2_a21o_1 _20175_ (.A2(_09900_),
    .A1(net770),
    .B1(net982),
    .X(_03930_));
 sg13g2_nor3_1 _20176_ (.A(net1033),
    .B(net769),
    .C(_09900_),
    .Y(_03931_));
 sg13g2_a21oi_1 _20177_ (.A1(net1033),
    .A2(_03930_),
    .Y(_03932_),
    .B1(_03931_));
 sg13g2_buf_1 _20178_ (.A(net947),
    .X(_03933_));
 sg13g2_a22oi_1 _20179_ (.Y(_03934_),
    .B1(\top_ihp.wb_emem.cmd[39] ),
    .B2(net832),
    .A2(\top_ihp.wb_emem.cmd[38] ),
    .A1(net906));
 sg13g2_o21ai_1 _20180_ (.B1(_03934_),
    .Y(_02484_),
    .A1(net831),
    .A2(_03932_));
 sg13g2_nand2_1 _20181_ (.Y(_03935_),
    .A(\top_ihp.wb_dati_ram[26] ),
    .B(net866));
 sg13g2_nand3_1 _20182_ (.B(_07657_),
    .C(net818),
    .A(\top_ihp.oisc.wb_dat_o[27] ),
    .Y(_03936_));
 sg13g2_a21oi_1 _20183_ (.A1(_03935_),
    .A2(_03936_),
    .Y(_03937_),
    .B1(_03827_));
 sg13g2_a21o_1 _20184_ (.A2(net835),
    .A1(\top_ihp.wb_dati_ram[27] ),
    .B1(_03937_),
    .X(_02485_));
 sg13g2_a21o_1 _20185_ (.A2(_09917_),
    .A1(net777),
    .B1(net912),
    .X(_03938_));
 sg13g2_nor3_1 _20186_ (.A(net1015),
    .B(net734),
    .C(_09917_),
    .Y(_03939_));
 sg13g2_a21oi_1 _20187_ (.A1(net1015),
    .A2(_03938_),
    .Y(_03940_),
    .B1(_03939_));
 sg13g2_a22oi_1 _20188_ (.Y(_03941_),
    .B1(\top_ihp.wb_emem.cmd[40] ),
    .B2(net832),
    .A2(\top_ihp.wb_emem.cmd[39] ),
    .A1(net906));
 sg13g2_o21ai_1 _20189_ (.B1(_03941_),
    .Y(_02486_),
    .A1(net831),
    .A2(_03940_));
 sg13g2_xnor2_1 _20190_ (.Y(_03942_),
    .A(_07548_),
    .B(_09937_));
 sg13g2_a21o_1 _20191_ (.A2(_03942_),
    .A1(net770),
    .B1(net982),
    .X(_03943_));
 sg13g2_nor3_1 _20192_ (.A(net1032),
    .B(net769),
    .C(_03942_),
    .Y(_03944_));
 sg13g2_a21oi_1 _20193_ (.A1(net1032),
    .A2(_03943_),
    .Y(_03945_),
    .B1(_03944_));
 sg13g2_buf_1 _20194_ (.A(net947),
    .X(_03946_));
 sg13g2_a22oi_1 _20195_ (.Y(_03947_),
    .B1(\top_ihp.wb_emem.cmd[41] ),
    .B2(_03921_),
    .A2(\top_ihp.wb_emem.cmd[40] ),
    .A1(net905));
 sg13g2_o21ai_1 _20196_ (.B1(_03947_),
    .Y(_02487_),
    .A1(net831),
    .A2(_03945_));
 sg13g2_xnor2_1 _20197_ (.Y(_03948_),
    .A(_07535_),
    .B(_09263_));
 sg13g2_nor2_1 _20198_ (.A(_07534_),
    .B(net734),
    .Y(_03949_));
 sg13g2_o21ai_1 _20199_ (.B1(net940),
    .Y(_03950_),
    .A1(net769),
    .A2(_03948_));
 sg13g2_a22oi_1 _20200_ (.Y(_03951_),
    .B1(_03950_),
    .B2(_07534_),
    .A2(_03949_),
    .A1(_03948_));
 sg13g2_a22oi_1 _20201_ (.Y(_03952_),
    .B1(\top_ihp.wb_emem.cmd[42] ),
    .B2(net832),
    .A2(\top_ihp.wb_emem.cmd[41] ),
    .A1(net905));
 sg13g2_o21ai_1 _20202_ (.B1(_03952_),
    .Y(_02488_),
    .A1(net831),
    .A2(_03951_));
 sg13g2_a22oi_1 _20203_ (.Y(_03953_),
    .B1(net777),
    .B2(_09292_),
    .A2(_07531_),
    .A1(net912));
 sg13g2_a22oi_1 _20204_ (.Y(_03954_),
    .B1(\top_ihp.wb_emem.cmd[43] ),
    .B2(_03921_),
    .A2(\top_ihp.wb_emem.cmd[42] ),
    .A1(net905));
 sg13g2_o21ai_1 _20205_ (.B1(_03954_),
    .Y(_02489_),
    .A1(net831),
    .A2(_03953_));
 sg13g2_nand2_1 _20206_ (.Y(_03955_),
    .A(net912),
    .B(_07528_));
 sg13g2_o21ai_1 _20207_ (.B1(_03955_),
    .Y(_03956_),
    .A1(net734),
    .A2(_09325_));
 sg13g2_nand2_1 _20208_ (.Y(_03957_),
    .A(_03810_),
    .B(_03956_));
 sg13g2_a22oi_1 _20209_ (.Y(_03958_),
    .B1(\top_ihp.wb_emem.cmd[44] ),
    .B2(net833),
    .A2(\top_ihp.wb_emem.cmd[43] ),
    .A1(net906));
 sg13g2_nand2_1 _20210_ (.Y(_02490_),
    .A(_03957_),
    .B(_03958_));
 sg13g2_xor2_1 _20211_ (.B(_07884_),
    .A(_07526_),
    .X(_03959_));
 sg13g2_nor2_1 _20212_ (.A(net1034),
    .B(net769),
    .Y(_03960_));
 sg13g2_o21ai_1 _20213_ (.B1(net940),
    .Y(_03961_),
    .A1(net769),
    .A2(_03959_));
 sg13g2_a22oi_1 _20214_ (.Y(_03962_),
    .B1(_03961_),
    .B2(net1034),
    .A2(_03960_),
    .A1(_03959_));
 sg13g2_a22oi_1 _20215_ (.Y(_03963_),
    .B1(\top_ihp.wb_emem.cmd[45] ),
    .B2(net832),
    .A2(\top_ihp.wb_emem.cmd[44] ),
    .A1(net905));
 sg13g2_o21ai_1 _20216_ (.B1(_03963_),
    .Y(_02491_),
    .A1(net831),
    .A2(_03962_));
 sg13g2_xnor2_1 _20217_ (.Y(_03964_),
    .A(_07522_),
    .B(_09396_));
 sg13g2_a21o_1 _20218_ (.A2(_03964_),
    .A1(net770),
    .B1(net982),
    .X(_03965_));
 sg13g2_nor3_1 _20219_ (.A(_07521_),
    .B(net769),
    .C(_03964_),
    .Y(_03966_));
 sg13g2_a21oi_1 _20220_ (.A1(_07521_),
    .A2(_03965_),
    .Y(_03967_),
    .B1(_03966_));
 sg13g2_a22oi_1 _20221_ (.Y(_03968_),
    .B1(\top_ihp.wb_emem.cmd[46] ),
    .B2(_03818_),
    .A2(\top_ihp.wb_emem.cmd[45] ),
    .A1(net905));
 sg13g2_o21ai_1 _20222_ (.B1(_03968_),
    .Y(_02492_),
    .A1(net831),
    .A2(_03967_));
 sg13g2_o21ai_1 _20223_ (.B1(net940),
    .Y(_03969_),
    .A1(net734),
    .A2(_09411_));
 sg13g2_nor2_1 _20224_ (.A(net1036),
    .B(net734),
    .Y(_03970_));
 sg13g2_a22oi_1 _20225_ (.Y(_03971_),
    .B1(_03970_),
    .B2(_09411_),
    .A2(_03969_),
    .A1(net1036));
 sg13g2_a22oi_1 _20226_ (.Y(_03972_),
    .B1(\top_ihp.wb_emem.cmd[47] ),
    .B2(net855),
    .A2(\top_ihp.wb_emem.cmd[46] ),
    .A1(net905));
 sg13g2_o21ai_1 _20227_ (.B1(_03972_),
    .Y(_02493_),
    .A1(net831),
    .A2(_03971_));
 sg13g2_xnor2_1 _20228_ (.Y(_03973_),
    .A(_07508_),
    .B(_09423_));
 sg13g2_a21oi_1 _20229_ (.A1(net777),
    .A2(_03973_),
    .Y(_03974_),
    .B1(net912));
 sg13g2_or3_1 _20230_ (.A(_07507_),
    .B(net734),
    .C(_03973_),
    .X(_03975_));
 sg13g2_o21ai_1 _20231_ (.B1(_03975_),
    .Y(_03976_),
    .A1(_07905_),
    .A2(_03974_));
 sg13g2_inv_1 _20232_ (.Y(_03977_),
    .A(\top_ihp.wb_emem.cmd[47] ));
 sg13g2_a22oi_1 _20233_ (.Y(_03978_),
    .B1(_00214_),
    .B2(net855),
    .A2(_03977_),
    .A1(_03946_));
 sg13g2_o21ai_1 _20234_ (.B1(_03978_),
    .Y(_02494_),
    .A1(_03929_),
    .A2(_03976_));
 sg13g2_a22oi_1 _20235_ (.Y(_03979_),
    .B1(net777),
    .B2(_09453_),
    .A2(net1035),
    .A1(net912));
 sg13g2_a22oi_1 _20236_ (.Y(_03980_),
    .B1(\top_ihp.wb_emem.cmd[49] ),
    .B2(net855),
    .A2(\top_ihp.wb_emem.cmd[48] ),
    .A1(net905));
 sg13g2_o21ai_1 _20237_ (.B1(_03980_),
    .Y(_02495_),
    .A1(_03929_),
    .A2(_03979_));
 sg13g2_and2_1 _20238_ (.A(\top_ihp.oisc.wb_dat_o[28] ),
    .B(net837),
    .X(_03981_));
 sg13g2_a221oi_1 _20239_ (.B2(net820),
    .C1(net857),
    .B1(_03981_),
    .A1(\top_ihp.wb_dati_ram[27] ),
    .Y(_03982_),
    .A2(_03852_));
 sg13g2_a21oi_1 _20240_ (.A1(_09336_),
    .A2(net834),
    .Y(_02496_),
    .B1(_03982_));
 sg13g2_xnor2_1 _20241_ (.Y(_03983_),
    .A(_07890_),
    .B(_09466_));
 sg13g2_a21o_1 _20242_ (.A2(_03983_),
    .A1(_03892_),
    .B1(net982),
    .X(_03984_));
 sg13g2_nor3_1 _20243_ (.A(net1043),
    .B(_03900_),
    .C(_03983_),
    .Y(_03985_));
 sg13g2_a21oi_1 _20244_ (.A1(net1043),
    .A2(_03984_),
    .Y(_03986_),
    .B1(_03985_));
 sg13g2_a22oi_1 _20245_ (.Y(_03987_),
    .B1(\top_ihp.wb_emem.cmd[50] ),
    .B2(net855),
    .A2(\top_ihp.wb_emem.cmd[49] ),
    .A1(net905));
 sg13g2_o21ai_1 _20246_ (.B1(_03987_),
    .Y(_02497_),
    .A1(net851),
    .A2(_03986_));
 sg13g2_a22oi_1 _20247_ (.Y(_03988_),
    .B1(_07441_),
    .B2(_09494_),
    .A2(net1042),
    .A1(net912));
 sg13g2_nor2_1 _20248_ (.A(_03918_),
    .B(\top_ihp.wb_emem.cmd[50] ),
    .Y(_03989_));
 sg13g2_a221oi_1 _20249_ (.B2(_03810_),
    .C1(_03989_),
    .B1(_03988_),
    .A1(_00215_),
    .Y(_03990_),
    .A2(_03801_));
 sg13g2_inv_1 _20250_ (.Y(_02498_),
    .A(_03990_));
 sg13g2_o21ai_1 _20251_ (.B1(net777),
    .Y(_03991_),
    .A1(_09560_),
    .A2(_09561_));
 sg13g2_o21ai_1 _20252_ (.B1(_03991_),
    .Y(_03992_),
    .A1(_08169_),
    .A2(_07451_));
 sg13g2_inv_1 _20253_ (.Y(_03993_),
    .A(\top_ihp.wb_emem.cmd[51] ));
 sg13g2_a22oi_1 _20254_ (.Y(_03994_),
    .B1(_00216_),
    .B2(net855),
    .A2(_03993_),
    .A1(_03946_));
 sg13g2_o21ai_1 _20255_ (.B1(_03994_),
    .Y(_02499_),
    .A1(net851),
    .A2(_03992_));
 sg13g2_o21ai_1 _20256_ (.B1(net940),
    .Y(_03995_),
    .A1(_03925_),
    .A2(_09592_));
 sg13g2_nand2_1 _20257_ (.Y(_03996_),
    .A(_07441_),
    .B(_09592_));
 sg13g2_nor2_1 _20258_ (.A(_07461_),
    .B(_03996_),
    .Y(_03997_));
 sg13g2_a21oi_1 _20259_ (.A1(_07461_),
    .A2(_03995_),
    .Y(_03998_),
    .B1(_03997_));
 sg13g2_a22oi_1 _20260_ (.Y(_03999_),
    .B1(\top_ihp.wb_emem.cmd[53] ),
    .B2(net855),
    .A2(\top_ihp.wb_emem.cmd[52] ),
    .A1(net947));
 sg13g2_o21ai_1 _20261_ (.B1(_03999_),
    .Y(_02500_),
    .A1(net851),
    .A2(_03998_));
 sg13g2_nand3b_1 _20262_ (.B(_07470_),
    .C(_09609_),
    .Y(_04000_),
    .A_N(net1044));
 sg13g2_o21ai_1 _20263_ (.B1(net1044),
    .Y(_04001_),
    .A1(_07602_),
    .A2(_09611_));
 sg13g2_a21oi_1 _20264_ (.A1(_04000_),
    .A2(_04001_),
    .Y(_04002_),
    .B1(net734));
 sg13g2_nand3_1 _20265_ (.B(_04000_),
    .C(_04001_),
    .A(net770),
    .Y(_04003_));
 sg13g2_a21oi_1 _20266_ (.A1(_08169_),
    .A2(_04003_),
    .Y(_04004_),
    .B1(_07801_));
 sg13g2_a21oi_1 _20267_ (.A1(_07801_),
    .A2(_04002_),
    .Y(_04005_),
    .B1(_04004_));
 sg13g2_a22oi_1 _20268_ (.Y(_04006_),
    .B1(\top_ihp.wb_emem.cmd[54] ),
    .B2(net855),
    .A2(\top_ihp.wb_emem.cmd[53] ),
    .A1(_03917_));
 sg13g2_o21ai_1 _20269_ (.B1(_04006_),
    .Y(_02501_),
    .A1(_03884_),
    .A2(_04005_));
 sg13g2_nand2_1 _20270_ (.Y(_04007_),
    .A(_03683_),
    .B(_07442_));
 sg13g2_o21ai_1 _20271_ (.B1(_04007_),
    .Y(_04008_),
    .A1(_03925_),
    .A2(_09639_));
 sg13g2_inv_1 _20272_ (.Y(_04009_),
    .A(\top_ihp.wb_emem.cmd[54] ));
 sg13g2_a22oi_1 _20273_ (.Y(_04010_),
    .B1(_00217_),
    .B2(net855),
    .A2(_04009_),
    .A1(net947));
 sg13g2_o21ai_1 _20274_ (.B1(_04010_),
    .Y(_02502_),
    .A1(_03884_),
    .A2(_04008_));
 sg13g2_inv_1 _20275_ (.Y(_04011_),
    .A(\top_ihp.wb_emem.cmd[56] ));
 sg13g2_buf_1 _20276_ (.A(_08182_),
    .X(_04012_));
 sg13g2_o21ai_1 _20277_ (.B1(net907),
    .Y(_04013_),
    .A1(net946),
    .A2(net869));
 sg13g2_nand2_1 _20278_ (.Y(_04014_),
    .A(\top_ihp.wb_emem.cmd[55] ),
    .B(net866));
 sg13g2_o21ai_1 _20279_ (.B1(_04014_),
    .Y(_04015_),
    .A1(net820),
    .A2(net850));
 sg13g2_nand2_1 _20280_ (.Y(_04016_),
    .A(_04013_),
    .B(_04015_));
 sg13g2_o21ai_1 _20281_ (.B1(_04016_),
    .Y(_02503_),
    .A1(_04011_),
    .A2(_04013_));
 sg13g2_a22oi_1 _20282_ (.Y(_04017_),
    .B1(_00218_),
    .B2(net835),
    .A2(_04011_),
    .A1(net906));
 sg13g2_inv_1 _20283_ (.Y(_02504_),
    .A(_04017_));
 sg13g2_o21ai_1 _20284_ (.B1(net850),
    .Y(_04018_),
    .A1(net907),
    .A2(\top_ihp.wb_emem.cmd[57] ));
 sg13g2_a21oi_1 _20285_ (.A1(_00219_),
    .A2(net832),
    .Y(_04019_),
    .B1(_04018_));
 sg13g2_inv_1 _20286_ (.Y(_02505_),
    .A(_04019_));
 sg13g2_a22oi_1 _20287_ (.Y(_04020_),
    .B1(\top_ihp.wb_emem.cmd[59] ),
    .B2(_03862_),
    .A2(\top_ihp.wb_emem.cmd[58] ),
    .A1(net906));
 sg13g2_inv_1 _20288_ (.Y(_02506_),
    .A(_04020_));
 sg13g2_nand2_1 _20289_ (.Y(_04021_),
    .A(\top_ihp.wb_dati_ram[28] ),
    .B(net866));
 sg13g2_nand3_1 _20290_ (.B(_07657_),
    .C(net818),
    .A(\top_ihp.oisc.wb_dat_o[29] ),
    .Y(_04022_));
 sg13g2_a21oi_1 _20291_ (.A1(_04021_),
    .A2(_04022_),
    .Y(_04023_),
    .B1(_03827_));
 sg13g2_a21o_1 _20292_ (.A2(net835),
    .A1(\top_ihp.wb_dati_ram[29] ),
    .B1(_04023_),
    .X(_02507_));
 sg13g2_a22oi_1 _20293_ (.Y(_04024_),
    .B1(\top_ihp.wb_emem.cmd[60] ),
    .B2(_03862_),
    .A2(\top_ihp.wb_emem.cmd[59] ),
    .A1(net906));
 sg13g2_inv_1 _20294_ (.Y(_02508_),
    .A(_04024_));
 sg13g2_o21ai_1 _20295_ (.B1(net850),
    .Y(_04025_),
    .A1(net907),
    .A2(\top_ihp.wb_emem.cmd[60] ));
 sg13g2_a21oi_1 _20296_ (.A1(_00220_),
    .A2(net832),
    .Y(_04026_),
    .B1(_04025_));
 sg13g2_inv_1 _20297_ (.Y(_02509_),
    .A(_04026_));
 sg13g2_o21ai_1 _20298_ (.B1(net850),
    .Y(_04027_),
    .A1(net907),
    .A2(\top_ihp.wb_emem.cmd[61] ));
 sg13g2_a21oi_1 _20299_ (.A1(_00221_),
    .A2(net832),
    .Y(_04028_),
    .B1(_04027_));
 sg13g2_inv_1 _20300_ (.Y(_02510_),
    .A(_04028_));
 sg13g2_a22oi_1 _20301_ (.Y(_04029_),
    .B1(\top_ihp.wb_emem.cmd[63] ),
    .B2(net833),
    .A2(\top_ihp.wb_emem.cmd[62] ),
    .A1(_03933_));
 sg13g2_inv_1 _20302_ (.Y(_02511_),
    .A(_04029_));
 sg13g2_and2_1 _20303_ (.A(\top_ihp.oisc.wb_dat_o[30] ),
    .B(net837),
    .X(_04030_));
 sg13g2_a221oi_1 _20304_ (.B2(_03807_),
    .C1(net857),
    .B1(_04030_),
    .A1(\top_ihp.wb_dati_ram[29] ),
    .Y(_04031_),
    .A2(_03852_));
 sg13g2_a21oi_1 _20305_ (.A1(_09386_),
    .A2(net834),
    .Y(_02512_),
    .B1(_04031_));
 sg13g2_and2_1 _20306_ (.A(\top_ihp.oisc.wb_dat_o[31] ),
    .B(_03809_),
    .X(_04032_));
 sg13g2_a221oi_1 _20307_ (.B2(net820),
    .C1(net857),
    .B1(_04032_),
    .A1(\top_ihp.wb_dati_ram[30] ),
    .Y(_04033_),
    .A2(net852));
 sg13g2_a21oi_1 _20308_ (.A1(_09231_),
    .A2(net834),
    .Y(_02513_),
    .B1(_04033_));
 sg13g2_and2_1 _20309_ (.A(\top_ihp.oisc.wb_dat_o[16] ),
    .B(net837),
    .X(_04034_));
 sg13g2_a221oi_1 _20310_ (.B2(net820),
    .C1(_03812_),
    .B1(_04034_),
    .A1(\top_ihp.wb_dati_ram[31] ),
    .Y(_04035_),
    .A2(net850));
 sg13g2_a21oi_1 _20311_ (.A1(_09129_),
    .A2(_03857_),
    .Y(_02514_),
    .B1(_04035_));
 sg13g2_and2_1 _20312_ (.A(\top_ihp.oisc.wb_dat_o[17] ),
    .B(_03809_),
    .X(_04036_));
 sg13g2_a221oi_1 _20313_ (.B2(_03807_),
    .C1(_03812_),
    .B1(_04036_),
    .A1(\top_ihp.wb_dati_ram[16] ),
    .Y(_04037_),
    .A2(net850));
 sg13g2_a21oi_1 _20314_ (.A1(_09445_),
    .A2(net834),
    .Y(_02515_),
    .B1(_04037_));
 sg13g2_xnor2_1 _20315_ (.Y(_04038_),
    .A(_03792_),
    .B(\top_ihp.wb_emem.nbits[6] ));
 sg13g2_buf_1 _20316_ (.A(\top_ihp.wb_emem.nbits[3] ),
    .X(_04039_));
 sg13g2_buf_2 _20317_ (.A(\top_ihp.wb_emem.nbits[4] ),
    .X(_04040_));
 sg13g2_buf_1 _20318_ (.A(\top_ihp.wb_emem.nbits[5] ),
    .X(_04041_));
 sg13g2_inv_1 _20319_ (.Y(_04042_),
    .A(_04041_));
 sg13g2_nor3_1 _20320_ (.A(_04039_),
    .B(_04040_),
    .C(_04042_),
    .Y(_04043_));
 sg13g2_a21oi_1 _20321_ (.A1(_04039_),
    .A2(_04040_),
    .Y(_04044_),
    .B1(_04043_));
 sg13g2_xor2_1 _20322_ (.B(_04040_),
    .A(_04039_),
    .X(_04045_));
 sg13g2_nor2_1 _20323_ (.A(_03783_),
    .B(_04045_),
    .Y(_04046_));
 sg13g2_a21oi_1 _20324_ (.A1(_03783_),
    .A2(_04044_),
    .Y(_04047_),
    .B1(_04046_));
 sg13g2_nor2b_1 _20325_ (.A(_04041_),
    .B_N(\top_ihp.wb_emem.nbits[6] ),
    .Y(_04048_));
 sg13g2_nor4_1 _20326_ (.A(_03787_),
    .B(_03792_),
    .C(_04039_),
    .D(_04040_),
    .Y(_04049_));
 sg13g2_a22oi_1 _20327_ (.Y(_04050_),
    .B1(_04048_),
    .B2(_04049_),
    .A2(_04047_),
    .A1(_04038_));
 sg13g2_xnor2_1 _20328_ (.Y(_04051_),
    .A(_03791_),
    .B(_04041_));
 sg13g2_inv_1 _20329_ (.Y(_04052_),
    .A(_04039_));
 sg13g2_nor2_1 _20330_ (.A(_03777_),
    .B(_04052_),
    .Y(_04053_));
 sg13g2_xor2_1 _20331_ (.B(_04051_),
    .A(_04040_),
    .X(_04054_));
 sg13g2_nor2_1 _20332_ (.A(_04039_),
    .B(_04054_),
    .Y(_04055_));
 sg13g2_a22oi_1 _20333_ (.Y(_04056_),
    .B1(_04055_),
    .B2(_03777_),
    .A2(_04053_),
    .A1(_04051_));
 sg13g2_nor4_1 _20334_ (.A(\top_ihp.wb_emem.bit_counter[7] ),
    .B(_03780_),
    .C(_04050_),
    .D(_04056_),
    .Y(_04057_));
 sg13g2_a21o_1 _20335_ (.A2(_03771_),
    .A1(_08180_),
    .B1(_04057_),
    .X(_02516_));
 sg13g2_buf_1 _20336_ (.A(\top_ihp.wb_emem.last_wait ),
    .X(_04058_));
 sg13g2_inv_1 _20337_ (.Y(_04059_),
    .A(_04058_));
 sg13g2_xor2_1 _20338_ (.B(net1013),
    .A(_08185_),
    .X(_04060_));
 sg13g2_and2_1 _20339_ (.A(_08184_),
    .B(_04060_),
    .X(_04061_));
 sg13g2_buf_2 _20340_ (.A(_04061_),
    .X(_04062_));
 sg13g2_inv_1 _20341_ (.Y(_04063_),
    .A(\top_ihp.wb_emem.wait_counter[3] ));
 sg13g2_buf_1 _20342_ (.A(\top_ihp.wb_emem.wait_counter[1] ),
    .X(_04064_));
 sg13g2_buf_2 _20343_ (.A(\top_ihp.wb_emem.wait_counter[0] ),
    .X(_04065_));
 sg13g2_nand3_1 _20344_ (.B(_04065_),
    .C(\top_ihp.wb_emem.wait_counter[2] ),
    .A(_04064_),
    .Y(_04066_));
 sg13g2_nor2_1 _20345_ (.A(_04063_),
    .B(_04066_),
    .Y(_04067_));
 sg13g2_buf_1 _20346_ (.A(\top_ihp.wb_emem.wait_counter[5] ),
    .X(_04068_));
 sg13g2_buf_1 _20347_ (.A(\top_ihp.wb_emem.wait_counter[4] ),
    .X(_04069_));
 sg13g2_buf_1 _20348_ (.A(\top_ihp.wb_emem.wait_counter[6] ),
    .X(_04070_));
 sg13g2_nor4_1 _20349_ (.A(_04068_),
    .B(_04069_),
    .C(\top_ihp.wb_emem.wait_counter[7] ),
    .D(_04070_),
    .Y(_04071_));
 sg13g2_nand3_1 _20350_ (.B(_04071_),
    .C(_04062_),
    .A(_04067_),
    .Y(_04072_));
 sg13g2_o21ai_1 _20351_ (.B1(_04072_),
    .Y(_02517_),
    .A1(_04059_),
    .A2(_04062_));
 sg13g2_buf_1 _20352_ (.A(_08185_),
    .X(_04073_));
 sg13g2_inv_1 _20353_ (.Y(_04074_),
    .A(_08186_));
 sg13g2_nand2_1 _20354_ (.Y(_04075_),
    .A(net945),
    .B(_04074_));
 sg13g2_nand3_1 _20355_ (.B(_08184_),
    .C(_04075_),
    .A(_08939_),
    .Y(_04076_));
 sg13g2_buf_1 _20356_ (.A(_04076_),
    .X(_04077_));
 sg13g2_nand2_1 _20357_ (.Y(_04078_),
    .A(_08939_),
    .B(net837));
 sg13g2_inv_1 _20358_ (.Y(_04079_),
    .A(_04078_));
 sg13g2_nand3_1 _20359_ (.B(_07658_),
    .C(_09158_),
    .A(_07824_),
    .Y(_04080_));
 sg13g2_a22oi_1 _20360_ (.Y(_02518_),
    .B1(_04079_),
    .B2(_04080_),
    .A2(_04077_),
    .A1(_04052_));
 sg13g2_nand2_1 _20361_ (.Y(_04081_),
    .A(_04040_),
    .B(_04077_));
 sg13g2_and3_1 _20362_ (.X(_04082_),
    .A(_09240_),
    .B(_07826_),
    .C(_07830_));
 sg13g2_buf_1 _20363_ (.A(_04082_),
    .X(_04083_));
 sg13g2_buf_1 _20364_ (.A(net816),
    .X(_04084_));
 sg13g2_nand3_1 _20365_ (.B(_04079_),
    .C(_04084_),
    .A(net806),
    .Y(_04085_));
 sg13g2_nand2_1 _20366_ (.Y(_02519_),
    .A(_04081_),
    .B(_04085_));
 sg13g2_nand3_1 _20367_ (.B(_07830_),
    .C(_04079_),
    .A(net806),
    .Y(_04086_));
 sg13g2_nand2_1 _20368_ (.Y(_04087_),
    .A(_04041_),
    .B(_04077_));
 sg13g2_nand2_1 _20369_ (.Y(_02520_),
    .A(_04086_),
    .B(_04087_));
 sg13g2_a21oi_1 _20370_ (.A1(net806),
    .A2(_07830_),
    .Y(_04088_),
    .B1(_04078_));
 sg13g2_a21o_1 _20371_ (.A2(_04077_),
    .A1(\top_ihp.wb_emem.nbits[6] ),
    .B1(_04088_),
    .X(_02521_));
 sg13g2_or2_1 _20372_ (.X(_04089_),
    .B(_08982_),
    .A(net769));
 sg13g2_a21oi_1 _20373_ (.A1(net912),
    .A2(_08946_),
    .Y(_04090_),
    .B1(_03804_));
 sg13g2_o21ai_1 _20374_ (.B1(_04090_),
    .Y(_04091_),
    .A1(_09772_),
    .A2(_04089_));
 sg13g2_nor2_1 _20375_ (.A(net1013),
    .B(net947),
    .Y(_04092_));
 sg13g2_a22oi_1 _20376_ (.Y(_04093_),
    .B1(_04058_),
    .B2(_04092_),
    .A2(net946),
    .A1(net1013));
 sg13g2_nand2b_1 _20377_ (.Y(_04094_),
    .B(net945),
    .A_N(_04093_));
 sg13g2_nor2_1 _20378_ (.A(net945),
    .B(net946),
    .Y(_04095_));
 sg13g2_o21ai_1 _20379_ (.B1(net1013),
    .Y(_04096_),
    .A1(net947),
    .A2(_04095_));
 sg13g2_nand2_1 _20380_ (.Y(_04097_),
    .A(net946),
    .B(_04092_));
 sg13g2_nand4_1 _20381_ (.B(_04094_),
    .C(_04096_),
    .A(_04091_),
    .Y(_02522_),
    .D(_04097_));
 sg13g2_inv_1 _20382_ (.Y(_04098_),
    .A(net945));
 sg13g2_nor3_1 _20383_ (.A(net1013),
    .B(_08182_),
    .C(_04058_),
    .Y(_04099_));
 sg13g2_a21oi_1 _20384_ (.A1(net1013),
    .A2(_04012_),
    .Y(_04100_),
    .B1(_04099_));
 sg13g2_nand2_1 _20385_ (.Y(_04101_),
    .A(net946),
    .B(_08180_));
 sg13g2_nor2_1 _20386_ (.A(_04074_),
    .B(_04058_),
    .Y(_04102_));
 sg13g2_a22oi_1 _20387_ (.Y(_04103_),
    .B1(_04102_),
    .B2(_04095_),
    .A2(_04101_),
    .A1(_08181_));
 sg13g2_o21ai_1 _20388_ (.B1(_04103_),
    .Y(_04104_),
    .A1(_04098_),
    .A2(_04100_));
 sg13g2_nand2b_1 _20389_ (.Y(_04105_),
    .B(_04091_),
    .A_N(_04104_));
 sg13g2_nor3_1 _20390_ (.A(net945),
    .B(_04074_),
    .C(_03798_),
    .Y(_04106_));
 sg13g2_a21oi_1 _20391_ (.A1(net945),
    .A2(_03798_),
    .Y(_04107_),
    .B1(_04106_));
 sg13g2_nand3_1 _20392_ (.B(_04074_),
    .C(net946),
    .A(_04073_),
    .Y(_04108_));
 sg13g2_o21ai_1 _20393_ (.B1(_04108_),
    .Y(_04109_),
    .A1(net947),
    .A2(_04107_));
 sg13g2_a21o_1 _20394_ (.A2(_04105_),
    .A1(_04073_),
    .B1(_04109_),
    .X(_02523_));
 sg13g2_nor2_1 _20395_ (.A(_08188_),
    .B(_04095_),
    .Y(_04110_));
 sg13g2_o21ai_1 _20396_ (.B1(net906),
    .Y(_04111_),
    .A1(_03798_),
    .A2(_04104_));
 sg13g2_o21ai_1 _20397_ (.B1(_04111_),
    .Y(_02524_),
    .A1(_04105_),
    .A2(_04110_));
 sg13g2_nand2_1 _20398_ (.Y(_04112_),
    .A(net907),
    .B(_04110_));
 sg13g2_mux2_1 _20399_ (.A0(_04112_),
    .A1(_04012_),
    .S(_04105_),
    .X(_02525_));
 sg13g2_inv_1 _20400_ (.Y(_04113_),
    .A(_04065_));
 sg13g2_o21ai_1 _20401_ (.B1(_04065_),
    .Y(_04114_),
    .A1(net945),
    .A2(_03798_));
 sg13g2_nor3_1 _20402_ (.A(net947),
    .B(net946),
    .C(_00139_),
    .Y(_04115_));
 sg13g2_mux2_1 _20403_ (.A0(_04113_),
    .A1(_04115_),
    .S(_04060_),
    .X(_04116_));
 sg13g2_a221oi_1 _20404_ (.B2(net906),
    .C1(_04116_),
    .B1(_04114_),
    .A1(net946),
    .Y(_02526_),
    .A2(_04113_));
 sg13g2_nand2_1 _20405_ (.Y(_04117_),
    .A(_04065_),
    .B(_04062_));
 sg13g2_o21ai_1 _20406_ (.B1(_03763_),
    .Y(_04118_),
    .A1(_04074_),
    .A2(net868));
 sg13g2_nor2_1 _20407_ (.A(net868),
    .B(_04075_),
    .Y(_04119_));
 sg13g2_a21oi_1 _20408_ (.A1(_04098_),
    .A2(_04118_),
    .Y(_04120_),
    .B1(_04119_));
 sg13g2_buf_1 _20409_ (.A(_04120_),
    .X(_04121_));
 sg13g2_nand2_1 _20410_ (.Y(_04122_),
    .A(_08184_),
    .B(_04060_));
 sg13g2_buf_1 _20411_ (.A(_04122_),
    .X(_04123_));
 sg13g2_nor2_1 _20412_ (.A(_04065_),
    .B(_04123_),
    .Y(_04124_));
 sg13g2_o21ai_1 _20413_ (.B1(_04064_),
    .Y(_04125_),
    .A1(_04121_),
    .A2(_04124_));
 sg13g2_o21ai_1 _20414_ (.B1(_04125_),
    .Y(_02527_),
    .A1(_04064_),
    .A2(_04117_));
 sg13g2_nand3_1 _20415_ (.B(_04065_),
    .C(_04062_),
    .A(_04064_),
    .Y(_04126_));
 sg13g2_a21oi_1 _20416_ (.A1(_04064_),
    .A2(_04065_),
    .Y(_04127_),
    .B1(_04123_));
 sg13g2_o21ai_1 _20417_ (.B1(\top_ihp.wb_emem.wait_counter[2] ),
    .Y(_04128_),
    .A1(_04121_),
    .A2(_04127_));
 sg13g2_o21ai_1 _20418_ (.B1(_04128_),
    .Y(_02528_),
    .A1(\top_ihp.wb_emem.wait_counter[2] ),
    .A2(_04126_));
 sg13g2_xnor2_1 _20419_ (.Y(_04129_),
    .A(_04063_),
    .B(_04066_));
 sg13g2_nand2_1 _20420_ (.Y(_04130_),
    .A(\top_ihp.wb_emem.wait_counter[3] ),
    .B(_04121_));
 sg13g2_o21ai_1 _20421_ (.B1(_04130_),
    .Y(_02529_),
    .A1(_04123_),
    .A2(_04129_));
 sg13g2_nand2_1 _20422_ (.Y(_04131_),
    .A(_04067_),
    .B(_04062_));
 sg13g2_nor2_1 _20423_ (.A(_04067_),
    .B(_04123_),
    .Y(_04132_));
 sg13g2_o21ai_1 _20424_ (.B1(_04069_),
    .Y(_04133_),
    .A1(_04121_),
    .A2(_04132_));
 sg13g2_o21ai_1 _20425_ (.B1(_04133_),
    .Y(_02530_),
    .A1(_04069_),
    .A2(_04131_));
 sg13g2_and2_1 _20426_ (.A(_04069_),
    .B(_04067_),
    .X(_04134_));
 sg13g2_buf_1 _20427_ (.A(_04134_),
    .X(_04135_));
 sg13g2_nand2_1 _20428_ (.Y(_04136_),
    .A(_04062_),
    .B(_04135_));
 sg13g2_nor2_1 _20429_ (.A(_04123_),
    .B(_04135_),
    .Y(_04137_));
 sg13g2_o21ai_1 _20430_ (.B1(_04068_),
    .Y(_04138_),
    .A1(_04121_),
    .A2(_04137_));
 sg13g2_o21ai_1 _20431_ (.B1(_04138_),
    .Y(_02531_),
    .A1(_04068_),
    .A2(_04136_));
 sg13g2_nand2_1 _20432_ (.Y(_04139_),
    .A(_04068_),
    .B(_04135_));
 sg13g2_xor2_1 _20433_ (.B(_04139_),
    .A(_04070_),
    .X(_04140_));
 sg13g2_nand2_1 _20434_ (.Y(_04141_),
    .A(_04070_),
    .B(_04121_));
 sg13g2_o21ai_1 _20435_ (.B1(_04141_),
    .Y(_02532_),
    .A1(_04123_),
    .A2(_04140_));
 sg13g2_o21ai_1 _20436_ (.B1(\top_ihp.wb_emem.wait_counter[7] ),
    .Y(_04142_),
    .A1(net945),
    .A2(_03763_));
 sg13g2_nand4_1 _20437_ (.B(_04070_),
    .C(_04062_),
    .A(_04068_),
    .Y(_04143_),
    .D(_04135_));
 sg13g2_mux2_1 _20438_ (.A0(\top_ihp.wb_emem.wait_counter[7] ),
    .A1(_04142_),
    .S(_04143_),
    .X(_04144_));
 sg13g2_inv_1 _20439_ (.Y(_02533_),
    .A(_04144_));
 sg13g2_mux4_1 _20440_ (.S0(_08173_),
    .A0(net8),
    .A1(net7),
    .A2(net6),
    .A3(net5),
    .S1(_08178_),
    .X(_04145_));
 sg13g2_nand2_1 _20441_ (.Y(_04146_),
    .A(_07673_),
    .B(_00003_));
 sg13g2_mux2_1 _20442_ (.A0(_04145_),
    .A1(\top_ihp.wb_dati_gpio[0] ),
    .S(_04146_),
    .X(_02534_));
 sg13g2_nor3_2 _20443_ (.A(_07677_),
    .B(_07673_),
    .C(_07712_),
    .Y(_04147_));
 sg13g2_nand3_1 _20444_ (.B(_08178_),
    .C(_04147_),
    .A(_08173_),
    .Y(_04148_));
 sg13g2_mux2_1 _20445_ (.A0(_03712_),
    .A1(\top_ihp.gpio_o_1 ),
    .S(_04148_),
    .X(_02535_));
 sg13g2_nand2_1 _20446_ (.Y(_04149_),
    .A(\top_ihp.oisc.wb_adr_o[0] ),
    .B(_08178_));
 sg13g2_mux2_1 _20447_ (.A0(_03712_),
    .A1(\top_ihp.gpio_o_2 ),
    .S(_04149_),
    .X(_04150_));
 sg13g2_inv_1 _20448_ (.Y(_04151_),
    .A(_04150_));
 sg13g2_mux2_1 _20449_ (.A0(_00222_),
    .A1(_04151_),
    .S(_04147_),
    .X(_02536_));
 sg13g2_inv_1 _20450_ (.Y(_04152_),
    .A(_00091_));
 sg13g2_nand3_1 _20451_ (.B(\top_ihp.oisc.wb_adr_o[1] ),
    .C(_04147_),
    .A(_08173_),
    .Y(_04153_));
 sg13g2_mux2_1 _20452_ (.A0(_04152_),
    .A1(\top_ihp.gpio_o_3 ),
    .S(_04153_),
    .X(_02537_));
 sg13g2_nor2_1 _20453_ (.A(_08173_),
    .B(_08178_),
    .Y(_04154_));
 sg13g2_mux2_1 _20454_ (.A0(\top_ihp.gpio_o_4 ),
    .A1(_03712_),
    .S(_04154_),
    .X(_04155_));
 sg13g2_inv_1 _20455_ (.Y(_04156_),
    .A(_04155_));
 sg13g2_mux2_1 _20456_ (.A0(_00223_),
    .A1(_04156_),
    .S(_04147_),
    .X(_02538_));
 sg13g2_nand2_1 _20457_ (.Y(_04157_),
    .A(_07713_),
    .B(_07741_));
 sg13g2_or2_1 _20458_ (.X(_04158_),
    .B(_07750_),
    .A(net884));
 sg13g2_buf_1 _20459_ (.A(_04158_),
    .X(_04159_));
 sg13g2_buf_1 _20460_ (.A(_04159_),
    .X(_04160_));
 sg13g2_buf_1 _20461_ (.A(net830),
    .X(_04161_));
 sg13g2_nand2_1 _20462_ (.Y(_04162_),
    .A(_04157_),
    .B(net815));
 sg13g2_nor3_1 _20463_ (.A(_07714_),
    .B(_07708_),
    .C(_07656_),
    .Y(_04163_));
 sg13g2_nor2_1 _20464_ (.A(net884),
    .B(_07750_),
    .Y(_04164_));
 sg13g2_nand3_1 _20465_ (.B(_07673_),
    .C(_07716_),
    .A(_07713_),
    .Y(_04165_));
 sg13g2_o21ai_1 _20466_ (.B1(_04165_),
    .Y(_04166_),
    .A1(_07713_),
    .A2(_04164_));
 sg13g2_a21oi_1 _20467_ (.A1(_07738_),
    .A2(_04163_),
    .Y(_04167_),
    .B1(_04166_));
 sg13g2_buf_1 _20468_ (.A(_04167_),
    .X(_04168_));
 sg13g2_buf_1 _20469_ (.A(_04168_),
    .X(_04169_));
 sg13g2_nand2_1 _20470_ (.Y(_04170_),
    .A(_07746_),
    .B(_04169_));
 sg13g2_o21ai_1 _20471_ (.B1(_04170_),
    .Y(_02539_),
    .A1(_07746_),
    .A2(_04162_));
 sg13g2_buf_1 _20472_ (.A(_04168_),
    .X(_04171_));
 sg13g2_buf_1 _20473_ (.A(_04171_),
    .X(_04172_));
 sg13g2_nor2b_1 _20474_ (.A(_07752_),
    .B_N(_09274_),
    .Y(_04173_));
 sg13g2_o21ai_1 _20475_ (.B1(_07754_),
    .Y(_04174_),
    .A1(_07750_),
    .A2(_04173_));
 sg13g2_nor2_1 _20476_ (.A(_07750_),
    .B(_04173_),
    .Y(_04175_));
 sg13g2_nor2b_1 _20477_ (.A(_04175_),
    .B_N(_07746_),
    .Y(_04176_));
 sg13g2_o21ai_1 _20478_ (.B1(_07745_),
    .Y(_04177_),
    .A1(_04171_),
    .A2(_04176_));
 sg13g2_o21ai_1 _20479_ (.B1(_04177_),
    .Y(_02540_),
    .A1(net628),
    .A2(_04174_));
 sg13g2_a21o_1 _20480_ (.A2(_07749_),
    .A1(_07752_),
    .B1(_04175_),
    .X(_04178_));
 sg13g2_buf_1 _20481_ (.A(_04178_),
    .X(_04179_));
 sg13g2_a21o_1 _20482_ (.A2(_04163_),
    .A1(_07738_),
    .B1(_04166_),
    .X(_04180_));
 sg13g2_buf_1 _20483_ (.A(_04180_),
    .X(_04181_));
 sg13g2_buf_1 _20484_ (.A(_04181_),
    .X(_04182_));
 sg13g2_nor3_1 _20485_ (.A(_07746_),
    .B(_07745_),
    .C(_07742_),
    .Y(_04183_));
 sg13g2_nor2b_1 _20486_ (.A(_07754_),
    .B_N(_07742_),
    .Y(_04184_));
 sg13g2_a21oi_1 _20487_ (.A1(_04182_),
    .A2(_04183_),
    .Y(_04185_),
    .B1(_04184_));
 sg13g2_nand2_1 _20488_ (.Y(_04186_),
    .A(_07742_),
    .B(_04169_));
 sg13g2_o21ai_1 _20489_ (.B1(_04186_),
    .Y(_02541_),
    .A1(_04179_),
    .A2(_04185_));
 sg13g2_nor2_1 _20490_ (.A(_04179_),
    .B(_04183_),
    .Y(_04187_));
 sg13g2_o21ai_1 _20491_ (.B1(\top_ihp.wb_imem.bits_left[3] ),
    .Y(_04188_),
    .A1(net661),
    .A2(_04187_));
 sg13g2_nor2b_1 _20492_ (.A(\top_ihp.wb_imem.bits_left[3] ),
    .B_N(_04183_),
    .Y(_04189_));
 sg13g2_nand2_1 _20493_ (.Y(_04190_),
    .A(_04181_),
    .B(_04189_));
 sg13g2_or2_1 _20494_ (.X(_04191_),
    .B(_04190_),
    .A(_04179_));
 sg13g2_nand2_1 _20495_ (.Y(_02542_),
    .A(_04188_),
    .B(_04191_));
 sg13g2_nor2_1 _20496_ (.A(_04179_),
    .B(_04189_),
    .Y(_04192_));
 sg13g2_o21ai_1 _20497_ (.B1(_07743_),
    .Y(_04193_),
    .A1(net661),
    .A2(_04192_));
 sg13g2_o21ai_1 _20498_ (.B1(_04193_),
    .Y(_02543_),
    .A1(_07743_),
    .A2(_04191_));
 sg13g2_buf_1 _20499_ (.A(_04164_),
    .X(_04194_));
 sg13g2_a221oi_1 _20500_ (.B2(_07744_),
    .C1(_04194_),
    .B1(_07754_),
    .A1(_07750_),
    .Y(_04195_),
    .A2(_07749_));
 sg13g2_o21ai_1 _20501_ (.B1(\top_ihp.wb_imem.bits_left[5] ),
    .Y(_04196_),
    .A1(_07743_),
    .A2(_04190_));
 sg13g2_o21ai_1 _20502_ (.B1(_04196_),
    .Y(_02544_),
    .A1(net628),
    .A2(_04195_));
 sg13g2_a22oi_1 _20503_ (.Y(_04197_),
    .B1(\top_ihp.oisc.wb_adr_o[0] ),
    .B2(net849),
    .A2(net2),
    .A1(net884));
 sg13g2_nand2_1 _20504_ (.Y(_04198_),
    .A(\top_ihp.wb_dati_rom[24] ),
    .B(net662));
 sg13g2_o21ai_1 _20505_ (.B1(_04198_),
    .Y(_02545_),
    .A1(net628),
    .A2(_04197_));
 sg13g2_buf_1 _20506_ (.A(_04159_),
    .X(_04199_));
 sg13g2_nor2_1 _20507_ (.A(_03951_),
    .B(_04199_),
    .Y(_04200_));
 sg13g2_a21oi_1 _20508_ (.A1(\top_ihp.wb_dati_rom[17] ),
    .A2(_04161_),
    .Y(_04201_),
    .B1(_04200_));
 sg13g2_nand2_1 _20509_ (.Y(_04202_),
    .A(\top_ihp.wb_dati_rom[18] ),
    .B(net662));
 sg13g2_o21ai_1 _20510_ (.B1(_04202_),
    .Y(_02546_),
    .A1(net628),
    .A2(_04201_));
 sg13g2_nor2_1 _20511_ (.A(_03953_),
    .B(_04199_),
    .Y(_04203_));
 sg13g2_a21oi_1 _20512_ (.A1(\top_ihp.wb_dati_rom[18] ),
    .A2(_04161_),
    .Y(_04204_),
    .B1(_04203_));
 sg13g2_nand2_1 _20513_ (.Y(_04205_),
    .A(\top_ihp.wb_dati_rom[19] ),
    .B(net662));
 sg13g2_o21ai_1 _20514_ (.B1(_04205_),
    .Y(_02547_),
    .A1(net628),
    .A2(_04204_));
 sg13g2_buf_1 _20515_ (.A(net830),
    .X(_04206_));
 sg13g2_nand2b_1 _20516_ (.Y(_04207_),
    .B(_04160_),
    .A_N(\top_ihp.wb_dati_rom[19] ));
 sg13g2_o21ai_1 _20517_ (.B1(_04207_),
    .Y(_04208_),
    .A1(_03956_),
    .A2(_04206_));
 sg13g2_nand2_1 _20518_ (.Y(_04209_),
    .A(\top_ihp.wb_dati_rom[20] ),
    .B(net662));
 sg13g2_o21ai_1 _20519_ (.B1(_04209_),
    .Y(_02548_),
    .A1(net628),
    .A2(_04208_));
 sg13g2_nor2_1 _20520_ (.A(_03962_),
    .B(net829),
    .Y(_04210_));
 sg13g2_a21oi_1 _20521_ (.A1(\top_ihp.wb_dati_rom[20] ),
    .A2(net815),
    .Y(_04211_),
    .B1(_04210_));
 sg13g2_nand2_1 _20522_ (.Y(_04212_),
    .A(\top_ihp.wb_dati_rom[21] ),
    .B(net662));
 sg13g2_o21ai_1 _20523_ (.B1(_04212_),
    .Y(_02549_),
    .A1(_04172_),
    .A2(_04211_));
 sg13g2_nor2_1 _20524_ (.A(_03967_),
    .B(net829),
    .Y(_04213_));
 sg13g2_a21oi_1 _20525_ (.A1(\top_ihp.wb_dati_rom[21] ),
    .A2(net815),
    .Y(_04214_),
    .B1(_04213_));
 sg13g2_nand2_1 _20526_ (.Y(_04215_),
    .A(\top_ihp.wb_dati_rom[22] ),
    .B(net662));
 sg13g2_o21ai_1 _20527_ (.B1(_04215_),
    .Y(_02550_),
    .A1(_04172_),
    .A2(_04214_));
 sg13g2_nand2_1 _20528_ (.Y(_04216_),
    .A(\top_ihp.wb_dati_rom[22] ),
    .B(net830));
 sg13g2_o21ai_1 _20529_ (.B1(_04216_),
    .Y(_04217_),
    .A1(_03971_),
    .A2(net814));
 sg13g2_mux2_1 _20530_ (.A0(\top_ihp.wb_dati_rom[23] ),
    .A1(_04217_),
    .S(net660),
    .X(_02551_));
 sg13g2_nor2_1 _20531_ (.A(_03976_),
    .B(net815),
    .Y(_04218_));
 sg13g2_o21ai_1 _20532_ (.B1(net660),
    .Y(_04219_),
    .A1(\top_ihp.wb_dati_rom[23] ),
    .A2(net849));
 sg13g2_nand2_1 _20533_ (.Y(_04220_),
    .A(\top_ihp.wb_dati_rom[8] ),
    .B(net662));
 sg13g2_o21ai_1 _20534_ (.B1(_04220_),
    .Y(_02552_),
    .A1(_04218_),
    .A2(_04219_));
 sg13g2_buf_1 _20535_ (.A(net661),
    .X(_04221_));
 sg13g2_nor2_1 _20536_ (.A(_03979_),
    .B(net829),
    .Y(_04222_));
 sg13g2_a21oi_1 _20537_ (.A1(\top_ihp.wb_dati_rom[8] ),
    .A2(net815),
    .Y(_04223_),
    .B1(_04222_));
 sg13g2_nand2_1 _20538_ (.Y(_04224_),
    .A(\top_ihp.wb_dati_rom[9] ),
    .B(net662));
 sg13g2_o21ai_1 _20539_ (.B1(_04224_),
    .Y(_02553_),
    .A1(net627),
    .A2(_04223_));
 sg13g2_nor2_1 _20540_ (.A(_03986_),
    .B(net829),
    .Y(_04225_));
 sg13g2_a21oi_1 _20541_ (.A1(\top_ihp.wb_dati_rom[9] ),
    .A2(net815),
    .Y(_04226_),
    .B1(_04225_));
 sg13g2_buf_1 _20542_ (.A(_04168_),
    .X(_04227_));
 sg13g2_nand2_1 _20543_ (.Y(_04228_),
    .A(\top_ihp.wb_dati_rom[10] ),
    .B(net659));
 sg13g2_o21ai_1 _20544_ (.B1(_04228_),
    .Y(_02554_),
    .A1(net627),
    .A2(_04226_));
 sg13g2_nand2_1 _20545_ (.Y(_04229_),
    .A(\top_ihp.wb_dati_rom[10] ),
    .B(net830));
 sg13g2_o21ai_1 _20546_ (.B1(_04229_),
    .Y(_04230_),
    .A1(_03988_),
    .A2(net814));
 sg13g2_mux2_1 _20547_ (.A0(\top_ihp.wb_dati_rom[11] ),
    .A1(_04230_),
    .S(net660),
    .X(_02555_));
 sg13g2_nor2_1 _20548_ (.A(_08178_),
    .B(net829),
    .Y(_04231_));
 sg13g2_a21oi_1 _20549_ (.A1(\top_ihp.wb_dati_rom[24] ),
    .A2(_04206_),
    .Y(_04232_),
    .B1(_04231_));
 sg13g2_nand2_1 _20550_ (.Y(_04233_),
    .A(\top_ihp.wb_dati_rom[25] ),
    .B(net659));
 sg13g2_o21ai_1 _20551_ (.B1(_04233_),
    .Y(_02556_),
    .A1(net627),
    .A2(_04232_));
 sg13g2_nor2_1 _20552_ (.A(_03992_),
    .B(net815),
    .Y(_04234_));
 sg13g2_o21ai_1 _20553_ (.B1(net660),
    .Y(_04235_),
    .A1(\top_ihp.wb_dati_rom[11] ),
    .A2(net849));
 sg13g2_nand2_1 _20554_ (.Y(_04236_),
    .A(\top_ihp.wb_dati_rom[12] ),
    .B(net659));
 sg13g2_o21ai_1 _20555_ (.B1(_04236_),
    .Y(_02557_),
    .A1(_04234_),
    .A2(_04235_));
 sg13g2_nor2_1 _20556_ (.A(\top_ihp.wb_dati_rom[12] ),
    .B(net849),
    .Y(_04237_));
 sg13g2_a21oi_1 _20557_ (.A1(_03998_),
    .A2(net849),
    .Y(_04238_),
    .B1(_04237_));
 sg13g2_mux2_1 _20558_ (.A0(\top_ihp.wb_dati_rom[13] ),
    .A1(_04238_),
    .S(net660),
    .X(_02558_));
 sg13g2_nand2_1 _20559_ (.Y(_04239_),
    .A(\top_ihp.wb_dati_rom[13] ),
    .B(net830));
 sg13g2_o21ai_1 _20560_ (.B1(_04239_),
    .Y(_04240_),
    .A1(_04005_),
    .A2(net814));
 sg13g2_mux2_1 _20561_ (.A0(\top_ihp.wb_dati_rom[14] ),
    .A1(_04240_),
    .S(net660),
    .X(_02559_));
 sg13g2_nor2_1 _20562_ (.A(_04008_),
    .B(net815),
    .Y(_04241_));
 sg13g2_o21ai_1 _20563_ (.B1(net660),
    .Y(_04242_),
    .A1(\top_ihp.wb_dati_rom[14] ),
    .A2(_04194_));
 sg13g2_nand2_1 _20564_ (.Y(_04243_),
    .A(\top_ihp.wb_dati_rom[15] ),
    .B(net659));
 sg13g2_o21ai_1 _20565_ (.B1(_04243_),
    .Y(_02560_),
    .A1(_04241_),
    .A2(_04242_));
 sg13g2_inv_1 _20566_ (.Y(_04244_),
    .A(\top_ihp.wb_dati_rom[0] ));
 sg13g2_a21oi_1 _20567_ (.A1(_07713_),
    .A2(_07741_),
    .Y(_04245_),
    .B1(_04164_));
 sg13g2_buf_2 _20568_ (.A(_04245_),
    .X(_04246_));
 sg13g2_inv_1 _20569_ (.Y(_04247_),
    .A(\top_ihp.wb_dati_rom[15] ));
 sg13g2_a22oi_1 _20570_ (.Y(_02561_),
    .B1(_04246_),
    .B2(_04247_),
    .A2(net628),
    .A1(_04244_));
 sg13g2_inv_1 _20571_ (.Y(_04248_),
    .A(\top_ihp.wb_dati_rom[1] ));
 sg13g2_a22oi_1 _20572_ (.Y(_02562_),
    .B1(_04246_),
    .B2(_04244_),
    .A2(net628),
    .A1(_04248_));
 sg13g2_nand2_1 _20573_ (.Y(_04249_),
    .A(\top_ihp.wb_dati_rom[2] ),
    .B(_04227_));
 sg13g2_o21ai_1 _20574_ (.B1(_04249_),
    .Y(_02563_),
    .A1(_04248_),
    .A2(_04162_));
 sg13g2_inv_1 _20575_ (.Y(_04250_),
    .A(\top_ihp.wb_dati_rom[3] ));
 sg13g2_nand2_1 _20576_ (.Y(_04251_),
    .A(\top_ihp.wb_dati_rom[2] ),
    .B(_04246_));
 sg13g2_o21ai_1 _20577_ (.B1(_04251_),
    .Y(_02564_),
    .A1(_04250_),
    .A2(net660));
 sg13g2_nand2_1 _20578_ (.Y(_04252_),
    .A(\top_ihp.wb_dati_rom[4] ),
    .B(_04227_));
 sg13g2_o21ai_1 _20579_ (.B1(_04252_),
    .Y(_02565_),
    .A1(_04250_),
    .A2(_04162_));
 sg13g2_and2_1 _20580_ (.A(\top_ihp.wb_dati_rom[5] ),
    .B(net661),
    .X(_04253_));
 sg13g2_a21o_1 _20581_ (.A2(_04246_),
    .A1(\top_ihp.wb_dati_rom[4] ),
    .B1(_04253_),
    .X(_02566_));
 sg13g2_nor2_1 _20582_ (.A(_03895_),
    .B(net829),
    .Y(_04254_));
 sg13g2_a21oi_1 _20583_ (.A1(\top_ihp.wb_dati_rom[25] ),
    .A2(net814),
    .Y(_04255_),
    .B1(_04254_));
 sg13g2_nand2_1 _20584_ (.Y(_04256_),
    .A(\top_ihp.wb_dati_rom[26] ),
    .B(net659));
 sg13g2_o21ai_1 _20585_ (.B1(_04256_),
    .Y(_02567_),
    .A1(_04221_),
    .A2(_04255_));
 sg13g2_and2_1 _20586_ (.A(\top_ihp.wb_dati_rom[6] ),
    .B(net661),
    .X(_04257_));
 sg13g2_a21o_1 _20587_ (.A2(_04246_),
    .A1(\top_ihp.wb_dati_rom[5] ),
    .B1(_04257_),
    .X(_02568_));
 sg13g2_and2_1 _20588_ (.A(\top_ihp.wb_dati_rom[7] ),
    .B(_04168_),
    .X(_04258_));
 sg13g2_a21o_1 _20589_ (.A2(_04246_),
    .A1(\top_ihp.wb_dati_rom[6] ),
    .B1(_04258_),
    .X(_02569_));
 sg13g2_nor2_1 _20590_ (.A(_03902_),
    .B(net829),
    .Y(_04259_));
 sg13g2_a21oi_1 _20591_ (.A1(\top_ihp.wb_dati_rom[26] ),
    .A2(net814),
    .Y(_04260_),
    .B1(_04259_));
 sg13g2_nand2_1 _20592_ (.Y(_04261_),
    .A(\top_ihp.wb_dati_rom[27] ),
    .B(net659));
 sg13g2_o21ai_1 _20593_ (.B1(_04261_),
    .Y(_02570_),
    .A1(_04221_),
    .A2(_04260_));
 sg13g2_and2_1 _20594_ (.A(\top_ihp.wb_dati_rom[27] ),
    .B(net830),
    .X(_04262_));
 sg13g2_a21oi_1 _20595_ (.A1(_03909_),
    .A2(net849),
    .Y(_04263_),
    .B1(_04262_));
 sg13g2_nand2_1 _20596_ (.Y(_04264_),
    .A(\top_ihp.wb_dati_rom[28] ),
    .B(net659));
 sg13g2_o21ai_1 _20597_ (.B1(_04264_),
    .Y(_02571_),
    .A1(net627),
    .A2(_04263_));
 sg13g2_and2_1 _20598_ (.A(\top_ihp.wb_dati_rom[28] ),
    .B(_04160_),
    .X(_04265_));
 sg13g2_a21oi_1 _20599_ (.A1(_03916_),
    .A2(net849),
    .Y(_04266_),
    .B1(_04265_));
 sg13g2_nand2_1 _20600_ (.Y(_04267_),
    .A(\top_ihp.wb_dati_rom[29] ),
    .B(net659));
 sg13g2_o21ai_1 _20601_ (.B1(_04267_),
    .Y(_02572_),
    .A1(net627),
    .A2(_04266_));
 sg13g2_nor2_1 _20602_ (.A(_03927_),
    .B(net829),
    .Y(_04268_));
 sg13g2_a21oi_1 _20603_ (.A1(\top_ihp.wb_dati_rom[29] ),
    .A2(net814),
    .Y(_04269_),
    .B1(_04268_));
 sg13g2_nand2_1 _20604_ (.Y(_04270_),
    .A(\top_ihp.wb_dati_rom[30] ),
    .B(net661));
 sg13g2_o21ai_1 _20605_ (.B1(_04270_),
    .Y(_02573_),
    .A1(net627),
    .A2(_04269_));
 sg13g2_nor2_1 _20606_ (.A(_03932_),
    .B(net830),
    .Y(_04271_));
 sg13g2_a21oi_1 _20607_ (.A1(\top_ihp.wb_dati_rom[30] ),
    .A2(net814),
    .Y(_04272_),
    .B1(_04271_));
 sg13g2_nand2_1 _20608_ (.Y(_04273_),
    .A(\top_ihp.wb_dati_rom[31] ),
    .B(net661));
 sg13g2_o21ai_1 _20609_ (.B1(_04273_),
    .Y(_02574_),
    .A1(net627),
    .A2(_04272_));
 sg13g2_nor2_1 _20610_ (.A(\top_ihp.wb_dati_rom[31] ),
    .B(_04164_),
    .Y(_04274_));
 sg13g2_a21oi_1 _20611_ (.A1(_03940_),
    .A2(net849),
    .Y(_04275_),
    .B1(_04274_));
 sg13g2_mux2_1 _20612_ (.A0(\top_ihp.wb_dati_rom[16] ),
    .A1(_04275_),
    .S(_04182_),
    .X(_02575_));
 sg13g2_nor2_1 _20613_ (.A(_03945_),
    .B(net830),
    .Y(_04276_));
 sg13g2_a21oi_1 _20614_ (.A1(\top_ihp.wb_dati_rom[16] ),
    .A2(net814),
    .Y(_04277_),
    .B1(_04276_));
 sg13g2_nand2_1 _20615_ (.Y(_04278_),
    .A(\top_ihp.wb_dati_rom[17] ),
    .B(net661));
 sg13g2_o21ai_1 _20616_ (.B1(_04278_),
    .Y(_02576_),
    .A1(net627),
    .A2(_04277_));
 sg13g2_nand4_1 _20617_ (.B(_07752_),
    .C(_07758_),
    .A(_09274_),
    .Y(_04279_),
    .D(_04157_));
 sg13g2_nand3_1 _20618_ (.B(_00224_),
    .C(_07741_),
    .A(_07713_),
    .Y(_04280_));
 sg13g2_nand3b_1 _20619_ (.B(_00224_),
    .C(net884),
    .Y(_04281_),
    .A_N(_07758_));
 sg13g2_nand2_1 _20620_ (.Y(_04282_),
    .A(_07713_),
    .B(_07752_));
 sg13g2_nand2_1 _20621_ (.Y(_04283_),
    .A(_07714_),
    .B(_00224_));
 sg13g2_o21ai_1 _20622_ (.B1(_04283_),
    .Y(_04284_),
    .A1(_07741_),
    .A2(_04282_));
 sg13g2_nand2b_1 _20623_ (.Y(_04285_),
    .B(_04284_),
    .A_N(net884));
 sg13g2_nand4_1 _20624_ (.B(_04280_),
    .C(_04281_),
    .A(_04279_),
    .Y(_02577_),
    .D(_04285_));
 sg13g2_nand2_1 _20625_ (.Y(_04286_),
    .A(_07651_),
    .B(_07664_));
 sg13g2_nand2_1 _20626_ (.Y(_04287_),
    .A(net807),
    .B(_07656_));
 sg13g2_inv_1 _20627_ (.Y(_04288_),
    .A(_00078_));
 sg13g2_a21oi_1 _20628_ (.A1(_07649_),
    .A2(_07656_),
    .Y(_04289_),
    .B1(_04288_));
 sg13g2_o21ai_1 _20629_ (.B1(_04289_),
    .Y(_04290_),
    .A1(_09671_),
    .A2(_04287_));
 sg13g2_buf_2 _20630_ (.A(_04290_),
    .X(_04291_));
 sg13g2_and2_1 _20631_ (.A(_04286_),
    .B(_04291_),
    .X(_04292_));
 sg13g2_buf_8 _20632_ (.A(_04292_),
    .X(_04293_));
 sg13g2_nand2_1 _20633_ (.Y(_04294_),
    .A(net983),
    .B(_04293_));
 sg13g2_nand2_1 _20634_ (.Y(_04295_),
    .A(_04286_),
    .B(_04291_));
 sg13g2_buf_2 _20635_ (.A(_04295_),
    .X(_04296_));
 sg13g2_buf_8 _20636_ (.A(_04296_),
    .X(_04297_));
 sg13g2_nand2_1 _20637_ (.Y(_04298_),
    .A(_07660_),
    .B(_04297_));
 sg13g2_o21ai_1 _20638_ (.B1(_04298_),
    .Y(_02578_),
    .A1(_07660_),
    .A2(_04294_));
 sg13g2_buf_1 _20639_ (.A(_04296_),
    .X(_04299_));
 sg13g2_or2_1 _20640_ (.X(_04300_),
    .B(\top_ihp.wb_spi.bits_left[1] ),
    .A(_07660_));
 sg13g2_buf_1 _20641_ (.A(_04300_),
    .X(_04301_));
 sg13g2_or2_1 _20642_ (.X(_04302_),
    .B(_04301_),
    .A(_07652_));
 sg13g2_buf_1 _20643_ (.A(_04302_),
    .X(_04303_));
 sg13g2_and2_1 _20644_ (.A(_07660_),
    .B(net1014),
    .X(_04304_));
 sg13g2_o21ai_1 _20645_ (.B1(\top_ihp.wb_spi.bits_left[1] ),
    .Y(_04305_),
    .A1(_04296_),
    .A2(_04304_));
 sg13g2_o21ai_1 _20646_ (.B1(_04305_),
    .Y(_02579_),
    .A1(net625),
    .A2(_04303_));
 sg13g2_nor3_1 _20647_ (.A(_07662_),
    .B(_07664_),
    .C(_04303_),
    .Y(_04306_));
 sg13g2_o21ai_1 _20648_ (.B1(net1014),
    .Y(_04307_),
    .A1(_07664_),
    .A2(_04301_));
 sg13g2_inv_1 _20649_ (.Y(_04308_),
    .A(_07662_));
 sg13g2_a21oi_1 _20650_ (.A1(_04291_),
    .A2(_04307_),
    .Y(_04309_),
    .B1(_04308_));
 sg13g2_a21o_1 _20651_ (.A2(_04306_),
    .A1(_04291_),
    .B1(_04309_),
    .X(_02580_));
 sg13g2_and3_1 _20652_ (.X(_04310_),
    .A(_07824_),
    .B(_07826_),
    .C(_09158_));
 sg13g2_buf_1 _20653_ (.A(_04310_),
    .X(_04311_));
 sg13g2_nor3_1 _20654_ (.A(_07662_),
    .B(\top_ihp.wb_spi.bits_left[3] ),
    .C(_04303_),
    .Y(_04312_));
 sg13g2_a21oi_1 _20655_ (.A1(_07652_),
    .A2(_04311_),
    .Y(_04313_),
    .B1(_04312_));
 sg13g2_nor3_1 _20656_ (.A(_07662_),
    .B(_07664_),
    .C(_04301_),
    .Y(_04314_));
 sg13g2_buf_1 _20657_ (.A(_07651_),
    .X(_04315_));
 sg13g2_nand2b_1 _20658_ (.Y(_04316_),
    .B(_04315_),
    .A_N(_04314_));
 sg13g2_inv_1 _20659_ (.Y(_04317_),
    .A(\top_ihp.wb_spi.bits_left[3] ));
 sg13g2_a21o_1 _20660_ (.A2(_04316_),
    .A1(_04291_),
    .B1(_04317_),
    .X(_04318_));
 sg13g2_o21ai_1 _20661_ (.B1(_04318_),
    .Y(_02581_),
    .A1(_04299_),
    .A2(_04313_));
 sg13g2_buf_8 _20662_ (.A(_04293_),
    .X(_04319_));
 sg13g2_buf_1 _20663_ (.A(net1014),
    .X(_04320_));
 sg13g2_nand2_1 _20664_ (.Y(_04321_),
    .A(_07666_),
    .B(_04312_));
 sg13g2_o21ai_1 _20665_ (.B1(_04321_),
    .Y(_04322_),
    .A1(net944),
    .A2(net801));
 sg13g2_buf_1 _20666_ (.A(net1014),
    .X(_04323_));
 sg13g2_nand2_1 _20667_ (.Y(_04324_),
    .A(_04317_),
    .B(_04314_));
 sg13g2_nand2_1 _20668_ (.Y(_04325_),
    .A(net943),
    .B(_04324_));
 sg13g2_a21oi_1 _20669_ (.A1(_04291_),
    .A2(_04325_),
    .Y(_04326_),
    .B1(_07666_));
 sg13g2_a21oi_1 _20670_ (.A1(net624),
    .A2(_04322_),
    .Y(_02582_),
    .B1(_04326_));
 sg13g2_buf_1 _20671_ (.A(_07828_),
    .X(_04327_));
 sg13g2_a22oi_1 _20672_ (.Y(_04328_),
    .B1(_04312_),
    .B2(_07667_),
    .A2(net800),
    .A1(_07652_));
 sg13g2_o21ai_1 _20673_ (.B1(net1014),
    .Y(_04329_),
    .A1(_07666_),
    .A2(_04324_));
 sg13g2_nand2_1 _20674_ (.Y(_04330_),
    .A(_04291_),
    .B(_04329_));
 sg13g2_nand2_1 _20675_ (.Y(_04331_),
    .A(\top_ihp.wb_spi.bits_left[5] ),
    .B(_04330_));
 sg13g2_o21ai_1 _20676_ (.B1(_04331_),
    .Y(_02583_),
    .A1(_04299_),
    .A2(_04328_));
 sg13g2_buf_1 _20677_ (.A(net800),
    .X(_04332_));
 sg13g2_buf_1 _20678_ (.A(_07651_),
    .X(_04333_));
 sg13g2_nor2_1 _20679_ (.A(_04333_),
    .B(_00091_),
    .Y(_04334_));
 sg13g2_a22oi_1 _20680_ (.Y(_04335_),
    .B1(_04332_),
    .B2(_04334_),
    .A2(net4),
    .A1(net983));
 sg13g2_buf_8 _20681_ (.A(_04293_),
    .X(_04336_));
 sg13g2_nor2_1 _20682_ (.A(\top_ihp.wb_dati_spi[0] ),
    .B(net623),
    .Y(_04337_));
 sg13g2_a21oi_1 _20683_ (.A1(_04319_),
    .A2(_04335_),
    .Y(_02584_),
    .B1(_04337_));
 sg13g2_nor2b_1 _20684_ (.A(net943),
    .B_N(_03718_),
    .Y(_04338_));
 sg13g2_a22oi_1 _20685_ (.Y(_04339_),
    .B1(net768),
    .B2(_04338_),
    .A2(\top_ihp.wb_dati_spi[9] ),
    .A1(net983));
 sg13g2_nor2_1 _20686_ (.A(\top_ihp.wb_dati_spi[10] ),
    .B(net623),
    .Y(_04340_));
 sg13g2_a21oi_1 _20687_ (.A1(net624),
    .A2(_04339_),
    .Y(_02585_),
    .B1(_04340_));
 sg13g2_nor2b_1 _20688_ (.A(net943),
    .B_N(_03721_),
    .Y(_04341_));
 sg13g2_a22oi_1 _20689_ (.Y(_04342_),
    .B1(net768),
    .B2(_04341_),
    .A2(\top_ihp.wb_dati_spi[10] ),
    .A1(net983));
 sg13g2_nor2_1 _20690_ (.A(\top_ihp.wb_dati_spi[11] ),
    .B(net623),
    .Y(_04343_));
 sg13g2_a21oi_1 _20691_ (.A1(net624),
    .A2(_04342_),
    .Y(_02586_),
    .B1(_04343_));
 sg13g2_buf_1 _20692_ (.A(_07674_),
    .X(_04344_));
 sg13g2_nor2b_1 _20693_ (.A(net942),
    .B_N(_03723_),
    .Y(_04345_));
 sg13g2_a22oi_1 _20694_ (.Y(_04346_),
    .B1(net768),
    .B2(_04345_),
    .A2(\top_ihp.wb_dati_spi[11] ),
    .A1(net983));
 sg13g2_nor2_1 _20695_ (.A(\top_ihp.wb_dati_spi[12] ),
    .B(net623),
    .Y(_04347_));
 sg13g2_a21oi_1 _20696_ (.A1(net624),
    .A2(_04346_),
    .Y(_02587_),
    .B1(_04347_));
 sg13g2_nor2b_1 _20697_ (.A(net942),
    .B_N(_03725_),
    .Y(_04348_));
 sg13g2_a22oi_1 _20698_ (.Y(_04349_),
    .B1(net768),
    .B2(_04348_),
    .A2(net944),
    .A1(\top_ihp.wb_dati_spi[12] ));
 sg13g2_nor2_1 _20699_ (.A(\top_ihp.wb_dati_spi[13] ),
    .B(net623),
    .Y(_04350_));
 sg13g2_a21oi_1 _20700_ (.A1(net624),
    .A2(_04349_),
    .Y(_02588_),
    .B1(_04350_));
 sg13g2_nor2b_1 _20701_ (.A(net942),
    .B_N(_03727_),
    .Y(_04351_));
 sg13g2_a22oi_1 _20702_ (.Y(_04352_),
    .B1(net768),
    .B2(_04351_),
    .A2(_04320_),
    .A1(\top_ihp.wb_dati_spi[13] ));
 sg13g2_nor2_1 _20703_ (.A(\top_ihp.wb_dati_spi[14] ),
    .B(net623),
    .Y(_04353_));
 sg13g2_a21oi_1 _20704_ (.A1(net624),
    .A2(_04352_),
    .Y(_02589_),
    .B1(_04353_));
 sg13g2_nor2b_1 _20705_ (.A(net942),
    .B_N(_03728_),
    .Y(_04354_));
 sg13g2_a22oi_1 _20706_ (.Y(_04355_),
    .B1(net768),
    .B2(_04354_),
    .A2(_04320_),
    .A1(\top_ihp.wb_dati_spi[14] ));
 sg13g2_buf_8 _20707_ (.A(_04293_),
    .X(_04356_));
 sg13g2_nor2_1 _20708_ (.A(\top_ihp.wb_dati_spi[15] ),
    .B(net622),
    .Y(_04357_));
 sg13g2_a21oi_1 _20709_ (.A1(net624),
    .A2(_04355_),
    .Y(_02590_),
    .B1(_04357_));
 sg13g2_nor2_1 _20710_ (.A(_07652_),
    .B(\top_ihp.wb_dati_spi[15] ),
    .Y(_04358_));
 sg13g2_buf_1 _20711_ (.A(_07828_),
    .X(_04359_));
 sg13g2_a221oi_1 _20712_ (.B2(_04152_),
    .C1(net1014),
    .B1(net801),
    .A1(\top_ihp.oisc.wb_dat_o[16] ),
    .Y(_04360_),
    .A2(_04359_));
 sg13g2_nor3_1 _20713_ (.A(_04296_),
    .B(_04358_),
    .C(_04360_),
    .Y(_04361_));
 sg13g2_a21o_1 _20714_ (.A2(_04297_),
    .A1(\top_ihp.wb_dati_spi[16] ),
    .B1(_04361_),
    .X(_02591_));
 sg13g2_inv_1 _20715_ (.Y(_04362_),
    .A(_00092_));
 sg13g2_a22oi_1 _20716_ (.Y(_04363_),
    .B1(_04084_),
    .B2(_04362_),
    .A2(net800),
    .A1(\top_ihp.oisc.wb_dat_o[17] ));
 sg13g2_nand2_1 _20717_ (.Y(_04364_),
    .A(_04344_),
    .B(\top_ihp.wb_dati_spi[16] ));
 sg13g2_o21ai_1 _20718_ (.B1(_04364_),
    .Y(_04365_),
    .A1(net943),
    .A2(_04363_));
 sg13g2_buf_8 _20719_ (.A(_04293_),
    .X(_04366_));
 sg13g2_mux2_1 _20720_ (.A0(\top_ihp.wb_dati_spi[17] ),
    .A1(_04365_),
    .S(_04366_),
    .X(_02592_));
 sg13g2_inv_1 _20721_ (.Y(_04367_),
    .A(_00093_));
 sg13g2_a22oi_1 _20722_ (.Y(_04368_),
    .B1(net801),
    .B2(_04367_),
    .A2(net800),
    .A1(\top_ihp.oisc.wb_dat_o[18] ));
 sg13g2_nand2_1 _20723_ (.Y(_04369_),
    .A(net942),
    .B(\top_ihp.wb_dati_spi[17] ));
 sg13g2_o21ai_1 _20724_ (.B1(_04369_),
    .Y(_04370_),
    .A1(net943),
    .A2(_04368_));
 sg13g2_mux2_1 _20725_ (.A0(\top_ihp.wb_dati_spi[18] ),
    .A1(_04370_),
    .S(net621),
    .X(_02593_));
 sg13g2_inv_1 _20726_ (.Y(_04371_),
    .A(_00094_));
 sg13g2_a22oi_1 _20727_ (.Y(_04372_),
    .B1(net801),
    .B2(_04371_),
    .A2(net799),
    .A1(\top_ihp.oisc.wb_dat_o[19] ));
 sg13g2_nand2_1 _20728_ (.Y(_04373_),
    .A(net942),
    .B(\top_ihp.wb_dati_spi[18] ));
 sg13g2_o21ai_1 _20729_ (.B1(_04373_),
    .Y(_04374_),
    .A1(net943),
    .A2(_04372_));
 sg13g2_mux2_1 _20730_ (.A0(\top_ihp.wb_dati_spi[19] ),
    .A1(_04374_),
    .S(_04366_),
    .X(_02594_));
 sg13g2_nor2_1 _20731_ (.A(_04333_),
    .B(_00092_),
    .Y(_04375_));
 sg13g2_a22oi_1 _20732_ (.Y(_04376_),
    .B1(_04332_),
    .B2(_04375_),
    .A2(\top_ihp.wb_dati_spi[0] ),
    .A1(net983));
 sg13g2_nor2_1 _20733_ (.A(\top_ihp.wb_dati_spi[1] ),
    .B(_04356_),
    .Y(_04377_));
 sg13g2_a21oi_1 _20734_ (.A1(_04319_),
    .A2(_04376_),
    .Y(_02595_),
    .B1(_04377_));
 sg13g2_inv_1 _20735_ (.Y(_04378_),
    .A(_00095_));
 sg13g2_a22oi_1 _20736_ (.Y(_04379_),
    .B1(net801),
    .B2(_04378_),
    .A2(_04359_),
    .A1(\top_ihp.oisc.wb_dat_o[20] ));
 sg13g2_nand2_1 _20737_ (.Y(_04380_),
    .A(_04344_),
    .B(\top_ihp.wb_dati_spi[19] ));
 sg13g2_o21ai_1 _20738_ (.B1(_04380_),
    .Y(_04381_),
    .A1(net943),
    .A2(_04379_));
 sg13g2_mux2_1 _20739_ (.A0(\top_ihp.wb_dati_spi[20] ),
    .A1(_04381_),
    .S(net623),
    .X(_02596_));
 sg13g2_inv_1 _20740_ (.Y(_04382_),
    .A(_00096_));
 sg13g2_a22oi_1 _20741_ (.Y(_04383_),
    .B1(net801),
    .B2(_04382_),
    .A2(net799),
    .A1(\top_ihp.oisc.wb_dat_o[21] ));
 sg13g2_nand2_1 _20742_ (.Y(_04384_),
    .A(net986),
    .B(\top_ihp.wb_dati_spi[20] ));
 sg13g2_o21ai_1 _20743_ (.B1(_04384_),
    .Y(_04385_),
    .A1(net943),
    .A2(_04383_));
 sg13g2_mux2_1 _20744_ (.A0(\top_ihp.wb_dati_spi[21] ),
    .A1(_04385_),
    .S(net623),
    .X(_02597_));
 sg13g2_inv_1 _20745_ (.Y(_04386_),
    .A(_00097_));
 sg13g2_a22oi_1 _20746_ (.Y(_04387_),
    .B1(net801),
    .B2(_04386_),
    .A2(net799),
    .A1(\top_ihp.oisc.wb_dat_o[22] ));
 sg13g2_nand2_1 _20747_ (.Y(_04388_),
    .A(net986),
    .B(\top_ihp.wb_dati_spi[21] ));
 sg13g2_o21ai_1 _20748_ (.B1(_04388_),
    .Y(_04389_),
    .A1(_04323_),
    .A2(_04387_));
 sg13g2_mux2_1 _20749_ (.A0(\top_ihp.wb_dati_spi[22] ),
    .A1(_04389_),
    .S(_04336_),
    .X(_02598_));
 sg13g2_inv_1 _20750_ (.Y(_04390_),
    .A(_00098_));
 sg13g2_a22oi_1 _20751_ (.Y(_04391_),
    .B1(net801),
    .B2(_04390_),
    .A2(net799),
    .A1(\top_ihp.oisc.wb_dat_o[23] ));
 sg13g2_nand2_1 _20752_ (.Y(_04392_),
    .A(net986),
    .B(\top_ihp.wb_dati_spi[22] ));
 sg13g2_o21ai_1 _20753_ (.B1(_04392_),
    .Y(_04393_),
    .A1(_04323_),
    .A2(_04391_));
 sg13g2_mux2_1 _20754_ (.A0(\top_ihp.wb_dati_spi[23] ),
    .A1(_04393_),
    .S(_04336_),
    .X(_02599_));
 sg13g2_buf_1 _20755_ (.A(net1014),
    .X(_04394_));
 sg13g2_nand2_1 _20756_ (.Y(_04395_),
    .A(\top_ihp.oisc.wb_dat_o[24] ),
    .B(net799));
 sg13g2_a22oi_1 _20757_ (.Y(_04396_),
    .B1(net813),
    .B2(_03712_),
    .A2(net816),
    .A1(_03758_));
 sg13g2_a21oi_1 _20758_ (.A1(_04395_),
    .A2(_04396_),
    .Y(_04397_),
    .B1(net987));
 sg13g2_a21oi_1 _20759_ (.A1(net941),
    .A2(\top_ihp.wb_dati_spi[23] ),
    .Y(_04398_),
    .B1(_04397_));
 sg13g2_nand2_1 _20760_ (.Y(_04399_),
    .A(\top_ihp.wb_dati_spi[24] ),
    .B(net626));
 sg13g2_o21ai_1 _20761_ (.B1(_04399_),
    .Y(_02600_),
    .A1(net625),
    .A2(_04398_));
 sg13g2_nand2_1 _20762_ (.Y(_04400_),
    .A(\top_ihp.oisc.wb_dat_o[25] ),
    .B(net799));
 sg13g2_a22oi_1 _20763_ (.Y(_04401_),
    .B1(net813),
    .B2(_03735_),
    .A2(_04083_),
    .A1(_03760_));
 sg13g2_a21oi_1 _20764_ (.A1(_04400_),
    .A2(_04401_),
    .Y(_04402_),
    .B1(net987));
 sg13g2_a21oi_1 _20765_ (.A1(net941),
    .A2(\top_ihp.wb_dati_spi[24] ),
    .Y(_04403_),
    .B1(_04402_));
 sg13g2_nand2_1 _20766_ (.Y(_04404_),
    .A(\top_ihp.wb_dati_spi[25] ),
    .B(net626));
 sg13g2_o21ai_1 _20767_ (.B1(_04404_),
    .Y(_02601_),
    .A1(net625),
    .A2(_04403_));
 sg13g2_nand2_1 _20768_ (.Y(_04405_),
    .A(\top_ihp.oisc.wb_dat_o[26] ),
    .B(net799));
 sg13g2_a22oi_1 _20769_ (.Y(_04406_),
    .B1(net813),
    .B2(_03745_),
    .A2(net816),
    .A1(_03718_));
 sg13g2_a21oi_1 _20770_ (.A1(_04405_),
    .A2(_04406_),
    .Y(_04407_),
    .B1(net987));
 sg13g2_a21oi_1 _20771_ (.A1(net944),
    .A2(\top_ihp.wb_dati_spi[25] ),
    .Y(_04408_),
    .B1(_04407_));
 sg13g2_nand2_1 _20772_ (.Y(_04409_),
    .A(\top_ihp.wb_dati_spi[26] ),
    .B(net626));
 sg13g2_o21ai_1 _20773_ (.B1(_04409_),
    .Y(_02602_),
    .A1(net625),
    .A2(_04408_));
 sg13g2_nand2_1 _20774_ (.Y(_04410_),
    .A(\top_ihp.oisc.wb_dat_o[27] ),
    .B(net799));
 sg13g2_a22oi_1 _20775_ (.Y(_04411_),
    .B1(net813),
    .B2(_03748_),
    .A2(net816),
    .A1(_03721_));
 sg13g2_a21oi_1 _20776_ (.A1(_04410_),
    .A2(_04411_),
    .Y(_04412_),
    .B1(net987));
 sg13g2_a21oi_1 _20777_ (.A1(net944),
    .A2(\top_ihp.wb_dati_spi[26] ),
    .Y(_04413_),
    .B1(_04412_));
 sg13g2_nand2_1 _20778_ (.Y(_04414_),
    .A(\top_ihp.wb_dati_spi[27] ),
    .B(net626));
 sg13g2_o21ai_1 _20779_ (.B1(_04414_),
    .Y(_02603_),
    .A1(net625),
    .A2(_04413_));
 sg13g2_nand2_1 _20780_ (.Y(_04415_),
    .A(\top_ihp.oisc.wb_dat_o[28] ),
    .B(_07828_));
 sg13g2_a22oi_1 _20781_ (.Y(_04416_),
    .B1(net813),
    .B2(_03750_),
    .A2(net816),
    .A1(_03723_));
 sg13g2_a21oi_1 _20782_ (.A1(_04415_),
    .A2(_04416_),
    .Y(_04417_),
    .B1(net987));
 sg13g2_a21oi_1 _20783_ (.A1(net944),
    .A2(\top_ihp.wb_dati_spi[27] ),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_nand2_1 _20784_ (.Y(_04419_),
    .A(\top_ihp.wb_dati_spi[28] ),
    .B(net626));
 sg13g2_o21ai_1 _20785_ (.B1(_04419_),
    .Y(_02604_),
    .A1(net625),
    .A2(_04418_));
 sg13g2_nand2_1 _20786_ (.Y(_04420_),
    .A(\top_ihp.oisc.wb_dat_o[29] ),
    .B(_07828_));
 sg13g2_a22oi_1 _20787_ (.Y(_04421_),
    .B1(net813),
    .B2(_03752_),
    .A2(net816),
    .A1(_03725_));
 sg13g2_a21oi_1 _20788_ (.A1(_04420_),
    .A2(_04421_),
    .Y(_04422_),
    .B1(net987));
 sg13g2_a21oi_1 _20789_ (.A1(net944),
    .A2(\top_ihp.wb_dati_spi[28] ),
    .Y(_04423_),
    .B1(_04422_));
 sg13g2_nand2_1 _20790_ (.Y(_04424_),
    .A(\top_ihp.wb_dati_spi[29] ),
    .B(net626));
 sg13g2_o21ai_1 _20791_ (.B1(_04424_),
    .Y(_02605_),
    .A1(net625),
    .A2(_04423_));
 sg13g2_nor2_1 _20792_ (.A(net986),
    .B(_00093_),
    .Y(_04425_));
 sg13g2_a22oi_1 _20793_ (.Y(_04426_),
    .B1(net768),
    .B2(_04425_),
    .A2(\top_ihp.wb_dati_spi[1] ),
    .A1(net941));
 sg13g2_nor2_1 _20794_ (.A(\top_ihp.wb_dati_spi[2] ),
    .B(net622),
    .Y(_04427_));
 sg13g2_a21oi_1 _20795_ (.A1(net624),
    .A2(_04426_),
    .Y(_02606_),
    .B1(_04427_));
 sg13g2_nand2_1 _20796_ (.Y(_04428_),
    .A(\top_ihp.oisc.wb_dat_o[30] ),
    .B(_07828_));
 sg13g2_a22oi_1 _20797_ (.Y(_04429_),
    .B1(net813),
    .B2(_03754_),
    .A2(net816),
    .A1(_03727_));
 sg13g2_a21oi_1 _20798_ (.A1(_04428_),
    .A2(_04429_),
    .Y(_04430_),
    .B1(net987));
 sg13g2_a21oi_1 _20799_ (.A1(net944),
    .A2(\top_ihp.wb_dati_spi[29] ),
    .Y(_04431_),
    .B1(_04430_));
 sg13g2_nand2_1 _20800_ (.Y(_04432_),
    .A(\top_ihp.wb_dati_spi[30] ),
    .B(net626));
 sg13g2_o21ai_1 _20801_ (.B1(_04432_),
    .Y(_02607_),
    .A1(net625),
    .A2(_04431_));
 sg13g2_nand2_1 _20802_ (.Y(_04433_),
    .A(\top_ihp.oisc.wb_dat_o[31] ),
    .B(_07828_));
 sg13g2_a22oi_1 _20803_ (.Y(_04434_),
    .B1(net813),
    .B2(_03756_),
    .A2(net816),
    .A1(_03728_));
 sg13g2_a21oi_1 _20804_ (.A1(_04433_),
    .A2(_04434_),
    .Y(_04435_),
    .B1(net987));
 sg13g2_a21oi_1 _20805_ (.A1(net944),
    .A2(\top_ihp.wb_dati_spi[30] ),
    .Y(_04436_),
    .B1(_04435_));
 sg13g2_nand2_1 _20806_ (.Y(_04437_),
    .A(\top_ihp.wb_dati_spi[31] ),
    .B(_04296_));
 sg13g2_o21ai_1 _20807_ (.B1(_04437_),
    .Y(_02608_),
    .A1(net626),
    .A2(_04436_));
 sg13g2_nor2_1 _20808_ (.A(net986),
    .B(_00094_),
    .Y(_04438_));
 sg13g2_a22oi_1 _20809_ (.Y(_04439_),
    .B1(net768),
    .B2(_04438_),
    .A2(\top_ihp.wb_dati_spi[2] ),
    .A1(net941));
 sg13g2_nor2_1 _20810_ (.A(\top_ihp.wb_dati_spi[3] ),
    .B(net622),
    .Y(_04440_));
 sg13g2_a21oi_1 _20811_ (.A1(net621),
    .A2(_04439_),
    .Y(_02609_),
    .B1(_04440_));
 sg13g2_nor2_1 _20812_ (.A(net986),
    .B(_00095_),
    .Y(_04441_));
 sg13g2_a22oi_1 _20813_ (.Y(_04442_),
    .B1(net800),
    .B2(_04441_),
    .A2(\top_ihp.wb_dati_spi[3] ),
    .A1(net941));
 sg13g2_nor2_1 _20814_ (.A(\top_ihp.wb_dati_spi[4] ),
    .B(net622),
    .Y(_04443_));
 sg13g2_a21oi_1 _20815_ (.A1(net621),
    .A2(_04442_),
    .Y(_02610_),
    .B1(_04443_));
 sg13g2_nor2_1 _20816_ (.A(net986),
    .B(_00096_),
    .Y(_04444_));
 sg13g2_a22oi_1 _20817_ (.Y(_04445_),
    .B1(net800),
    .B2(_04444_),
    .A2(\top_ihp.wb_dati_spi[4] ),
    .A1(net941));
 sg13g2_nor2_1 _20818_ (.A(\top_ihp.wb_dati_spi[5] ),
    .B(net622),
    .Y(_04446_));
 sg13g2_a21oi_1 _20819_ (.A1(net621),
    .A2(_04445_),
    .Y(_02611_),
    .B1(_04446_));
 sg13g2_nor2_1 _20820_ (.A(net986),
    .B(_00097_),
    .Y(_04447_));
 sg13g2_a22oi_1 _20821_ (.Y(_04448_),
    .B1(_04327_),
    .B2(_04447_),
    .A2(\top_ihp.wb_dati_spi[5] ),
    .A1(_04394_));
 sg13g2_nor2_1 _20822_ (.A(\top_ihp.wb_dati_spi[6] ),
    .B(net622),
    .Y(_04449_));
 sg13g2_a21oi_1 _20823_ (.A1(net621),
    .A2(_04448_),
    .Y(_02612_),
    .B1(_04449_));
 sg13g2_nor2_1 _20824_ (.A(_04315_),
    .B(_00098_),
    .Y(_04450_));
 sg13g2_a22oi_1 _20825_ (.Y(_04451_),
    .B1(net800),
    .B2(_04450_),
    .A2(\top_ihp.wb_dati_spi[6] ),
    .A1(net941));
 sg13g2_nor2_1 _20826_ (.A(\top_ihp.wb_dati_spi[7] ),
    .B(net622),
    .Y(_04452_));
 sg13g2_a21oi_1 _20827_ (.A1(net621),
    .A2(_04451_),
    .Y(_02613_),
    .B1(_04452_));
 sg13g2_nor2b_1 _20828_ (.A(net942),
    .B_N(_03758_),
    .Y(_04453_));
 sg13g2_a22oi_1 _20829_ (.Y(_04454_),
    .B1(_04327_),
    .B2(_04453_),
    .A2(\top_ihp.wb_dati_spi[7] ),
    .A1(_04394_));
 sg13g2_nor2_1 _20830_ (.A(\top_ihp.wb_dati_spi[8] ),
    .B(_04356_),
    .Y(_04455_));
 sg13g2_a21oi_1 _20831_ (.A1(net621),
    .A2(_04454_),
    .Y(_02614_),
    .B1(_04455_));
 sg13g2_nor2b_1 _20832_ (.A(net942),
    .B_N(_03760_),
    .Y(_04456_));
 sg13g2_a22oi_1 _20833_ (.Y(_04457_),
    .B1(net800),
    .B2(_04456_),
    .A2(\top_ihp.wb_dati_spi[8] ),
    .A1(net941));
 sg13g2_nor2_1 _20834_ (.A(\top_ihp.wb_dati_spi[9] ),
    .B(net622),
    .Y(_04458_));
 sg13g2_a21oi_1 _20835_ (.A1(net621),
    .A2(_04457_),
    .Y(_02615_),
    .B1(_04458_));
 sg13g2_nor2_1 _20836_ (.A(net983),
    .B(_03909_),
    .Y(_04459_));
 sg13g2_nand2_1 _20837_ (.Y(_04460_),
    .A(_07674_),
    .B(_07650_));
 sg13g2_o21ai_1 _20838_ (.B1(_07671_),
    .Y(_04461_),
    .A1(_04288_),
    .A2(_07656_));
 sg13g2_a21oi_2 _20839_ (.B1(_07670_),
    .Y(_04462_),
    .A2(_04461_),
    .A1(_04460_));
 sg13g2_mux2_1 _20840_ (.A0(_00225_),
    .A1(_04459_),
    .S(_04462_),
    .X(_02616_));
 sg13g2_nor2_1 _20841_ (.A(_07675_),
    .B(_03916_),
    .Y(_04463_));
 sg13g2_mux2_1 _20842_ (.A0(_00226_),
    .A1(_04463_),
    .S(_04462_),
    .X(_02617_));
 sg13g2_and2_1 _20843_ (.A(_07652_),
    .B(_03927_),
    .X(_04464_));
 sg13g2_mux2_1 _20844_ (.A0(_00227_),
    .A1(_04464_),
    .S(_04462_),
    .X(_02618_));
 sg13g2_buf_1 _20845_ (.A(\top_ihp.wb_uart.state[1] ),
    .X(_04465_));
 sg13g2_buf_1 _20846_ (.A(\top_ihp.wb_uart.rx_ready ),
    .X(_04466_));
 sg13g2_buf_1 _20847_ (.A(\top_ihp.wb_uart.tx_ready ),
    .X(_04467_));
 sg13g2_buf_1 _20848_ (.A(\top_ihp.wb_uart.state[0] ),
    .X(_04468_));
 sg13g2_nor2b_1 _20849_ (.A(_04465_),
    .B_N(_04468_),
    .Y(_04469_));
 sg13g2_a22oi_1 _20850_ (.Y(_04470_),
    .B1(_04467_),
    .B2(_04469_),
    .A2(_04466_),
    .A1(_04465_));
 sg13g2_nor2_1 _20851_ (.A(_08939_),
    .B(net992),
    .Y(_04471_));
 sg13g2_a21oi_1 _20852_ (.A1(_08939_),
    .A2(_04470_),
    .Y(_02619_),
    .B1(_04471_));
 sg13g2_mux2_1 _20853_ (.A0(_08083_),
    .A1(_04467_),
    .S(_04468_),
    .X(_04472_));
 sg13g2_nand3b_1 _20854_ (.B(_04468_),
    .C(_04465_),
    .Y(_04473_),
    .A_N(_04466_));
 sg13g2_o21ai_1 _20855_ (.B1(_04473_),
    .Y(_02620_),
    .A1(_04465_),
    .A2(_04472_));
 sg13g2_or2_1 _20856_ (.X(_04474_),
    .B(_04468_),
    .A(_04465_));
 sg13g2_nand2b_1 _20857_ (.Y(_04475_),
    .B(_04465_),
    .A_N(_04466_));
 sg13g2_o21ai_1 _20858_ (.B1(_04475_),
    .Y(_02621_),
    .A1(_07922_),
    .A2(_04474_));
 sg13g2_xnor2_1 _20859_ (.Y(_04476_),
    .A(_07928_),
    .B(net877));
 sg13g2_nor2_1 _20860_ (.A(_07943_),
    .B(_04476_),
    .Y(_02622_));
 sg13g2_inv_1 _20861_ (.Y(_04477_),
    .A(_07929_));
 sg13g2_nand2_1 _20862_ (.Y(_04478_),
    .A(_07928_),
    .B(net877));
 sg13g2_xnor2_1 _20863_ (.Y(_04479_),
    .A(_04477_),
    .B(_04478_));
 sg13g2_nor2_1 _20864_ (.A(_07943_),
    .B(_04479_),
    .Y(_02623_));
 sg13g2_nand3_1 _20865_ (.B(_07929_),
    .C(_07799_),
    .A(_07928_),
    .Y(_04480_));
 sg13g2_xor2_1 _20866_ (.B(_04480_),
    .A(_07926_),
    .X(_04481_));
 sg13g2_nor2_1 _20867_ (.A(_07943_),
    .B(_04481_),
    .Y(_02624_));
 sg13g2_nor3_1 _20868_ (.A(_04477_),
    .B(_00089_),
    .C(_07927_),
    .Y(_04482_));
 sg13g2_xnor2_1 _20869_ (.Y(_04483_),
    .A(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .B(_04482_));
 sg13g2_nor2_1 _20870_ (.A(_07943_),
    .B(_04483_),
    .Y(_02625_));
 sg13g2_inv_1 _20871_ (.Y(_04484_),
    .A(_07943_));
 sg13g2_and2_1 _20872_ (.A(_07795_),
    .B(_07794_),
    .X(_04485_));
 sg13g2_nor3_1 _20873_ (.A(_07787_),
    .B(_07777_),
    .C(_07784_),
    .Y(_04486_));
 sg13g2_nand4_1 _20874_ (.B(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ),
    .C(_07790_),
    .A(_07788_),
    .Y(_04487_),
    .D(_07791_));
 sg13g2_nor3_1 _20875_ (.A(_07786_),
    .B(_07796_),
    .C(_04487_),
    .Y(_04488_));
 sg13g2_nand4_1 _20876_ (.B(_04485_),
    .C(_04486_),
    .A(_04484_),
    .Y(_04489_),
    .D(_04488_));
 sg13g2_buf_1 _20877_ (.A(_04489_),
    .X(_04490_));
 sg13g2_nor2_1 _20878_ (.A(_07926_),
    .B(_04490_),
    .Y(_04491_));
 sg13g2_nor2_1 _20879_ (.A(_07928_),
    .B(_07929_),
    .Y(_04492_));
 sg13g2_nand2_1 _20880_ (.Y(_04493_),
    .A(_04491_),
    .B(_04492_));
 sg13g2_nand2_1 _20881_ (.Y(_04494_),
    .A(_00089_),
    .B(_07936_));
 sg13g2_nand2_1 _20882_ (.Y(_04495_),
    .A(\top_ihp.wb_dati_uart[0] ),
    .B(_04493_));
 sg13g2_o21ai_1 _20883_ (.B1(_04495_),
    .Y(_02626_),
    .A1(_04493_),
    .A2(_04494_));
 sg13g2_nand3_1 _20884_ (.B(_04477_),
    .C(_04491_),
    .A(_07928_),
    .Y(_04496_));
 sg13g2_nand2_1 _20885_ (.Y(_04497_),
    .A(\top_ihp.wb_dati_uart[1] ),
    .B(_04496_));
 sg13g2_o21ai_1 _20886_ (.B1(_04497_),
    .Y(_02627_),
    .A1(_07937_),
    .A2(_04496_));
 sg13g2_inv_1 _20887_ (.Y(_04498_),
    .A(_07928_));
 sg13g2_nand3_1 _20888_ (.B(_07929_),
    .C(_04491_),
    .A(_04498_),
    .Y(_04499_));
 sg13g2_nand2_1 _20889_ (.Y(_04500_),
    .A(\top_ihp.wb_dati_uart[2] ),
    .B(_04499_));
 sg13g2_o21ai_1 _20890_ (.B1(_04500_),
    .Y(_02628_),
    .A1(_07937_),
    .A2(_04499_));
 sg13g2_nand2b_1 _20891_ (.Y(_04501_),
    .B(_04491_),
    .A_N(_07930_));
 sg13g2_nand2_1 _20892_ (.Y(_04502_),
    .A(\top_ihp.wb_dati_uart[3] ),
    .B(_04501_));
 sg13g2_o21ai_1 _20893_ (.B1(_04502_),
    .Y(_02629_),
    .A1(_07937_),
    .A2(_04501_));
 sg13g2_inv_1 _20894_ (.Y(_04503_),
    .A(_04490_));
 sg13g2_nand2_1 _20895_ (.Y(_04504_),
    .A(_07926_),
    .B(_04503_));
 sg13g2_nand2_1 _20896_ (.Y(_04505_),
    .A(_07936_),
    .B(_04492_));
 sg13g2_nand2_1 _20897_ (.Y(_04506_),
    .A(_07926_),
    .B(_04492_));
 sg13g2_o21ai_1 _20898_ (.B1(_04506_),
    .Y(_04507_),
    .A1(_07926_),
    .A2(_07930_));
 sg13g2_nand2_1 _20899_ (.Y(_04508_),
    .A(_00089_),
    .B(_04507_));
 sg13g2_o21ai_1 _20900_ (.B1(\top_ihp.wb_dati_uart[4] ),
    .Y(_04509_),
    .A1(_04490_),
    .A2(_04508_));
 sg13g2_o21ai_1 _20901_ (.B1(_04509_),
    .Y(_02630_),
    .A1(_04504_),
    .A2(_04505_));
 sg13g2_nor3_1 _20902_ (.A(_04498_),
    .B(_07929_),
    .C(_04504_),
    .Y(_04510_));
 sg13g2_mux2_1 _20903_ (.A0(\top_ihp.wb_dati_uart[5] ),
    .A1(_07936_),
    .S(_04510_),
    .X(_02631_));
 sg13g2_nor3_1 _20904_ (.A(_07928_),
    .B(_04477_),
    .C(_04504_),
    .Y(_04511_));
 sg13g2_mux2_1 _20905_ (.A0(\top_ihp.wb_dati_uart[6] ),
    .A1(_07936_),
    .S(_04511_),
    .X(_02632_));
 sg13g2_nor2_1 _20906_ (.A(_07930_),
    .B(_04504_),
    .Y(_04512_));
 sg13g2_mux2_1 _20907_ (.A0(\top_ihp.wb_dati_uart[7] ),
    .A1(_07936_),
    .S(_04512_),
    .X(_02633_));
 sg13g2_nand2_1 _20908_ (.Y(_04513_),
    .A(_07925_),
    .B(_07944_));
 sg13g2_a21oi_1 _20909_ (.A1(_07788_),
    .A2(_00079_),
    .Y(_04514_),
    .B1(_07976_));
 sg13g2_a21o_1 _20910_ (.A2(_04514_),
    .A1(_07796_),
    .B1(_04488_),
    .X(_04515_));
 sg13g2_a22oi_1 _20911_ (.Y(_04516_),
    .B1(_04515_),
    .B2(_04485_),
    .A2(_04514_),
    .A1(_04487_));
 sg13g2_a21oi_1 _20912_ (.A1(_04486_),
    .A2(_04516_),
    .Y(_04517_),
    .B1(_07945_));
 sg13g2_a21o_1 _20913_ (.A2(_04513_),
    .A1(_04466_),
    .B1(_04517_),
    .X(_02634_));
 sg13g2_nand2_2 _20914_ (.Y(_04518_),
    .A(net1024),
    .B(_08041_));
 sg13g2_xnor2_1 _20915_ (.Y(_04519_),
    .A(_08043_),
    .B(_08079_));
 sg13g2_nor2_1 _20916_ (.A(_04518_),
    .B(_04519_),
    .Y(_02635_));
 sg13g2_nand2_1 _20917_ (.Y(_04520_),
    .A(_08043_),
    .B(_08079_));
 sg13g2_xor2_1 _20918_ (.B(_04520_),
    .A(_08044_),
    .X(_04521_));
 sg13g2_nor2_1 _20919_ (.A(_04518_),
    .B(_04521_),
    .Y(_02636_));
 sg13g2_o21ai_1 _20920_ (.B1(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .Y(_04522_),
    .A1(_08060_),
    .A2(_08077_));
 sg13g2_nand2_1 _20921_ (.Y(_04523_),
    .A(_08043_),
    .B(_08044_));
 sg13g2_xor2_1 _20922_ (.B(_04523_),
    .A(_00090_),
    .X(_04524_));
 sg13g2_nand2_1 _20923_ (.Y(_04525_),
    .A(_08079_),
    .B(_04524_));
 sg13g2_a21oi_1 _20924_ (.A1(_04522_),
    .A2(_04525_),
    .Y(_02637_),
    .B1(_04518_));
 sg13g2_xor2_1 _20925_ (.B(_08080_),
    .A(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ),
    .X(_04526_));
 sg13g2_nor2_1 _20926_ (.A(_04518_),
    .B(_04526_),
    .Y(_02638_));
 sg13g2_mux2_1 _20927_ (.A0(_03712_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ),
    .S(_08090_),
    .X(_02639_));
 sg13g2_mux2_1 _20928_ (.A0(_03735_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ),
    .S(net551),
    .X(_02640_));
 sg13g2_mux2_1 _20929_ (.A0(_03745_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ),
    .S(net551),
    .X(_02641_));
 sg13g2_mux2_1 _20930_ (.A0(_03748_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ),
    .S(net551),
    .X(_02642_));
 sg13g2_mux2_1 _20931_ (.A0(_03750_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ),
    .S(net551),
    .X(_02643_));
 sg13g2_mux2_1 _20932_ (.A0(_03752_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ),
    .S(net551),
    .X(_02644_));
 sg13g2_mux2_1 _20933_ (.A0(_03754_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ),
    .S(net551),
    .X(_02645_));
 sg13g2_mux2_1 _20934_ (.A0(_03756_),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ),
    .S(net551),
    .X(_02646_));
 sg13g2_nand2b_1 _20935_ (.Y(_04527_),
    .B(_08040_),
    .A_N(_04467_));
 sg13g2_o21ai_1 _20936_ (.B1(_04527_),
    .Y(_04528_),
    .A1(_08040_),
    .A2(_08083_));
 sg13g2_o21ai_1 _20937_ (.B1(net1024),
    .Y(_04529_),
    .A1(_04467_),
    .A2(_08087_));
 sg13g2_o21ai_1 _20938_ (.B1(_04529_),
    .Y(_02647_),
    .A1(net1024),
    .A2(_04528_));
 sg13g2_nand2_1 _20939_ (.Y(_04530_),
    .A(_09734_),
    .B(_09825_));
 sg13g2_buf_2 _20940_ (.A(_04530_),
    .X(_04531_));
 sg13g2_buf_1 _20941_ (.A(net804),
    .X(_04532_));
 sg13g2_buf_1 _20942_ (.A(_09383_),
    .X(_04533_));
 sg13g2_buf_1 _20943_ (.A(_09827_),
    .X(_04534_));
 sg13g2_nor3_1 _20944_ (.A(net980),
    .B(_09844_),
    .C(_09848_),
    .Y(_04535_));
 sg13g2_a221oi_1 _20945_ (.B2(_09363_),
    .C1(_04535_),
    .B1(net804),
    .A1(_09152_),
    .Y(_04536_),
    .A2(\top_ihp.wb_dati_uart[5] ));
 sg13g2_nand3_1 _20946_ (.B(_09883_),
    .C(_09884_),
    .A(_09389_),
    .Y(_04537_));
 sg13g2_nor4_1 _20947_ (.A(_09732_),
    .B(net732),
    .C(_04536_),
    .D(_04537_),
    .Y(_04538_));
 sg13g2_nor3_1 _20948_ (.A(_08218_),
    .B(_09818_),
    .C(_09822_),
    .Y(_04539_));
 sg13g2_a221oi_1 _20949_ (.B2(_09851_),
    .C1(_04539_),
    .B1(_09850_),
    .A1(_09152_),
    .Y(_04540_),
    .A2(\top_ihp.wb_dati_uart[4] ));
 sg13g2_buf_1 _20950_ (.A(_04540_),
    .X(_04541_));
 sg13g2_and2_1 _20951_ (.A(_09885_),
    .B(_04541_),
    .X(_04542_));
 sg13g2_o21ai_1 _20952_ (.B1(_09790_),
    .Y(_04543_),
    .A1(_04538_),
    .A2(_04542_));
 sg13g2_buf_2 _20953_ (.A(_04543_),
    .X(_04544_));
 sg13g2_inv_2 _20954_ (.Y(_04545_),
    .A(_04544_));
 sg13g2_nor2_1 _20955_ (.A(net733),
    .B(_04545_),
    .Y(_04546_));
 sg13g2_buf_1 _20956_ (.A(_09357_),
    .X(_04547_));
 sg13g2_nor2_1 _20957_ (.A(_04536_),
    .B(_04537_),
    .Y(_04548_));
 sg13g2_a221oi_1 _20958_ (.B2(_04548_),
    .C1(_09391_),
    .B1(_09790_),
    .A1(net767),
    .Y(_04549_),
    .A2(net798));
 sg13g2_a21oi_1 _20959_ (.A1(net767),
    .A2(_04546_),
    .Y(_04550_),
    .B1(_04549_));
 sg13g2_nor3_1 _20960_ (.A(net804),
    .B(_09357_),
    .C(_09383_),
    .Y(_04551_));
 sg13g2_buf_1 _20961_ (.A(_09732_),
    .X(_04552_));
 sg13g2_nand2_1 _20962_ (.Y(_04553_),
    .A(_09827_),
    .B(_09853_));
 sg13g2_buf_2 _20963_ (.A(_04553_),
    .X(_04554_));
 sg13g2_nand2b_1 _20964_ (.Y(_04555_),
    .B(_09885_),
    .A_N(_09790_));
 sg13g2_nand4_1 _20965_ (.B(_09825_),
    .C(_09883_),
    .A(_09790_),
    .Y(_04556_),
    .D(_09884_));
 sg13g2_o21ai_1 _20966_ (.B1(_04556_),
    .Y(_04557_),
    .A1(_04554_),
    .A2(_04555_));
 sg13g2_buf_1 _20967_ (.A(_04557_),
    .X(_04558_));
 sg13g2_and2_1 _20968_ (.A(net708),
    .B(_04558_),
    .X(_04559_));
 sg13g2_nor2_2 _20969_ (.A(_04551_),
    .B(_04559_),
    .Y(_04560_));
 sg13g2_nand2_1 _20970_ (.Y(_04561_),
    .A(net798),
    .B(net733));
 sg13g2_buf_1 _20971_ (.A(_04544_),
    .X(_04562_));
 sg13g2_nand2_1 _20972_ (.Y(_04563_),
    .A(_09734_),
    .B(_04541_));
 sg13g2_or2_1 _20973_ (.X(_04564_),
    .B(_04563_),
    .A(net620));
 sg13g2_a21o_1 _20974_ (.A2(_04561_),
    .A1(_04560_),
    .B1(_04564_),
    .X(_04565_));
 sg13g2_o21ai_1 _20975_ (.B1(_04565_),
    .Y(_04566_),
    .A1(_04531_),
    .A2(_04550_));
 sg13g2_buf_1 _20976_ (.A(net771),
    .X(_04567_));
 sg13g2_mux2_1 _20977_ (.A0(\top_ihp.oisc.decoder.decoded[0] ),
    .A1(_04566_),
    .S(net731),
    .X(_00231_));
 sg13g2_a21oi_1 _20978_ (.A1(net767),
    .A2(net798),
    .Y(_04568_),
    .B1(_04563_));
 sg13g2_nand3_1 _20979_ (.B(_04546_),
    .C(_04568_),
    .A(net771),
    .Y(_04569_));
 sg13g2_o21ai_1 _20980_ (.B1(_04569_),
    .Y(_00232_),
    .A1(_07653_),
    .A2(net731));
 sg13g2_buf_1 _20981_ (.A(_09825_),
    .X(_04570_));
 sg13g2_buf_1 _20982_ (.A(_09363_),
    .X(_04571_));
 sg13g2_nor2_2 _20983_ (.A(net804),
    .B(_09383_),
    .Y(_04572_));
 sg13g2_o21ai_1 _20984_ (.B1(net736),
    .Y(_04573_),
    .A1(net766),
    .A2(_04572_));
 sg13g2_nor4_1 _20985_ (.A(_08223_),
    .B(net708),
    .C(net730),
    .D(_04573_),
    .Y(_04574_));
 sg13g2_a21o_1 _20986_ (.A2(net775),
    .A1(_07420_),
    .B1(_04574_),
    .X(_00233_));
 sg13g2_nor2_1 _20987_ (.A(_09058_),
    .B(net771),
    .Y(_04575_));
 sg13g2_o21ai_1 _20988_ (.B1(net708),
    .Y(_04576_),
    .A1(_04551_),
    .A2(_04558_));
 sg13g2_a21oi_1 _20989_ (.A1(net732),
    .A2(net736),
    .Y(_04577_),
    .B1(_04576_));
 sg13g2_a21oi_1 _20990_ (.A1(net732),
    .A2(_04573_),
    .Y(_04578_),
    .B1(net708));
 sg13g2_nor4_1 _20991_ (.A(net805),
    .B(_04545_),
    .C(_04577_),
    .D(_04578_),
    .Y(_04579_));
 sg13g2_buf_1 _20992_ (.A(_09734_),
    .X(_04580_));
 sg13g2_xnor2_1 _20993_ (.Y(_04581_),
    .A(net707),
    .B(net732));
 sg13g2_nor2_1 _20994_ (.A(_04560_),
    .B(_04581_),
    .Y(_04582_));
 sg13g2_nand2_1 _20995_ (.Y(_04583_),
    .A(net804),
    .B(_09363_));
 sg13g2_nor3_1 _20996_ (.A(_09391_),
    .B(_04531_),
    .C(_04583_),
    .Y(_04584_));
 sg13g2_or3_1 _20997_ (.A(net805),
    .B(_04544_),
    .C(_04584_),
    .X(_04585_));
 sg13g2_buf_1 _20998_ (.A(_04585_),
    .X(_04586_));
 sg13g2_a21oi_1 _20999_ (.A1(_09853_),
    .A2(_04582_),
    .Y(_04587_),
    .B1(_04586_));
 sg13g2_nor3_1 _21000_ (.A(_04575_),
    .B(_04579_),
    .C(_04587_),
    .Y(_00234_));
 sg13g2_nand3_1 _21001_ (.B(_04570_),
    .C(net736),
    .A(_04532_),
    .Y(_04588_));
 sg13g2_nand2_1 _21002_ (.Y(_04589_),
    .A(_09363_),
    .B(_09734_));
 sg13g2_a21oi_1 _21003_ (.A1(_04554_),
    .A2(_04588_),
    .Y(_04590_),
    .B1(_04589_));
 sg13g2_nor2_1 _21004_ (.A(net798),
    .B(_04534_),
    .Y(_04591_));
 sg13g2_nand2_1 _21005_ (.Y(_04592_),
    .A(_04552_),
    .B(_04591_));
 sg13g2_a21oi_1 _21006_ (.A1(_04563_),
    .A2(_04592_),
    .Y(_04593_),
    .B1(net767));
 sg13g2_nor2_1 _21007_ (.A(_04590_),
    .B(_04593_),
    .Y(_04594_));
 sg13g2_nor2_1 _21008_ (.A(net733),
    .B(_04594_),
    .Y(_04595_));
 sg13g2_and3_1 _21009_ (.X(_04596_),
    .A(_04552_),
    .B(_04570_),
    .C(_04558_));
 sg13g2_o21ai_1 _21010_ (.B1(net620),
    .Y(_04597_),
    .A1(_04595_),
    .A2(_04596_));
 sg13g2_a21oi_1 _21011_ (.A1(_09855_),
    .A2(_04584_),
    .Y(_04598_),
    .B1(_08223_));
 sg13g2_a22oi_1 _21012_ (.Y(_00235_),
    .B1(_04597_),
    .B2(_04598_),
    .A2(net738),
    .A1(_09114_));
 sg13g2_nand2_1 _21013_ (.Y(_04599_),
    .A(net804),
    .B(_04591_));
 sg13g2_o21ai_1 _21014_ (.B1(_04599_),
    .Y(_04600_),
    .A1(net730),
    .A2(_04544_));
 sg13g2_nand2_1 _21015_ (.Y(_04601_),
    .A(net733),
    .B(_04600_));
 sg13g2_nand2_1 _21016_ (.Y(_04602_),
    .A(net730),
    .B(_04572_));
 sg13g2_o21ai_1 _21017_ (.B1(_04602_),
    .Y(_04603_),
    .A1(net730),
    .A2(_04544_));
 sg13g2_a22oi_1 _21018_ (.Y(_04604_),
    .B1(_04603_),
    .B2(net766),
    .A2(net620),
    .A1(net730));
 sg13g2_a221oi_1 _21019_ (.B2(_04604_),
    .C1(net708),
    .B1(_04601_),
    .A1(_09850_),
    .Y(_04605_),
    .A2(_09851_));
 sg13g2_nor3_1 _21020_ (.A(_04580_),
    .B(net732),
    .C(_04560_),
    .Y(_04606_));
 sg13g2_o21ai_1 _21021_ (.B1(net771),
    .Y(_04607_),
    .A1(_04605_),
    .A2(_04606_));
 sg13g2_o21ai_1 _21022_ (.B1(_04607_),
    .Y(_00236_),
    .A1(_09119_),
    .A2(net731));
 sg13g2_nor2_1 _21023_ (.A(net708),
    .B(net732),
    .Y(_04608_));
 sg13g2_o21ai_1 _21024_ (.B1(_04608_),
    .Y(_04609_),
    .A1(net798),
    .A2(net733));
 sg13g2_o21ai_1 _21025_ (.B1(_04609_),
    .Y(_04610_),
    .A1(_04560_),
    .A2(_04581_));
 sg13g2_o21ai_1 _21026_ (.B1(net620),
    .Y(_04611_),
    .A1(_04531_),
    .A2(_04583_));
 sg13g2_a21oi_1 _21027_ (.A1(_09853_),
    .A2(_04610_),
    .Y(_04612_),
    .B1(_04611_));
 sg13g2_nand2_1 _21028_ (.Y(_04613_),
    .A(_09363_),
    .B(_04572_));
 sg13g2_nor3_1 _21029_ (.A(net736),
    .B(_04531_),
    .C(_04613_),
    .Y(_04614_));
 sg13g2_nand2_1 _21030_ (.Y(_04615_),
    .A(_09206_),
    .B(net805));
 sg13g2_o21ai_1 _21031_ (.B1(_04615_),
    .Y(_04616_),
    .A1(_04586_),
    .A2(_04614_));
 sg13g2_a21oi_1 _21032_ (.A1(net731),
    .A2(_04612_),
    .Y(_00237_),
    .B1(_04616_));
 sg13g2_nor2_1 _21033_ (.A(_04554_),
    .B(_04576_),
    .Y(_04617_));
 sg13g2_nor2_1 _21034_ (.A(_09391_),
    .B(_04563_),
    .Y(_04618_));
 sg13g2_nor3_1 _21035_ (.A(_04586_),
    .B(_04617_),
    .C(_04618_),
    .Y(_04619_));
 sg13g2_o21ai_1 _21036_ (.B1(_09383_),
    .Y(_04620_),
    .A1(_09732_),
    .A2(_04541_));
 sg13g2_nand2_1 _21037_ (.Y(_04621_),
    .A(net766),
    .B(_04620_));
 sg13g2_a21oi_1 _21038_ (.A1(net767),
    .A2(net708),
    .Y(_04622_),
    .B1(_04621_));
 sg13g2_xnor2_1 _21039_ (.Y(_04623_),
    .A(net732),
    .B(net736));
 sg13g2_or3_1 _21040_ (.A(net951),
    .B(_09326_),
    .C(_09330_),
    .X(_04624_));
 sg13g2_buf_2 _21041_ (.A(_04624_),
    .X(_04625_));
 sg13g2_nand2_1 _21042_ (.Y(_04626_),
    .A(_04625_),
    .B(_09825_));
 sg13g2_nand4_1 _21043_ (.B(net707),
    .C(_04620_),
    .A(net766),
    .Y(_04627_),
    .D(_04626_));
 sg13g2_o21ai_1 _21044_ (.B1(_04627_),
    .Y(_04628_),
    .A1(net707),
    .A2(_04623_));
 sg13g2_o21ai_1 _21045_ (.B1(_04628_),
    .Y(_04629_),
    .A1(_04558_),
    .A2(_04622_));
 sg13g2_nand2_1 _21046_ (.Y(_04630_),
    .A(_09383_),
    .B(_04534_));
 sg13g2_o21ai_1 _21047_ (.B1(_09391_),
    .Y(_04631_),
    .A1(_04532_),
    .A2(_04591_));
 sg13g2_nand3_1 _21048_ (.B(_04630_),
    .C(_04631_),
    .A(net707),
    .Y(_04632_));
 sg13g2_nand4_1 _21049_ (.B(net620),
    .C(_04629_),
    .A(_03696_),
    .Y(_04633_),
    .D(_04632_));
 sg13g2_o21ai_1 _21050_ (.B1(_04633_),
    .Y(_04634_),
    .A1(\top_ihp.oisc.decoder.decoded[1] ),
    .A2(net771));
 sg13g2_nor2_1 _21051_ (.A(_04619_),
    .B(_04634_),
    .Y(_00238_));
 sg13g2_nand3_1 _21052_ (.B(net736),
    .C(_04559_),
    .A(net730),
    .Y(_04635_));
 sg13g2_nand2_1 _21053_ (.Y(_04636_),
    .A(_09332_),
    .B(net730));
 sg13g2_nor4_1 _21054_ (.A(_09383_),
    .B(_09853_),
    .C(_04556_),
    .D(_04636_),
    .Y(_04637_));
 sg13g2_a21oi_1 _21055_ (.A1(_09383_),
    .A2(_09853_),
    .Y(_04638_),
    .B1(net730));
 sg13g2_nand4_1 _21056_ (.B(_09825_),
    .C(net736),
    .A(net708),
    .Y(_04639_),
    .D(_04572_));
 sg13g2_o21ai_1 _21057_ (.B1(_04639_),
    .Y(_04640_),
    .A1(_04625_),
    .A2(_04531_));
 sg13g2_a21o_1 _21058_ (.A2(_04638_),
    .A1(net707),
    .B1(_04640_),
    .X(_04641_));
 sg13g2_o21ai_1 _21059_ (.B1(net766),
    .Y(_04642_),
    .A1(_04637_),
    .A2(_04641_));
 sg13g2_nand4_1 _21060_ (.B(net707),
    .C(net732),
    .A(net798),
    .Y(_04643_),
    .D(_04572_));
 sg13g2_nand4_1 _21061_ (.B(_04635_),
    .C(_04642_),
    .A(net620),
    .Y(_04644_),
    .D(_04643_));
 sg13g2_o21ai_1 _21062_ (.B1(_04613_),
    .Y(_04645_),
    .A1(_04625_),
    .A2(_04630_));
 sg13g2_nand3_1 _21063_ (.B(_09853_),
    .C(_04645_),
    .A(_04580_),
    .Y(_04646_));
 sg13g2_a21oi_1 _21064_ (.A1(_04545_),
    .A2(_04646_),
    .Y(_04647_),
    .B1(net776));
 sg13g2_a22oi_1 _21065_ (.Y(_04648_),
    .B1(_04644_),
    .B2(_04647_),
    .A2(net776),
    .A1(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_inv_1 _21066_ (.Y(_00239_),
    .A(_04648_));
 sg13g2_xnor2_1 _21067_ (.Y(_04649_),
    .A(_04625_),
    .B(net798));
 sg13g2_a21oi_1 _21068_ (.A1(_04618_),
    .A2(_04649_),
    .Y(_04650_),
    .B1(_04617_));
 sg13g2_nor2_1 _21069_ (.A(net767),
    .B(net766),
    .Y(_04651_));
 sg13g2_a22oi_1 _21070_ (.Y(_04652_),
    .B1(_04651_),
    .B2(_04630_),
    .A2(_04638_),
    .A1(net766));
 sg13g2_nand3b_1 _21071_ (.B(net707),
    .C(net620),
    .Y(_04653_),
    .A_N(_04652_));
 sg13g2_o21ai_1 _21072_ (.B1(_04653_),
    .Y(_04654_),
    .A1(net620),
    .A2(_04650_));
 sg13g2_mux2_1 _21073_ (.A0(\top_ihp.oisc.decoder.decoded[3] ),
    .A1(_04654_),
    .S(_04567_),
    .X(_00240_));
 sg13g2_o21ai_1 _21074_ (.B1(_09332_),
    .Y(_04655_),
    .A1(_04541_),
    .A2(_04591_));
 sg13g2_o21ai_1 _21075_ (.B1(_04655_),
    .Y(_04656_),
    .A1(net798),
    .A2(_04554_));
 sg13g2_nand3_1 _21076_ (.B(net707),
    .C(_04656_),
    .A(net733),
    .Y(_04657_));
 sg13g2_o21ai_1 _21077_ (.B1(_04657_),
    .Y(_04658_),
    .A1(_04554_),
    .A2(_04560_));
 sg13g2_nor2_1 _21078_ (.A(_04571_),
    .B(_04531_),
    .Y(_04659_));
 sg13g2_or4_1 _21079_ (.A(_04545_),
    .B(_04584_),
    .C(_04617_),
    .D(_04659_),
    .X(_04660_));
 sg13g2_o21ai_1 _21080_ (.B1(_04660_),
    .Y(_04661_),
    .A1(_04562_),
    .A2(_04658_));
 sg13g2_nand2_1 _21081_ (.Y(_04662_),
    .A(\top_ihp.oisc.decoder.decoded[4] ),
    .B(_08225_));
 sg13g2_o21ai_1 _21082_ (.B1(_04662_),
    .Y(_00241_),
    .A1(net738),
    .A2(_04661_));
 sg13g2_nor2_1 _21083_ (.A(net733),
    .B(_04544_),
    .Y(_04663_));
 sg13g2_nor2_1 _21084_ (.A(net767),
    .B(_04554_),
    .Y(_04664_));
 sg13g2_nor2_1 _21085_ (.A(_04636_),
    .B(_04663_),
    .Y(_04665_));
 sg13g2_a21oi_1 _21086_ (.A1(_04663_),
    .A2(_04664_),
    .Y(_04666_),
    .B1(_04665_));
 sg13g2_nand4_1 _21087_ (.B(net733),
    .C(_04608_),
    .A(_04625_),
    .Y(_04667_),
    .D(_04562_));
 sg13g2_o21ai_1 _21088_ (.B1(_04667_),
    .Y(_04668_),
    .A1(_04589_),
    .A2(_04666_));
 sg13g2_mux2_1 _21089_ (.A0(\top_ihp.oisc.decoder.decoded[5] ),
    .A1(_04668_),
    .S(_04567_),
    .X(_00242_));
 sg13g2_inv_1 _21090_ (.Y(_04669_),
    .A(\top_ihp.oisc.decoder.decoded[6] ));
 sg13g2_nor2_1 _21091_ (.A(_04571_),
    .B(_04533_),
    .Y(_04670_));
 sg13g2_a21oi_1 _21092_ (.A1(_04625_),
    .A2(_04533_),
    .Y(_04671_),
    .B1(_04670_));
 sg13g2_nor3_1 _21093_ (.A(_04531_),
    .B(_04545_),
    .C(_04671_),
    .Y(_04672_));
 sg13g2_a21oi_1 _21094_ (.A1(_09391_),
    .A2(_04583_),
    .Y(_04673_),
    .B1(_04564_));
 sg13g2_nor3_1 _21095_ (.A(net776),
    .B(_04672_),
    .C(_04673_),
    .Y(_04674_));
 sg13g2_a21oi_1 _21096_ (.A1(_04669_),
    .A2(net738),
    .Y(_00243_),
    .B1(_04674_));
 sg13g2_o21ai_1 _21097_ (.B1(_04545_),
    .Y(_04675_),
    .A1(_04547_),
    .A2(_09391_));
 sg13g2_a22oi_1 _21098_ (.Y(_04676_),
    .B1(_04675_),
    .B2(net767),
    .A2(_04546_),
    .A1(_04547_));
 sg13g2_nor3_1 _21099_ (.A(net776),
    .B(_04531_),
    .C(_04676_),
    .Y(_04677_));
 sg13g2_a21o_1 _21100_ (.A2(_08225_),
    .A1(\top_ihp.oisc.decoder.decoded[7] ),
    .B1(_04677_),
    .X(_00244_));
 sg13g2_buf_1 _21101_ (.A(net771),
    .X(_04678_));
 sg13g2_mux2_1 _21102_ (.A0(_09096_),
    .A1(_09253_),
    .S(net729),
    .X(_00245_));
 sg13g2_mux2_1 _21103_ (.A0(_09087_),
    .A1(_09277_),
    .S(net729),
    .X(_00246_));
 sg13g2_nand2_1 _21104_ (.Y(_04679_),
    .A(net988),
    .B(net775));
 sg13g2_o21ai_1 _21105_ (.B1(_04679_),
    .Y(_00247_),
    .A1(net738),
    .A2(_04625_));
 sg13g2_nand2_1 _21106_ (.Y(_04680_),
    .A(net917),
    .B(net775));
 sg13g2_o21ai_1 _21107_ (.B1(_04680_),
    .Y(_00248_),
    .A1(net738),
    .A2(net766));
 sg13g2_nand2_1 _21108_ (.Y(_04681_),
    .A(_09241_),
    .B(net775));
 sg13g2_o21ai_1 _21109_ (.B1(_04681_),
    .Y(_00249_),
    .A1(net738),
    .A2(_09391_));
 sg13g2_inv_1 _21110_ (.Y(_04682_),
    .A(\top_ihp.oisc.decoder.instruction[16] ));
 sg13g2_or4_1 _21111_ (.A(_07647_),
    .B(_08243_),
    .C(_09131_),
    .D(_09133_),
    .X(_04683_));
 sg13g2_buf_1 _21112_ (.A(_04683_),
    .X(_04684_));
 sg13g2_o21ai_1 _21113_ (.B1(_04684_),
    .Y(_00250_),
    .A1(_04682_),
    .A2(net731));
 sg13g2_inv_1 _21114_ (.Y(_04685_),
    .A(\top_ihp.oisc.decoder.instruction[17] ));
 sg13g2_or4_1 _21115_ (.A(_07647_),
    .B(_08243_),
    .C(_09448_),
    .D(_09449_),
    .X(_04686_));
 sg13g2_buf_1 _21116_ (.A(_04686_),
    .X(_04687_));
 sg13g2_o21ai_1 _21117_ (.B1(_04687_),
    .Y(_00251_),
    .A1(_04685_),
    .A2(net731));
 sg13g2_inv_1 _21118_ (.Y(_04688_),
    .A(\top_ihp.oisc.decoder.instruction[18] ));
 sg13g2_or4_1 _21119_ (.A(_07647_),
    .B(_08243_),
    .C(_09471_),
    .D(_09472_),
    .X(_04689_));
 sg13g2_buf_1 _21120_ (.A(_04689_),
    .X(_04690_));
 sg13g2_o21ai_1 _21121_ (.B1(_04690_),
    .Y(_00252_),
    .A1(_04688_),
    .A2(net731));
 sg13g2_nor4_1 _21122_ (.A(net984),
    .B(net823),
    .C(_09499_),
    .D(_09501_),
    .Y(_04691_));
 sg13g2_a21o_1 _21123_ (.A2(net775),
    .A1(\top_ihp.oisc.decoder.instruction[19] ),
    .B1(_04691_),
    .X(_00253_));
 sg13g2_nand2_1 _21124_ (.Y(_04692_),
    .A(net771),
    .B(_09569_));
 sg13g2_o21ai_1 _21125_ (.B1(_04692_),
    .Y(_00254_),
    .A1(_09116_),
    .A2(net731));
 sg13g2_mux2_1 _21126_ (.A0(_09542_),
    .A1(_09589_),
    .S(net729),
    .X(_00255_));
 sg13g2_mux2_1 _21127_ (.A0(_09615_),
    .A1(_09606_),
    .S(_04678_),
    .X(_00256_));
 sg13g2_nand2_1 _21128_ (.Y(_04693_),
    .A(_09625_),
    .B(net775));
 sg13g2_o21ai_1 _21129_ (.B1(_04693_),
    .Y(_00257_),
    .A1(net738),
    .A2(_09217_));
 sg13g2_mux2_1 _21130_ (.A0(_09649_),
    .A1(_09172_),
    .S(net729),
    .X(_00258_));
 sg13g2_mux2_1 _21131_ (.A0(_09663_),
    .A1(_09520_),
    .S(net729),
    .X(_00259_));
 sg13g2_mux2_1 _21132_ (.A0(_09672_),
    .A1(_09257_),
    .S(net729),
    .X(_00260_));
 sg13g2_nand2_1 _21133_ (.Y(_04694_),
    .A(\top_ihp.oisc.decoder.instruction[27] ),
    .B(net776));
 sg13g2_o21ai_1 _21134_ (.B1(_04694_),
    .Y(_00261_),
    .A1(_08224_),
    .A2(_09285_));
 sg13g2_mux2_1 _21135_ (.A0(_09705_),
    .A1(_09340_),
    .S(net729),
    .X(_00262_));
 sg13g2_mux2_1 _21136_ (.A0(\top_ihp.oisc.decoder.instruction[29] ),
    .A1(_09361_),
    .S(net729),
    .X(_00263_));
 sg13g2_mux2_1 _21137_ (.A0(\top_ihp.oisc.decoder.instruction[30] ),
    .A1(_09389_),
    .S(_04678_),
    .X(_00264_));
 sg13g2_nand2_1 _21138_ (.Y(_04695_),
    .A(_09295_),
    .B(net776));
 sg13g2_o21ai_1 _21139_ (.B1(_04695_),
    .Y(_00265_),
    .A1(_08224_),
    .A2(_09235_));
 sg13g2_nand2_1 _21140_ (.Y(_04696_),
    .A(_09225_),
    .B(_09902_));
 sg13g2_mux2_1 _21141_ (.A0(_09074_),
    .A1(_04696_),
    .S(net771),
    .X(_00266_));
 sg13g2_mux2_1 _21142_ (.A0(_09055_),
    .A1(_09177_),
    .S(_03697_),
    .X(_00267_));
 sg13g2_nand2_1 _21143_ (.Y(_04697_),
    .A(_09099_),
    .B(net776));
 sg13g2_o21ai_1 _21144_ (.B1(_04697_),
    .Y(_00268_),
    .A1(net775),
    .A2(_09526_));
 sg13g2_nand3b_1 _21145_ (.B(_09061_),
    .C(\top_ihp.oisc.decoder.decoded[15] ),
    .Y(_04698_),
    .A_N(_09060_));
 sg13g2_buf_1 _21146_ (.A(_04698_),
    .X(_04699_));
 sg13g2_nand3b_1 _21147_ (.B(_04699_),
    .C(net998),
    .Y(_04700_),
    .A_N(_00099_));
 sg13g2_buf_1 _21148_ (.A(_04700_),
    .X(_04701_));
 sg13g2_inv_1 _21149_ (.Y(_04702_),
    .A(\top_ihp.oisc.micro_op[13] ));
 sg13g2_nand3b_1 _21150_ (.B(_07422_),
    .C(_08228_),
    .Y(_04703_),
    .A_N(_09070_));
 sg13g2_buf_1 _21151_ (.A(_04703_),
    .X(_04704_));
 sg13g2_or2_1 _21152_ (.X(_04705_),
    .B(_04704_),
    .A(_04702_));
 sg13g2_buf_1 _21153_ (.A(_04705_),
    .X(_04706_));
 sg13g2_nand2_1 _21154_ (.Y(_04707_),
    .A(_04701_),
    .B(_04706_));
 sg13g2_o21ai_1 _21155_ (.B1(_04707_),
    .Y(_04708_),
    .A1(net984),
    .A2(_08243_));
 sg13g2_a21oi_1 _21156_ (.A1(_04684_),
    .A2(_04708_),
    .Y(_04709_),
    .B1(_09089_));
 sg13g2_buf_8 _21157_ (.A(_04709_),
    .X(_04710_));
 sg13g2_nand2_1 _21158_ (.Y(_04711_),
    .A(_08228_),
    .B(_07422_));
 sg13g2_nor2_2 _21159_ (.A(_09070_),
    .B(_04711_),
    .Y(_04712_));
 sg13g2_and2_1 _21160_ (.A(net998),
    .B(_04699_),
    .X(_04713_));
 sg13g2_inv_1 _21161_ (.Y(_04714_),
    .A(_00101_));
 sg13g2_a22oi_1 _21162_ (.Y(_04715_),
    .B1(_04713_),
    .B2(_04714_),
    .A2(_04712_),
    .A1(\top_ihp.oisc.micro_op[15] ));
 sg13g2_buf_2 _21163_ (.A(_04715_),
    .X(_04716_));
 sg13g2_a21o_1 _21164_ (.A2(net845),
    .A1(_07417_),
    .B1(_04716_),
    .X(_04717_));
 sg13g2_buf_1 _21165_ (.A(_04717_),
    .X(_04718_));
 sg13g2_a21oi_1 _21166_ (.A1(_04690_),
    .A2(_04718_),
    .Y(_04719_),
    .B1(net997));
 sg13g2_buf_8 _21167_ (.A(_04719_),
    .X(_04720_));
 sg13g2_nor2_1 _21168_ (.A(net728),
    .B(net727),
    .Y(_04721_));
 sg13g2_buf_2 _21169_ (.A(_04721_),
    .X(_04722_));
 sg13g2_inv_1 _21170_ (.Y(_04723_),
    .A(_09089_));
 sg13g2_nand3_1 _21171_ (.B(_04723_),
    .C(net845),
    .A(net1017),
    .Y(_04724_));
 sg13g2_nand3_1 _21172_ (.B(\top_ihp.oisc.decoder.instruction[20] ),
    .C(_04699_),
    .A(net998),
    .Y(_04725_));
 sg13g2_buf_1 _21173_ (.A(_04725_),
    .X(_04726_));
 sg13g2_inv_1 _21174_ (.Y(_04727_),
    .A(\top_ihp.oisc.micro_op[12] ));
 sg13g2_or2_1 _21175_ (.X(_04728_),
    .B(_04704_),
    .A(_04727_));
 sg13g2_buf_1 _21176_ (.A(_04728_),
    .X(_04729_));
 sg13g2_and3_1 _21177_ (.X(_04730_),
    .A(_04723_),
    .B(_04726_),
    .C(_04729_));
 sg13g2_o21ai_1 _21178_ (.B1(_04730_),
    .Y(_04731_),
    .A1(net984),
    .A2(net823));
 sg13g2_o21ai_1 _21179_ (.B1(_04731_),
    .Y(_04732_),
    .A1(_09406_),
    .A2(_04724_));
 sg13g2_buf_2 _21180_ (.A(_04732_),
    .X(_04733_));
 sg13g2_a21oi_1 _21181_ (.A1(net728),
    .A2(net727),
    .Y(_04734_),
    .B1(_04733_));
 sg13g2_nor2_1 _21182_ (.A(_09083_),
    .B(_00102_),
    .Y(_04735_));
 sg13g2_nand2_1 _21183_ (.Y(_04736_),
    .A(_04699_),
    .B(_04735_));
 sg13g2_nand3_1 _21184_ (.B(_04712_),
    .C(_04736_),
    .A(net805),
    .Y(_04737_));
 sg13g2_inv_1 _21185_ (.Y(_04738_),
    .A(\top_ihp.oisc.micro_op[14] ));
 sg13g2_inv_1 _21186_ (.Y(_04739_),
    .A(_00100_));
 sg13g2_nand3_1 _21187_ (.B(_04739_),
    .C(_04699_),
    .A(_09071_),
    .Y(_04740_));
 sg13g2_o21ai_1 _21188_ (.B1(_04740_),
    .Y(_04741_),
    .A1(_04738_),
    .A2(_04704_));
 sg13g2_o21ai_1 _21189_ (.B1(_04741_),
    .Y(_04742_),
    .A1(_07647_),
    .A2(_08243_));
 sg13g2_a21oi_1 _21190_ (.A1(_04687_),
    .A2(_04742_),
    .Y(_04743_),
    .B1(_09089_));
 sg13g2_buf_8 _21191_ (.A(_04743_),
    .X(_04744_));
 sg13g2_a21oi_1 _21192_ (.A1(_04723_),
    .A2(_04737_),
    .Y(_04745_),
    .B1(net726));
 sg13g2_o21ai_1 _21193_ (.B1(_04745_),
    .Y(_04746_),
    .A1(_04722_),
    .A2(_04734_));
 sg13g2_a21o_1 _21194_ (.A2(_04708_),
    .A1(_04684_),
    .B1(net997),
    .X(_04747_));
 sg13g2_buf_4 _21195_ (.X(_04748_),
    .A(_04747_));
 sg13g2_or4_1 _21196_ (.A(net984),
    .B(net823),
    .C(_09499_),
    .D(_09501_),
    .X(_04749_));
 sg13g2_and2_1 _21197_ (.A(_04699_),
    .B(_04735_),
    .X(_04750_));
 sg13g2_buf_1 _21198_ (.A(_04750_),
    .X(_04751_));
 sg13g2_o21ai_1 _21199_ (.B1(_04751_),
    .Y(_04752_),
    .A1(net984),
    .A2(net823));
 sg13g2_a21oi_1 _21200_ (.A1(_04749_),
    .A2(_04752_),
    .Y(_04753_),
    .B1(net997));
 sg13g2_buf_1 _21201_ (.A(_04753_),
    .X(_04754_));
 sg13g2_nor2_1 _21202_ (.A(_04748_),
    .B(_04754_),
    .Y(_04755_));
 sg13g2_a21oi_1 _21203_ (.A1(net805),
    .A2(_04712_),
    .Y(_04756_),
    .B1(net997));
 sg13g2_nor2_1 _21204_ (.A(net727),
    .B(_04756_),
    .Y(_04757_));
 sg13g2_a21o_1 _21205_ (.A2(_04742_),
    .A1(_04687_),
    .B1(net997),
    .X(_04758_));
 sg13g2_buf_8 _21206_ (.A(_04758_),
    .X(_04759_));
 sg13g2_and3_1 _21207_ (.X(_04760_),
    .A(_04723_),
    .B(net724),
    .C(_04737_));
 sg13g2_o21ai_1 _21208_ (.B1(_04760_),
    .Y(_04761_),
    .A1(_04755_),
    .A2(_04757_));
 sg13g2_nor2_1 _21209_ (.A(net726),
    .B(_04748_),
    .Y(_04762_));
 sg13g2_buf_2 _21210_ (.A(_04762_),
    .X(_04763_));
 sg13g2_nor2_1 _21211_ (.A(net724),
    .B(net728),
    .Y(_04764_));
 sg13g2_buf_2 _21212_ (.A(_04764_),
    .X(_04765_));
 sg13g2_a21o_1 _21213_ (.A2(_04718_),
    .A1(_04690_),
    .B1(_09089_),
    .X(_04766_));
 sg13g2_buf_8 _21214_ (.A(_04766_),
    .X(_04767_));
 sg13g2_nor2_1 _21215_ (.A(_09089_),
    .B(_04704_),
    .Y(_04768_));
 sg13g2_nand4_1 _21216_ (.B(_04726_),
    .C(_04729_),
    .A(_04736_),
    .Y(_04769_),
    .D(_04768_));
 sg13g2_a21o_1 _21217_ (.A2(net845),
    .A1(_07417_),
    .B1(_04769_),
    .X(_04770_));
 sg13g2_buf_1 _21218_ (.A(_04770_),
    .X(_04771_));
 sg13g2_buf_8 _21219_ (.A(_04771_),
    .X(_04772_));
 sg13g2_nor2_1 _21220_ (.A(net723),
    .B(net765),
    .Y(_04773_));
 sg13g2_o21ai_1 _21221_ (.B1(_04773_),
    .Y(_04774_),
    .A1(_04763_),
    .A2(_04765_));
 sg13g2_nand3_1 _21222_ (.B(_04761_),
    .C(_04774_),
    .A(_04746_),
    .Y(_04775_));
 sg13g2_buf_8 _21223_ (.A(_04748_),
    .X(_04776_));
 sg13g2_buf_8 _21224_ (.A(net706),
    .X(_04777_));
 sg13g2_nor2_2 _21225_ (.A(_04716_),
    .B(net765),
    .Y(_04778_));
 sg13g2_nand2_1 _21226_ (.Y(_04779_),
    .A(_04726_),
    .B(_04729_));
 sg13g2_inv_1 _21227_ (.Y(_04780_),
    .A(_04768_));
 sg13g2_a21oi_1 _21228_ (.A1(_07418_),
    .A2(net845),
    .Y(_04781_),
    .B1(_04780_));
 sg13g2_buf_2 _21229_ (.A(_04781_),
    .X(_04782_));
 sg13g2_nand3_1 _21230_ (.B(_04779_),
    .C(_04782_),
    .A(_04751_),
    .Y(_04783_));
 sg13g2_buf_1 _21231_ (.A(_04783_),
    .X(_04784_));
 sg13g2_nor4_1 _21232_ (.A(_09071_),
    .B(_04727_),
    .C(_04711_),
    .D(_04751_),
    .Y(_04785_));
 sg13g2_a21oi_1 _21233_ (.A1(net805),
    .A2(_04785_),
    .Y(_04786_),
    .B1(_09090_));
 sg13g2_buf_2 _21234_ (.A(_04786_),
    .X(_04787_));
 sg13g2_o21ai_1 _21235_ (.B1(_04787_),
    .Y(_04788_),
    .A1(net727),
    .A2(_04784_));
 sg13g2_buf_8 _21236_ (.A(net724),
    .X(_04789_));
 sg13g2_mux2_1 _21237_ (.A0(_04778_),
    .A1(_04788_),
    .S(net705),
    .X(_04790_));
 sg13g2_nand2_1 _21238_ (.Y(_04791_),
    .A(net681),
    .B(_04790_));
 sg13g2_buf_8 _21239_ (.A(net724),
    .X(_04792_));
 sg13g2_or2_1 _21240_ (.X(_04793_),
    .B(_09501_),
    .A(_09499_));
 sg13g2_nor3_1 _21241_ (.A(net984),
    .B(_09089_),
    .C(net823),
    .Y(_04794_));
 sg13g2_nor3_1 _21242_ (.A(_09089_),
    .B(_04712_),
    .C(_04751_),
    .Y(_04795_));
 sg13g2_a22oi_1 _21243_ (.Y(_04796_),
    .B1(_04795_),
    .B2(_08222_),
    .A2(_04794_),
    .A1(_04793_));
 sg13g2_buf_2 _21244_ (.A(_04796_),
    .X(_04797_));
 sg13g2_nand2b_1 _21245_ (.Y(_04798_),
    .B(_04707_),
    .A_N(_04771_));
 sg13g2_buf_2 _21246_ (.A(_04798_),
    .X(_04799_));
 sg13g2_and3_1 _21247_ (.X(_04800_),
    .A(_04727_),
    .B(_04699_),
    .C(_04735_));
 sg13g2_buf_1 _21248_ (.A(_04800_),
    .X(_04801_));
 sg13g2_or2_1 _21249_ (.X(_04802_),
    .B(_04706_),
    .A(_04727_));
 sg13g2_a22oi_1 _21250_ (.Y(_04803_),
    .B1(_04726_),
    .B2(_04802_),
    .A2(_04706_),
    .A1(_00099_));
 sg13g2_o21ai_1 _21251_ (.B1(_04782_),
    .Y(_04804_),
    .A1(_04801_),
    .A2(_04803_));
 sg13g2_mux2_1 _21252_ (.A0(_04799_),
    .A1(_04804_),
    .S(net723),
    .X(_04805_));
 sg13g2_o21ai_1 _21253_ (.B1(_04805_),
    .Y(_04806_),
    .A1(net706),
    .A2(_04797_));
 sg13g2_nand2_1 _21254_ (.Y(_04807_),
    .A(net704),
    .B(_04806_));
 sg13g2_and3_1 _21255_ (.X(_04808_),
    .A(_04775_),
    .B(_04791_),
    .C(_04807_));
 sg13g2_buf_1 _21256_ (.A(_04808_),
    .X(_04809_));
 sg13g2_buf_8 _21257_ (.A(_04809_),
    .X(_04810_));
 sg13g2_buf_8 _21258_ (.A(_04810_),
    .X(_04811_));
 sg13g2_buf_8 _21259_ (.A(net726),
    .X(_04812_));
 sg13g2_buf_8 _21260_ (.A(net728),
    .X(_04813_));
 sg13g2_buf_1 _21261_ (.A(net723),
    .X(_04814_));
 sg13g2_nor4_1 _21262_ (.A(net703),
    .B(net702),
    .C(net701),
    .D(_04784_),
    .Y(_04815_));
 sg13g2_buf_2 _21263_ (.A(_04815_),
    .X(_04816_));
 sg13g2_buf_1 _21264_ (.A(_04816_),
    .X(_04817_));
 sg13g2_buf_8 _21265_ (.A(net727),
    .X(_04818_));
 sg13g2_nor4_1 _21266_ (.A(net726),
    .B(net702),
    .C(net700),
    .D(_04784_),
    .Y(_04819_));
 sg13g2_buf_1 _21267_ (.A(_04819_),
    .X(_04820_));
 sg13g2_buf_1 _21268_ (.A(_04820_),
    .X(_04821_));
 sg13g2_a22oi_1 _21269_ (.Y(_04822_),
    .B1(net618),
    .B2(\top_ihp.oisc.regs[17][0] ),
    .A2(_04817_),
    .A1(\top_ihp.oisc.regs[25][0] ));
 sg13g2_or2_1 _21270_ (.X(_04823_),
    .B(net765),
    .A(_04716_));
 sg13g2_buf_1 _21271_ (.A(_04823_),
    .X(_04824_));
 sg13g2_nor3_1 _21272_ (.A(net704),
    .B(net681),
    .C(_04824_),
    .Y(_04825_));
 sg13g2_buf_2 _21273_ (.A(_04825_),
    .X(_04826_));
 sg13g2_buf_8 _21274_ (.A(_04826_),
    .X(_04827_));
 sg13g2_buf_8 _21275_ (.A(net726),
    .X(_04828_));
 sg13g2_buf_2 _21276_ (.A(net723),
    .X(_04829_));
 sg13g2_nand4_1 _21277_ (.B(_04706_),
    .C(_04768_),
    .A(_04701_),
    .Y(_04830_),
    .D(_04801_));
 sg13g2_nand2b_1 _21278_ (.Y(_04831_),
    .B(_08222_),
    .A_N(_04830_));
 sg13g2_buf_1 _21279_ (.A(_04831_),
    .X(_04832_));
 sg13g2_nor3_2 _21280_ (.A(net699),
    .B(net698),
    .C(_04832_),
    .Y(_04833_));
 sg13g2_buf_2 _21281_ (.A(_04833_),
    .X(_04834_));
 sg13g2_a22oi_1 _21282_ (.Y(_04835_),
    .B1(_04834_),
    .B2(\top_ihp.oisc.regs[24][0] ),
    .A2(_04827_),
    .A1(\top_ihp.oisc.regs[14][0] ));
 sg13g2_and2_1 _21283_ (.A(_04822_),
    .B(_04835_),
    .X(_04836_));
 sg13g2_buf_1 _21284_ (.A(net724),
    .X(_04837_));
 sg13g2_a22oi_1 _21285_ (.Y(_04838_),
    .B1(_04794_),
    .B2(_08210_),
    .A2(_04730_),
    .A1(_08221_));
 sg13g2_buf_2 _21286_ (.A(_04838_),
    .X(_04839_));
 sg13g2_nand2b_1 _21287_ (.Y(_04840_),
    .B(_04839_),
    .A_N(_04797_));
 sg13g2_buf_2 _21288_ (.A(_04840_),
    .X(_04841_));
 sg13g2_nor4_1 _21289_ (.A(net697),
    .B(_04776_),
    .C(net701),
    .D(_04841_),
    .Y(_04842_));
 sg13g2_buf_2 _21290_ (.A(_04842_),
    .X(_04843_));
 sg13g2_buf_8 _21291_ (.A(_04843_),
    .X(_04844_));
 sg13g2_nor4_1 _21292_ (.A(_04789_),
    .B(net706),
    .C(net700),
    .D(_04787_),
    .Y(_04845_));
 sg13g2_buf_1 _21293_ (.A(_04845_),
    .X(_04846_));
 sg13g2_buf_1 _21294_ (.A(net657),
    .X(_04847_));
 sg13g2_nand2_1 _21295_ (.Y(_04848_),
    .A(_07475_),
    .B(net803));
 sg13g2_nor2_1 _21296_ (.A(net997),
    .B(_04716_),
    .Y(_04849_));
 sg13g2_a21oi_1 _21297_ (.A1(net1017),
    .A2(net845),
    .Y(_04850_),
    .B1(_04830_));
 sg13g2_buf_2 _21298_ (.A(_04850_),
    .X(_04851_));
 sg13g2_nor2b_1 _21299_ (.A(_04849_),
    .B_N(net797),
    .Y(_04852_));
 sg13g2_buf_2 _21300_ (.A(_04852_),
    .X(_04853_));
 sg13g2_and2_1 _21301_ (.A(net699),
    .B(net722),
    .X(_04854_));
 sg13g2_buf_1 _21302_ (.A(_04854_),
    .X(_04855_));
 sg13g2_nand2_1 _21303_ (.Y(_04856_),
    .A(\top_ihp.oisc.regs[20][0] ),
    .B(_04855_));
 sg13g2_nand2_1 _21304_ (.Y(_04857_),
    .A(_04848_),
    .B(_04856_));
 sg13g2_a221oi_1 _21305_ (.B2(\top_ihp.oisc.regs[7][0] ),
    .C1(_04857_),
    .B1(net617),
    .A1(\top_ihp.oisc.regs[47][0] ),
    .Y(_04858_),
    .A2(net476));
 sg13g2_a221oi_1 _21306_ (.B2(_09072_),
    .C1(_04736_),
    .B1(_08230_),
    .A1(net1017),
    .Y(_04859_),
    .A2(_08220_));
 sg13g2_o21ai_1 _21307_ (.B1(_04723_),
    .Y(_04860_),
    .A1(_04691_),
    .A2(_04859_));
 sg13g2_buf_2 _21308_ (.A(_04860_),
    .X(_04861_));
 sg13g2_nor3_2 _21309_ (.A(net728),
    .B(net727),
    .C(_04861_),
    .Y(_04862_));
 sg13g2_nor2_1 _21310_ (.A(net724),
    .B(_04733_),
    .Y(_04863_));
 sg13g2_and2_1 _21311_ (.A(_04862_),
    .B(_04863_),
    .X(_04864_));
 sg13g2_buf_2 _21312_ (.A(_04864_),
    .X(_04865_));
 sg13g2_buf_8 _21313_ (.A(_04865_),
    .X(_04866_));
 sg13g2_nor3_2 _21314_ (.A(_04748_),
    .B(net727),
    .C(_04861_),
    .Y(_04867_));
 sg13g2_and2_1 _21315_ (.A(_04863_),
    .B(_04867_),
    .X(_04868_));
 sg13g2_buf_2 _21316_ (.A(_04868_),
    .X(_04869_));
 sg13g2_buf_8 _21317_ (.A(_04869_),
    .X(_04870_));
 sg13g2_buf_8 _21318_ (.A(net615),
    .X(_04871_));
 sg13g2_a22oi_1 _21319_ (.Y(_04872_),
    .B1(net475),
    .B2(\top_ihp.oisc.regs[55][0] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][0] ));
 sg13g2_buf_8 _21320_ (.A(_04818_),
    .X(_04873_));
 sg13g2_nor4_1 _21321_ (.A(_04812_),
    .B(_04813_),
    .C(net680),
    .D(_04841_),
    .Y(_04874_));
 sg13g2_buf_2 _21322_ (.A(_04874_),
    .X(_04875_));
 sg13g2_buf_1 _21323_ (.A(_04875_),
    .X(_04876_));
 sg13g2_buf_1 _21324_ (.A(net681),
    .X(_04877_));
 sg13g2_buf_1 _21325_ (.A(_04784_),
    .X(_04878_));
 sg13g2_nor2_1 _21326_ (.A(_04812_),
    .B(_04814_),
    .Y(_04879_));
 sg13g2_buf_2 _21327_ (.A(_04879_),
    .X(_04880_));
 sg13g2_nor2_1 _21328_ (.A(_04789_),
    .B(net700),
    .Y(_04881_));
 sg13g2_buf_2 _21329_ (.A(_04881_),
    .X(_04882_));
 sg13g2_a22oi_1 _21330_ (.Y(_04883_),
    .B1(_04882_),
    .B2(\top_ihp.oisc.regs[23][0] ),
    .A2(_04880_),
    .A1(\top_ihp.oisc.regs[27][0] ));
 sg13g2_nor3_1 _21331_ (.A(_04877_),
    .B(net696),
    .C(_04883_),
    .Y(_04884_));
 sg13g2_a21oi_1 _21332_ (.A1(\top_ihp.oisc.regs[33][0] ),
    .A2(net474),
    .Y(_04885_),
    .B1(_04884_));
 sg13g2_nand4_1 _21333_ (.B(_04858_),
    .C(_04872_),
    .A(_04836_),
    .Y(_04886_),
    .D(_04885_));
 sg13g2_nor4_1 _21334_ (.A(net705),
    .B(net702),
    .C(net701),
    .D(_04787_),
    .Y(_04887_));
 sg13g2_buf_1 _21335_ (.A(_04887_),
    .X(_04888_));
 sg13g2_buf_2 _21336_ (.A(net655),
    .X(_04889_));
 sg13g2_buf_8 _21337_ (.A(_04889_),
    .X(_04890_));
 sg13g2_nor4_1 _21338_ (.A(net705),
    .B(net702),
    .C(net701),
    .D(net696),
    .Y(_04891_));
 sg13g2_buf_1 _21339_ (.A(_04891_),
    .X(_04892_));
 sg13g2_buf_1 _21340_ (.A(_04892_),
    .X(_04893_));
 sg13g2_buf_1 _21341_ (.A(net613),
    .X(_04894_));
 sg13g2_a22oi_1 _21342_ (.Y(_04895_),
    .B1(net472),
    .B2(\top_ihp.oisc.regs[29][0] ),
    .A2(net473),
    .A1(\top_ihp.oisc.regs[13][0] ));
 sg13g2_buf_1 _21343_ (.A(_04824_),
    .X(_04896_));
 sg13g2_nor3_1 _21344_ (.A(_04828_),
    .B(net681),
    .C(net679),
    .Y(_04897_));
 sg13g2_buf_2 _21345_ (.A(_04897_),
    .X(_04898_));
 sg13g2_buf_1 _21346_ (.A(_04898_),
    .X(_04899_));
 sg13g2_nor4_1 _21347_ (.A(net705),
    .B(net702),
    .C(net700),
    .D(net696),
    .Y(_04900_));
 sg13g2_buf_2 _21348_ (.A(_04900_),
    .X(_04901_));
 sg13g2_buf_8 _21349_ (.A(_04901_),
    .X(_04902_));
 sg13g2_buf_2 _21350_ (.A(net612),
    .X(_04903_));
 sg13g2_a22oi_1 _21351_ (.Y(_04904_),
    .B1(net470),
    .B2(\top_ihp.oisc.regs[21][0] ),
    .A2(net471),
    .A1(\top_ihp.oisc.regs[10][0] ));
 sg13g2_nor3_2 _21352_ (.A(net724),
    .B(net728),
    .C(_04787_),
    .Y(_04905_));
 sg13g2_and2_1 _21353_ (.A(net698),
    .B(_04905_),
    .X(_04906_));
 sg13g2_buf_1 _21354_ (.A(_04906_),
    .X(_04907_));
 sg13g2_buf_8 _21355_ (.A(_04907_),
    .X(_04908_));
 sg13g2_buf_8 _21356_ (.A(net611),
    .X(_04909_));
 sg13g2_buf_2 _21357_ (.A(net704),
    .X(_04910_));
 sg13g2_buf_1 _21358_ (.A(net678),
    .X(_04911_));
 sg13g2_mux2_1 _21359_ (.A0(\top_ihp.oisc.regs[22][0] ),
    .A1(\top_ihp.oisc.regs[18][0] ),
    .S(net654),
    .X(_04912_));
 sg13g2_nand2_1 _21360_ (.Y(_04913_),
    .A(_04702_),
    .B(_04701_));
 sg13g2_and2_1 _21361_ (.A(_04801_),
    .B(_04913_),
    .X(_04914_));
 sg13g2_and3_1 _21362_ (.X(_04915_),
    .A(_04716_),
    .B(_04782_),
    .C(_04914_));
 sg13g2_buf_1 _21363_ (.A(_04915_),
    .X(_04916_));
 sg13g2_buf_2 _21364_ (.A(net721),
    .X(_04917_));
 sg13g2_a22oi_1 _21365_ (.Y(_04918_),
    .B1(_04912_),
    .B2(net695),
    .A2(net469),
    .A1(\top_ihp.oisc.regs[5][0] ));
 sg13g2_nor4_1 _21366_ (.A(net697),
    .B(net681),
    .C(net680),
    .D(net765),
    .Y(_04919_));
 sg13g2_buf_1 _21367_ (.A(_04919_),
    .X(_04920_));
 sg13g2_buf_1 _21368_ (.A(net610),
    .X(_04921_));
 sg13g2_nand2_1 _21369_ (.Y(_04922_),
    .A(\top_ihp.oisc.regs[6][0] ),
    .B(net468));
 sg13g2_nand4_1 _21370_ (.B(_04904_),
    .C(_04918_),
    .A(_04895_),
    .Y(_04923_),
    .D(_04922_));
 sg13g2_nor4_1 _21371_ (.A(net705),
    .B(net706),
    .C(net701),
    .D(_04787_),
    .Y(_04924_));
 sg13g2_buf_1 _21372_ (.A(_04924_),
    .X(_04925_));
 sg13g2_buf_8 _21373_ (.A(net653),
    .X(_04926_));
 sg13g2_buf_1 _21374_ (.A(net609),
    .X(_04927_));
 sg13g2_nand2_1 _21375_ (.Y(_04928_),
    .A(_04801_),
    .B(_04913_));
 sg13g2_nor4_2 _21376_ (.A(_03696_),
    .B(_04716_),
    .C(_04780_),
    .Y(_04929_),
    .D(_04928_));
 sg13g2_buf_2 _21377_ (.A(_04929_),
    .X(_04930_));
 sg13g2_buf_1 _21378_ (.A(net678),
    .X(_04931_));
 sg13g2_mux2_1 _21379_ (.A0(\top_ihp.oisc.regs[30][0] ),
    .A1(\top_ihp.oisc.regs[26][0] ),
    .S(net652),
    .X(_04932_));
 sg13g2_a22oi_1 _21380_ (.Y(_04933_),
    .B1(net720),
    .B2(_04932_),
    .A2(_04927_),
    .A1(\top_ihp.oisc.regs[15][0] ));
 sg13g2_nor4_1 _21381_ (.A(net703),
    .B(net702),
    .C(net700),
    .D(_04787_),
    .Y(_04934_));
 sg13g2_buf_1 _21382_ (.A(_04934_),
    .X(_04935_));
 sg13g2_buf_1 _21383_ (.A(_04935_),
    .X(_04936_));
 sg13g2_buf_1 _21384_ (.A(net608),
    .X(_04937_));
 sg13g2_nor4_1 _21385_ (.A(net705),
    .B(net706),
    .C(net701),
    .D(net696),
    .Y(_04938_));
 sg13g2_buf_2 _21386_ (.A(_04938_),
    .X(_04939_));
 sg13g2_buf_8 _21387_ (.A(_04939_),
    .X(_04940_));
 sg13g2_buf_1 _21388_ (.A(net607),
    .X(_04941_));
 sg13g2_a22oi_1 _21389_ (.Y(_04942_),
    .B1(net465),
    .B2(\top_ihp.oisc.regs[31][0] ),
    .A2(net466),
    .A1(\top_ihp.oisc.regs[1][0] ));
 sg13g2_buf_1 _21390_ (.A(_04710_),
    .X(_04943_));
 sg13g2_buf_1 _21391_ (.A(_04943_),
    .X(_04944_));
 sg13g2_nor2_2 _21392_ (.A(net677),
    .B(net679),
    .Y(_04945_));
 sg13g2_mux2_1 _21393_ (.A0(\top_ihp.oisc.regs[12][0] ),
    .A1(\top_ihp.oisc.regs[8][0] ),
    .S(net654),
    .X(_04946_));
 sg13g2_nand2_2 _21394_ (.Y(_04947_),
    .A(net699),
    .B(net680));
 sg13g2_nor2_2 _21395_ (.A(_04832_),
    .B(_04947_),
    .Y(_04948_));
 sg13g2_buf_8 _21396_ (.A(_04948_),
    .X(_04949_));
 sg13g2_a22oi_1 _21397_ (.Y(_04950_),
    .B1(net464),
    .B2(\top_ihp.oisc.regs[28][0] ),
    .A2(_04946_),
    .A1(_04945_));
 sg13g2_nor3_1 _21398_ (.A(_04828_),
    .B(net680),
    .C(_04832_),
    .Y(_04951_));
 sg13g2_buf_2 _21399_ (.A(net725),
    .X(_04952_));
 sg13g2_buf_2 _21400_ (.A(net693),
    .X(_04953_));
 sg13g2_mux2_1 _21401_ (.A0(\top_ihp.oisc.regs[3][0] ),
    .A1(\top_ihp.oisc.regs[19][0] ),
    .S(net676),
    .X(_04954_));
 sg13g2_a22oi_1 _21402_ (.Y(_04955_),
    .B1(_04713_),
    .B2(_04739_),
    .A2(_04712_),
    .A1(\top_ihp.oisc.micro_op[14] ));
 sg13g2_and4_1 _21403_ (.A(_04955_),
    .B(_04716_),
    .C(_04782_),
    .D(_04803_),
    .X(_04956_));
 sg13g2_buf_2 _21404_ (.A(_04956_),
    .X(_04957_));
 sg13g2_buf_2 _21405_ (.A(_04957_),
    .X(_04958_));
 sg13g2_buf_1 _21406_ (.A(net692),
    .X(_04959_));
 sg13g2_a22oi_1 _21407_ (.Y(_04960_),
    .B1(_04954_),
    .B2(net675),
    .A2(_04951_),
    .A1(\top_ihp.oisc.regs[16][0] ));
 sg13g2_nand4_1 _21408_ (.B(_04942_),
    .C(_04950_),
    .A(_04933_),
    .Y(_04961_),
    .D(_04960_));
 sg13g2_nor4_1 _21409_ (.A(net80),
    .B(_04886_),
    .C(_04923_),
    .D(_04961_),
    .Y(_04962_));
 sg13g2_nor3_1 _21410_ (.A(net726),
    .B(_04839_),
    .C(_04797_),
    .Y(_04963_));
 sg13g2_and2_1 _21411_ (.A(_04722_),
    .B(_04963_),
    .X(_04964_));
 sg13g2_buf_2 _21412_ (.A(_04964_),
    .X(_04965_));
 sg13g2_buf_2 _21413_ (.A(_04965_),
    .X(_04966_));
 sg13g2_nor2_1 _21414_ (.A(_04759_),
    .B(_04839_),
    .Y(_04967_));
 sg13g2_and2_1 _21415_ (.A(_04867_),
    .B(_04967_),
    .X(_04968_));
 sg13g2_buf_2 _21416_ (.A(_04968_),
    .X(_04969_));
 sg13g2_buf_1 _21417_ (.A(_04969_),
    .X(_04970_));
 sg13g2_a22oi_1 _21418_ (.Y(_04971_),
    .B1(net606),
    .B2(\top_ihp.oisc.regs[54][0] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][0] ));
 sg13g2_nor2_2 _21419_ (.A(_04748_),
    .B(net723),
    .Y(_04972_));
 sg13g2_and2_1 _21420_ (.A(_04972_),
    .B(_04963_),
    .X(_04973_));
 sg13g2_buf_2 _21421_ (.A(_04973_),
    .X(_04974_));
 sg13g2_buf_8 _21422_ (.A(_04974_),
    .X(_04975_));
 sg13g2_nor2_1 _21423_ (.A(net726),
    .B(_04733_),
    .Y(_04976_));
 sg13g2_and2_1 _21424_ (.A(_04862_),
    .B(_04976_),
    .X(_04977_));
 sg13g2_buf_2 _21425_ (.A(_04977_),
    .X(_04978_));
 sg13g2_buf_2 _21426_ (.A(_04978_),
    .X(_04979_));
 sg13g2_a22oi_1 _21427_ (.Y(_04980_),
    .B1(net604),
    .B2(\top_ihp.oisc.regs[49][0] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][0] ));
 sg13g2_nor3_1 _21428_ (.A(net726),
    .B(net723),
    .C(_04861_),
    .Y(_04981_));
 sg13g2_and3_1 _21429_ (.X(_04982_),
    .A(_04943_),
    .B(_04733_),
    .C(_04981_));
 sg13g2_buf_2 _21430_ (.A(_04982_),
    .X(_04983_));
 sg13g2_buf_8 _21431_ (.A(_04983_),
    .X(_04984_));
 sg13g2_or2_1 _21432_ (.X(_04985_),
    .B(_04797_),
    .A(_04839_));
 sg13g2_buf_1 _21433_ (.A(_04985_),
    .X(_04986_));
 sg13g2_nor4_1 _21434_ (.A(net697),
    .B(net694),
    .C(net680),
    .D(_04986_),
    .Y(_04987_));
 sg13g2_buf_2 _21435_ (.A(_04987_),
    .X(_04988_));
 sg13g2_buf_8 _21436_ (.A(_04988_),
    .X(_04989_));
 sg13g2_a22oi_1 _21437_ (.Y(_04990_),
    .B1(net462),
    .B2(\top_ihp.oisc.regs[36][0] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[58][0] ));
 sg13g2_nor3_1 _21438_ (.A(_04759_),
    .B(_04748_),
    .C(net727),
    .Y(_04991_));
 sg13g2_buf_1 _21439_ (.A(_04991_),
    .X(_04992_));
 sg13g2_nor2b_1 _21440_ (.A(_04986_),
    .B_N(_04992_),
    .Y(_04993_));
 sg13g2_buf_2 _21441_ (.A(_04993_),
    .X(_04994_));
 sg13g2_buf_8 _21442_ (.A(_04994_),
    .X(_04995_));
 sg13g2_nor3_1 _21443_ (.A(_04748_),
    .B(net723),
    .C(_04861_),
    .Y(_04996_));
 sg13g2_and2_1 _21444_ (.A(_04976_),
    .B(_04996_),
    .X(_04997_));
 sg13g2_buf_2 _21445_ (.A(_04997_),
    .X(_04998_));
 sg13g2_buf_8 _21446_ (.A(_04998_),
    .X(_04999_));
 sg13g2_a22oi_1 _21447_ (.Y(_05000_),
    .B1(net602),
    .B2(\top_ihp.oisc.regs[59][0] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][0] ));
 sg13g2_nand4_1 _21448_ (.B(_04980_),
    .C(_04990_),
    .A(_04971_),
    .Y(_05001_),
    .D(_05000_));
 sg13g2_and3_1 _21449_ (.X(_05002_),
    .A(net704),
    .B(_04733_),
    .C(_04862_));
 sg13g2_buf_1 _21450_ (.A(_05002_),
    .X(_05003_));
 sg13g2_buf_1 _21451_ (.A(_05003_),
    .X(_05004_));
 sg13g2_nand2_1 _21452_ (.Y(_05005_),
    .A(\top_ihp.oisc.regs[48][0] ),
    .B(net601));
 sg13g2_nor3_1 _21453_ (.A(_04744_),
    .B(_04748_),
    .C(_04720_),
    .Y(_05006_));
 sg13g2_buf_2 _21454_ (.A(_05006_),
    .X(_05007_));
 sg13g2_nor2b_1 _21455_ (.A(net765),
    .B_N(_05007_),
    .Y(_05008_));
 sg13g2_buf_1 _21456_ (.A(_05008_),
    .X(_05009_));
 sg13g2_and2_1 _21457_ (.A(_04867_),
    .B(_04976_),
    .X(_05010_));
 sg13g2_buf_2 _21458_ (.A(_05010_),
    .X(_05011_));
 sg13g2_buf_2 _21459_ (.A(_05011_),
    .X(_05012_));
 sg13g2_a22oi_1 _21460_ (.Y(_05013_),
    .B1(net599),
    .B2(\top_ihp.oisc.regs[51][0] ),
    .A2(net600),
    .A1(\top_ihp.oisc.regs[2][0] ));
 sg13g2_nor4_1 _21461_ (.A(net705),
    .B(net702),
    .C(net700),
    .D(net765),
    .Y(_05014_));
 sg13g2_buf_2 _21462_ (.A(_05014_),
    .X(_05015_));
 sg13g2_buf_1 _21463_ (.A(_05015_),
    .X(_05016_));
 sg13g2_buf_1 _21464_ (.A(_04787_),
    .X(_05017_));
 sg13g2_nor4_1 _21465_ (.A(net703),
    .B(net706),
    .C(net698),
    .D(net691),
    .Y(_05018_));
 sg13g2_buf_1 _21466_ (.A(_05018_),
    .X(_05019_));
 sg13g2_nor4_1 _21467_ (.A(net703),
    .B(net702),
    .C(net701),
    .D(_04787_),
    .Y(_05020_));
 sg13g2_buf_1 _21468_ (.A(_05020_),
    .X(_05021_));
 sg13g2_buf_1 _21469_ (.A(_05021_),
    .X(_05022_));
 sg13g2_and2_1 _21470_ (.A(\top_ihp.oisc.regs[9][0] ),
    .B(net597),
    .X(_05023_));
 sg13g2_a221oi_1 _21471_ (.B2(\top_ihp.oisc.regs[11][0] ),
    .C1(_05023_),
    .B1(net651),
    .A1(\top_ihp.oisc.regs[4][0] ),
    .Y(_05024_),
    .A2(net598));
 sg13g2_nand2_1 _21472_ (.Y(_05025_),
    .A(net724),
    .B(net728));
 sg13g2_nor3_1 _21473_ (.A(_05025_),
    .B(net698),
    .C(_04841_),
    .Y(_05026_));
 sg13g2_buf_2 _21474_ (.A(_05026_),
    .X(_05027_));
 sg13g2_buf_8 _21475_ (.A(_05027_),
    .X(_05028_));
 sg13g2_and2_1 _21476_ (.A(_04863_),
    .B(_04996_),
    .X(_05029_));
 sg13g2_buf_8 _21477_ (.A(_05029_),
    .X(_05030_));
 sg13g2_buf_8 _21478_ (.A(_05030_),
    .X(_05031_));
 sg13g2_a22oi_1 _21479_ (.Y(_05032_),
    .B1(net596),
    .B2(\top_ihp.oisc.regs[63][0] ),
    .A2(net460),
    .A1(\top_ihp.oisc.regs[43][0] ));
 sg13g2_nand4_1 _21480_ (.B(_05013_),
    .C(_05024_),
    .A(_05005_),
    .Y(_05033_),
    .D(_05032_));
 sg13g2_and3_1 _21481_ (.X(_05034_),
    .A(_04777_),
    .B(_04733_),
    .C(_04981_));
 sg13g2_buf_2 _21482_ (.A(_05034_),
    .X(_05035_));
 sg13g2_buf_8 _21483_ (.A(_05035_),
    .X(_05036_));
 sg13g2_buf_8 _21484_ (.A(net459),
    .X(_05037_));
 sg13g2_and3_1 _21485_ (.X(_05038_),
    .A(_04792_),
    .B(_04733_),
    .C(_04867_));
 sg13g2_buf_2 _21486_ (.A(_05038_),
    .X(_05039_));
 sg13g2_buf_2 _21487_ (.A(_05039_),
    .X(_05040_));
 sg13g2_a22oi_1 _21488_ (.Y(_05041_),
    .B1(net595),
    .B2(\top_ihp.oisc.regs[50][0] ),
    .A2(net273),
    .A1(\top_ihp.oisc.regs[56][0] ));
 sg13g2_nor4_1 _21489_ (.A(net697),
    .B(_04813_),
    .C(_04814_),
    .D(_04986_),
    .Y(_05042_));
 sg13g2_buf_2 _21490_ (.A(_05042_),
    .X(_05043_));
 sg13g2_buf_8 _21491_ (.A(_05043_),
    .X(_05044_));
 sg13g2_and2_1 _21492_ (.A(_04967_),
    .B(_04996_),
    .X(_05045_));
 sg13g2_buf_1 _21493_ (.A(_05045_),
    .X(_05046_));
 sg13g2_buf_2 _21494_ (.A(_05046_),
    .X(_05047_));
 sg13g2_a22oi_1 _21495_ (.Y(_05048_),
    .B1(net594),
    .B2(\top_ihp.oisc.regs[62][0] ),
    .A2(net458),
    .A1(\top_ihp.oisc.regs[44][0] ));
 sg13g2_nor3_1 _21496_ (.A(net728),
    .B(net723),
    .C(_04861_),
    .Y(_05049_));
 sg13g2_and2_1 _21497_ (.A(_04863_),
    .B(_05049_),
    .X(_05050_));
 sg13g2_buf_8 _21498_ (.A(_05050_),
    .X(_05051_));
 sg13g2_buf_8 _21499_ (.A(_05051_),
    .X(_05052_));
 sg13g2_nor3_1 _21500_ (.A(_05025_),
    .B(_04873_),
    .C(_04841_),
    .Y(_05053_));
 sg13g2_buf_2 _21501_ (.A(_05053_),
    .X(_05054_));
 sg13g2_buf_2 _21502_ (.A(_05054_),
    .X(_05055_));
 sg13g2_a22oi_1 _21503_ (.Y(_05056_),
    .B1(net457),
    .B2(\top_ihp.oisc.regs[35][0] ),
    .A2(net593),
    .A1(\top_ihp.oisc.regs[61][0] ));
 sg13g2_nor4_1 _21504_ (.A(net697),
    .B(_04777_),
    .C(net698),
    .D(_04986_),
    .Y(_05057_));
 sg13g2_buf_2 _21505_ (.A(_05057_),
    .X(_05058_));
 sg13g2_buf_8 _21506_ (.A(_05058_),
    .X(_05059_));
 sg13g2_and2_1 _21507_ (.A(_04976_),
    .B(_05049_),
    .X(_05060_));
 sg13g2_buf_8 _21508_ (.A(_05060_),
    .X(_05061_));
 sg13g2_buf_1 _21509_ (.A(_05061_),
    .X(_05062_));
 sg13g2_a22oi_1 _21510_ (.Y(_05063_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][0] ),
    .A2(net456),
    .A1(\top_ihp.oisc.regs[46][0] ));
 sg13g2_nand4_1 _21511_ (.B(_05048_),
    .C(_05056_),
    .A(_05041_),
    .Y(_05064_),
    .D(_05063_));
 sg13g2_and2_1 _21512_ (.A(_04862_),
    .B(_04967_),
    .X(_05065_));
 sg13g2_buf_2 _21513_ (.A(_05065_),
    .X(_05066_));
 sg13g2_buf_8 _21514_ (.A(_05066_),
    .X(_05067_));
 sg13g2_buf_1 _21515_ (.A(net591),
    .X(_05068_));
 sg13g2_nor2_1 _21516_ (.A(_04776_),
    .B(net700),
    .Y(_05069_));
 sg13g2_and2_1 _21517_ (.A(_05069_),
    .B(_04963_),
    .X(_05070_));
 sg13g2_buf_2 _21518_ (.A(_05070_),
    .X(_05071_));
 sg13g2_buf_8 _21519_ (.A(_05071_),
    .X(_05072_));
 sg13g2_buf_8 _21520_ (.A(net454),
    .X(_05073_));
 sg13g2_a22oi_1 _21521_ (.Y(_05074_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][0] ),
    .A2(net455),
    .A1(\top_ihp.oisc.regs[52][0] ));
 sg13g2_nor4_1 _21522_ (.A(_04837_),
    .B(net694),
    .C(net698),
    .D(_04841_),
    .Y(_05075_));
 sg13g2_buf_2 _21523_ (.A(_05075_),
    .X(_05076_));
 sg13g2_buf_2 _21524_ (.A(_05076_),
    .X(_05077_));
 sg13g2_nor2b_1 _21525_ (.A(_04841_),
    .B_N(_04992_),
    .Y(_05078_));
 sg13g2_buf_2 _21526_ (.A(_05078_),
    .X(_05079_));
 sg13g2_buf_1 _21527_ (.A(_05079_),
    .X(_05080_));
 sg13g2_a22oi_1 _21528_ (.Y(_05081_),
    .B1(net452),
    .B2(\top_ihp.oisc.regs[39][0] ),
    .A2(net453),
    .A1(\top_ihp.oisc.regs[45][0] ));
 sg13g2_nor3_1 _21529_ (.A(_04744_),
    .B(_04710_),
    .C(_04767_),
    .Y(_05082_));
 sg13g2_buf_1 _21530_ (.A(_05082_),
    .X(_05083_));
 sg13g2_nor2b_1 _21531_ (.A(_04986_),
    .B_N(net673),
    .Y(_05084_));
 sg13g2_buf_2 _21532_ (.A(_05084_),
    .X(_05085_));
 sg13g2_buf_8 _21533_ (.A(_05085_),
    .X(_05086_));
 sg13g2_nor4_1 _21534_ (.A(_04837_),
    .B(net694),
    .C(net680),
    .D(_04841_),
    .Y(_05087_));
 sg13g2_buf_2 _21535_ (.A(_05087_),
    .X(_05088_));
 sg13g2_buf_8 _21536_ (.A(_05088_),
    .X(_05089_));
 sg13g2_buf_8 _21537_ (.A(net450),
    .X(_05090_));
 sg13g2_a22oi_1 _21538_ (.Y(_05091_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][0] ),
    .A2(net451),
    .A1(\top_ihp.oisc.regs[40][0] ));
 sg13g2_nor2b_1 _21539_ (.A(_04841_),
    .B_N(net673),
    .Y(_05092_));
 sg13g2_buf_2 _21540_ (.A(_05092_),
    .X(_05093_));
 sg13g2_buf_8 _21541_ (.A(_05093_),
    .X(_05094_));
 sg13g2_and2_1 _21542_ (.A(_04967_),
    .B(_05049_),
    .X(_05095_));
 sg13g2_buf_2 _21543_ (.A(_05095_),
    .X(_05096_));
 sg13g2_buf_1 _21544_ (.A(_05096_),
    .X(_05097_));
 sg13g2_a22oi_1 _21545_ (.Y(_05098_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][0] ),
    .A2(net449),
    .A1(\top_ihp.oisc.regs[41][0] ));
 sg13g2_nand4_1 _21546_ (.B(_05081_),
    .C(_05091_),
    .A(_05074_),
    .Y(_05099_),
    .D(_05098_));
 sg13g2_nor4_2 _21547_ (.A(_05001_),
    .B(_05033_),
    .C(_05064_),
    .Y(_05100_),
    .D(_05099_));
 sg13g2_buf_8 _21548_ (.A(_04810_),
    .X(_05101_));
 sg13g2_a21oi_1 _21549_ (.A1(_04751_),
    .A2(_04782_),
    .Y(_05102_),
    .B1(net803));
 sg13g2_nand2b_1 _21550_ (.Y(_05103_),
    .B(_05102_),
    .A_N(_04965_));
 sg13g2_buf_2 _21551_ (.A(_05103_),
    .X(_05104_));
 sg13g2_buf_8 _21552_ (.A(_05104_),
    .X(_05105_));
 sg13g2_a21o_1 _21553_ (.A2(net79),
    .A1(_09053_),
    .B1(net154),
    .X(_05106_));
 sg13g2_a22oi_1 _21554_ (.Y(_00294_),
    .B1(_05106_),
    .B2(_04848_),
    .A2(_05100_),
    .A1(_04962_));
 sg13g2_buf_8 _21555_ (.A(net456),
    .X(_05107_));
 sg13g2_a22oi_1 _21556_ (.Y(_05108_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][10] ),
    .A2(net270),
    .A1(\top_ihp.oisc.regs[46][10] ));
 sg13g2_buf_1 _21557_ (.A(net615),
    .X(_05109_));
 sg13g2_buf_8 _21558_ (.A(_05028_),
    .X(_05110_));
 sg13g2_a22oi_1 _21559_ (.Y(_05111_),
    .B1(net269),
    .B2(\top_ihp.oisc.regs[43][10] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][10] ));
 sg13g2_buf_1 _21560_ (.A(_05054_),
    .X(_05112_));
 sg13g2_a22oi_1 _21561_ (.Y(_05113_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][10] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[35][10] ));
 sg13g2_buf_8 _21562_ (.A(net458),
    .X(_05114_));
 sg13g2_buf_8 _21563_ (.A(_05096_),
    .X(_05115_));
 sg13g2_buf_8 _21564_ (.A(net589),
    .X(_05116_));
 sg13g2_a22oi_1 _21565_ (.Y(_05117_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][10] ),
    .A2(net268),
    .A1(\top_ihp.oisc.regs[44][10] ));
 sg13g2_nand4_1 _21566_ (.B(_05111_),
    .C(_05113_),
    .A(_05108_),
    .Y(_05118_),
    .D(_05117_));
 sg13g2_buf_1 _21567_ (.A(net765),
    .X(_05119_));
 sg13g2_a22oi_1 _21568_ (.Y(_05120_),
    .B1(net673),
    .B2(\top_ihp.oisc.regs[8][10] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[6][10] ));
 sg13g2_mux2_1 _21569_ (.A0(\top_ihp.oisc.regs[26][10] ),
    .A1(\top_ihp.oisc.regs[18][10] ),
    .S(net698),
    .X(_05121_));
 sg13g2_buf_2 _21570_ (.A(net704),
    .X(_05122_));
 sg13g2_a22oi_1 _21571_ (.Y(_05123_),
    .B1(_05121_),
    .B2(net672),
    .A2(_04882_),
    .A1(\top_ihp.oisc.regs[22][10] ));
 sg13g2_and2_1 _21572_ (.A(_04782_),
    .B(_04914_),
    .X(_05124_));
 sg13g2_buf_1 _21573_ (.A(_05124_),
    .X(_05125_));
 sg13g2_buf_1 _21574_ (.A(_05125_),
    .X(_05126_));
 sg13g2_buf_1 _21575_ (.A(_05126_),
    .X(_05127_));
 sg13g2_nand2b_1 _21576_ (.Y(_05128_),
    .B(_05127_),
    .A_N(_05123_));
 sg13g2_o21ai_1 _21577_ (.B1(_05128_),
    .Y(_05129_),
    .A1(net719),
    .A2(_05120_));
 sg13g2_buf_2 _21578_ (.A(_04832_),
    .X(_05130_));
 sg13g2_buf_1 _21579_ (.A(_04880_),
    .X(_05131_));
 sg13g2_buf_8 _21580_ (.A(_04829_),
    .X(_05132_));
 sg13g2_mux2_1 _21581_ (.A0(\top_ihp.oisc.regs[28][10] ),
    .A1(\top_ihp.oisc.regs[20][10] ),
    .S(net670),
    .X(_05133_));
 sg13g2_buf_2 _21582_ (.A(net699),
    .X(_05134_));
 sg13g2_buf_1 _21583_ (.A(net669),
    .X(_05135_));
 sg13g2_a22oi_1 _21584_ (.Y(_05136_),
    .B1(_05133_),
    .B2(net650),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[24][10] ));
 sg13g2_nor2_1 _21585_ (.A(net689),
    .B(_05136_),
    .Y(_05137_));
 sg13g2_a22oi_1 _21586_ (.Y(_05138_),
    .B1(_04898_),
    .B2(\top_ihp.oisc.regs[10][10] ),
    .A2(net477),
    .A1(\top_ihp.oisc.regs[14][10] ));
 sg13g2_buf_2 _21587_ (.A(_04845_),
    .X(_05139_));
 sg13g2_nor4_1 _21588_ (.A(net705),
    .B(net706),
    .C(net700),
    .D(net696),
    .Y(_05140_));
 sg13g2_buf_1 _21589_ (.A(_05140_),
    .X(_05141_));
 sg13g2_buf_8 _21590_ (.A(net648),
    .X(_05142_));
 sg13g2_a22oi_1 _21591_ (.Y(_05143_),
    .B1(net587),
    .B2(\top_ihp.oisc.regs[23][10] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][10] ));
 sg13g2_buf_1 _21592_ (.A(_04820_),
    .X(_05144_));
 sg13g2_a22oi_1 _21593_ (.Y(_05145_),
    .B1(net613),
    .B2(\top_ihp.oisc.regs[29][10] ),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][10] ));
 sg13g2_buf_1 _21594_ (.A(_05018_),
    .X(_05146_));
 sg13g2_a22oi_1 _21595_ (.Y(_05147_),
    .B1(net647),
    .B2(\top_ihp.oisc.regs[11][10] ),
    .A2(net653),
    .A1(\top_ihp.oisc.regs[15][10] ));
 sg13g2_nand4_1 _21596_ (.B(_05143_),
    .C(_05145_),
    .A(_05138_),
    .Y(_05148_),
    .D(_05147_));
 sg13g2_nor3_1 _21597_ (.A(net704),
    .B(net694),
    .C(net679),
    .Y(_05149_));
 sg13g2_buf_1 _21598_ (.A(_05149_),
    .X(_05150_));
 sg13g2_nand2_1 _21599_ (.Y(_05151_),
    .A(\top_ihp.oisc.regs[12][10] ),
    .B(net585));
 sg13g2_nor4_1 _21600_ (.A(net703),
    .B(net706),
    .C(net701),
    .D(net696),
    .Y(_05152_));
 sg13g2_buf_1 _21601_ (.A(_05152_),
    .X(_05153_));
 sg13g2_buf_1 _21602_ (.A(_05153_),
    .X(_05154_));
 sg13g2_a22oi_1 _21603_ (.Y(_05155_),
    .B1(net584),
    .B2(\top_ihp.oisc.regs[27][10] ),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[5][10] ));
 sg13g2_mux2_1 _21604_ (.A0(\top_ihp.oisc.regs[3][10] ),
    .A1(\top_ihp.oisc.regs[19][10] ),
    .S(net693),
    .X(_05156_));
 sg13g2_a22oi_1 _21605_ (.Y(_05157_),
    .B1(_05156_),
    .B2(net692),
    .A2(net597),
    .A1(\top_ihp.oisc.regs[9][10] ));
 sg13g2_buf_1 _21606_ (.A(_04901_),
    .X(_05158_));
 sg13g2_a22oi_1 _21607_ (.Y(_05159_),
    .B1(net608),
    .B2(\top_ihp.oisc.regs[1][10] ),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][10] ));
 sg13g2_nand4_1 _21608_ (.B(_05155_),
    .C(_05157_),
    .A(_05151_),
    .Y(_05160_),
    .D(_05159_));
 sg13g2_or4_1 _21609_ (.A(_05129_),
    .B(_05137_),
    .C(_05148_),
    .D(_05160_),
    .X(_05161_));
 sg13g2_nor3_1 _21610_ (.A(net79),
    .B(_05118_),
    .C(_05161_),
    .Y(_05162_));
 sg13g2_a22oi_1 _21611_ (.Y(_05163_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][10] ),
    .A2(net604),
    .A1(\top_ihp.oisc.regs[49][10] ));
 sg13g2_buf_2 _21612_ (.A(_05079_),
    .X(_05164_));
 sg13g2_a22oi_1 _21613_ (.Y(_05165_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][10] ),
    .A2(net593),
    .A1(\top_ihp.oisc.regs[61][10] ));
 sg13g2_buf_1 _21614_ (.A(_05046_),
    .X(_05166_));
 sg13g2_a22oi_1 _21615_ (.Y(_05167_),
    .B1(_05166_),
    .B2(\top_ihp.oisc.regs[62][10] ),
    .A2(net459),
    .A1(\top_ihp.oisc.regs[56][10] ));
 sg13g2_a22oi_1 _21616_ (.Y(_05168_),
    .B1(net602),
    .B2(\top_ihp.oisc.regs[59][10] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][10] ));
 sg13g2_nand4_1 _21617_ (.B(_05165_),
    .C(_05167_),
    .A(_05163_),
    .Y(_05169_),
    .D(_05168_));
 sg13g2_buf_8 _21618_ (.A(_04995_),
    .X(_05170_));
 sg13g2_buf_8 _21619_ (.A(net591),
    .X(_05171_));
 sg13g2_a22oi_1 _21620_ (.Y(_05172_),
    .B1(_05171_),
    .B2(\top_ihp.oisc.regs[52][10] ),
    .A2(net267),
    .A1(\top_ihp.oisc.regs[38][10] ));
 sg13g2_buf_8 _21621_ (.A(net616),
    .X(_05173_));
 sg13g2_buf_2 _21622_ (.A(_05011_),
    .X(_05174_));
 sg13g2_a22oi_1 _21623_ (.Y(_05175_),
    .B1(_05174_),
    .B2(\top_ihp.oisc.regs[51][10] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][10] ));
 sg13g2_nand2_1 _21624_ (.Y(_05176_),
    .A(_05172_),
    .B(_05175_));
 sg13g2_buf_8 _21625_ (.A(net603),
    .X(_05177_));
 sg13g2_a22oi_1 _21626_ (.Y(_05178_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[58][10] ),
    .A2(net606),
    .A1(\top_ihp.oisc.regs[54][10] ));
 sg13g2_buf_1 _21627_ (.A(_04875_),
    .X(_05179_));
 sg13g2_buf_1 _21628_ (.A(net600),
    .X(_05180_));
 sg13g2_a22oi_1 _21629_ (.Y(_05181_),
    .B1(net440),
    .B2(\top_ihp.oisc.regs[2][10] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][10] ));
 sg13g2_buf_1 _21630_ (.A(_04974_),
    .X(_05182_));
 sg13g2_buf_1 _21631_ (.A(_05003_),
    .X(_05183_));
 sg13g2_a22oi_1 _21632_ (.Y(_05184_),
    .B1(net579),
    .B2(\top_ihp.oisc.regs[48][10] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][10] ));
 sg13g2_buf_1 _21633_ (.A(_05039_),
    .X(_05185_));
 sg13g2_a22oi_1 _21634_ (.Y(_05186_),
    .B1(net578),
    .B2(\top_ihp.oisc.regs[50][10] ),
    .A2(net462),
    .A1(\top_ihp.oisc.regs[36][10] ));
 sg13g2_nand4_1 _21635_ (.B(_05181_),
    .C(_05184_),
    .A(_05178_),
    .Y(_05187_),
    .D(_05186_));
 sg13g2_buf_8 _21636_ (.A(net596),
    .X(_05188_));
 sg13g2_buf_8 _21637_ (.A(net449),
    .X(_05189_));
 sg13g2_a22oi_1 _21638_ (.Y(_05190_),
    .B1(_05189_),
    .B2(\top_ihp.oisc.regs[41][10] ),
    .A2(_05188_),
    .A1(\top_ihp.oisc.regs[63][10] ));
 sg13g2_buf_8 _21639_ (.A(net476),
    .X(_05191_));
 sg13g2_buf_8 _21640_ (.A(_05076_),
    .X(_05192_));
 sg13g2_buf_8 _21641_ (.A(net438),
    .X(_05193_));
 sg13g2_a22oi_1 _21642_ (.Y(_05194_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][10] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][10] ));
 sg13g2_a22oi_1 _21643_ (.Y(_05195_),
    .B1(net607),
    .B2(\top_ihp.oisc.regs[31][10] ),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][10] ));
 sg13g2_buf_1 _21644_ (.A(_05015_),
    .X(_05196_));
 sg13g2_a22oi_1 _21645_ (.Y(_05197_),
    .B1(net577),
    .B2(\top_ihp.oisc.regs[4][10] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][10] ));
 sg13g2_and2_1 _21646_ (.A(_05195_),
    .B(_05197_),
    .X(_05198_));
 sg13g2_and2_1 _21647_ (.A(net703),
    .B(_04929_),
    .X(_05199_));
 sg13g2_buf_1 _21648_ (.A(_05199_),
    .X(_05200_));
 sg13g2_buf_2 _21649_ (.A(net646),
    .X(_05201_));
 sg13g2_buf_1 _21650_ (.A(net803),
    .X(_05202_));
 sg13g2_and2_1 _21651_ (.A(net697),
    .B(net722),
    .X(_05203_));
 sg13g2_buf_1 _21652_ (.A(_05203_),
    .X(_05204_));
 sg13g2_a22oi_1 _21653_ (.Y(_05205_),
    .B1(net645),
    .B2(\top_ihp.oisc.regs[16][10] ),
    .A2(net764),
    .A1(_07534_));
 sg13g2_inv_1 _21654_ (.Y(_05206_),
    .A(_05205_));
 sg13g2_a221oi_1 _21655_ (.B2(\top_ihp.oisc.regs[30][10] ),
    .C1(_05206_),
    .B1(_05201_),
    .A1(\top_ihp.oisc.regs[40][10] ),
    .Y(_05207_),
    .A2(net451));
 sg13g2_nand4_1 _21656_ (.B(_05194_),
    .C(_05198_),
    .A(_05190_),
    .Y(_05208_),
    .D(_05207_));
 sg13g2_nor4_2 _21657_ (.A(_05169_),
    .B(_05176_),
    .C(_05187_),
    .Y(_05209_),
    .D(_05208_));
 sg13g2_buf_8 _21658_ (.A(_04810_),
    .X(_05210_));
 sg13g2_buf_8 _21659_ (.A(_05104_),
    .X(_05211_));
 sg13g2_a21oi_1 _21660_ (.A1(_00117_),
    .A2(_05210_),
    .Y(_05212_),
    .B1(net153));
 sg13g2_a21oi_1 _21661_ (.A1(_07534_),
    .A2(net709),
    .Y(_05213_),
    .B1(_05212_));
 sg13g2_a21oi_1 _21662_ (.A1(_05162_),
    .A2(_05209_),
    .Y(_00295_),
    .B1(_05213_));
 sg13g2_buf_8 _21663_ (.A(_04969_),
    .X(_05214_));
 sg13g2_buf_8 _21664_ (.A(net575),
    .X(_05215_));
 sg13g2_a22oi_1 _21665_ (.Y(_05216_),
    .B1(net267),
    .B2(\top_ihp.oisc.regs[38][11] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[54][11] ));
 sg13g2_buf_2 _21666_ (.A(_04875_),
    .X(_05217_));
 sg13g2_a22oi_1 _21667_ (.Y(_05218_),
    .B1(net436),
    .B2(\top_ihp.oisc.regs[33][11] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][11] ));
 sg13g2_buf_8 _21668_ (.A(net451),
    .X(_05219_));
 sg13g2_a22oi_1 _21669_ (.Y(_05220_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][11] ),
    .A2(net578),
    .A1(\top_ihp.oisc.regs[50][11] ));
 sg13g2_buf_2 _21670_ (.A(_05079_),
    .X(_05221_));
 sg13g2_a22oi_1 _21671_ (.Y(_05222_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][11] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][11] ));
 sg13g2_nand4_1 _21672_ (.B(_05218_),
    .C(_05220_),
    .A(_05216_),
    .Y(_05223_),
    .D(_05222_));
 sg13g2_buf_8 _21673_ (.A(net462),
    .X(_05224_));
 sg13g2_a22oi_1 _21674_ (.Y(_05225_),
    .B1(net270),
    .B2(\top_ihp.oisc.regs[46][11] ),
    .A2(net262),
    .A1(\top_ihp.oisc.regs[36][11] ));
 sg13g2_buf_2 _21675_ (.A(_04965_),
    .X(_05226_));
 sg13g2_a22oi_1 _21676_ (.Y(_05227_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][11] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[32][11] ));
 sg13g2_a22oi_1 _21677_ (.Y(_05228_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][11] ),
    .A2(net581),
    .A1(\top_ihp.oisc.regs[51][11] ));
 sg13g2_a22oi_1 _21678_ (.Y(_05229_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[52][11] ),
    .A2(net594),
    .A1(\top_ihp.oisc.regs[62][11] ));
 sg13g2_nand4_1 _21679_ (.B(_05227_),
    .C(_05228_),
    .A(_05225_),
    .Y(_05230_),
    .D(_05229_));
 sg13g2_a22oi_1 _21680_ (.Y(_05231_),
    .B1(net454),
    .B2(\top_ihp.oisc.regs[34][11] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][11] ));
 sg13g2_a22oi_1 _21681_ (.Y(_05232_),
    .B1(net460),
    .B2(\top_ihp.oisc.regs[43][11] ),
    .A2(_04998_),
    .A1(\top_ihp.oisc.regs[59][11] ));
 sg13g2_nand2_1 _21682_ (.Y(_05233_),
    .A(_05231_),
    .B(_05232_));
 sg13g2_a22oi_1 _21683_ (.Y(_05234_),
    .B1(_05035_),
    .B2(\top_ihp.oisc.regs[56][11] ),
    .A2(_04978_),
    .A1(\top_ihp.oisc.regs[49][11] ));
 sg13g2_nand2_1 _21684_ (.Y(_05235_),
    .A(\top_ihp.oisc.regs[61][11] ),
    .B(net593));
 sg13g2_and2_1 _21685_ (.A(net697),
    .B(_04929_),
    .X(_05236_));
 sg13g2_buf_2 _21686_ (.A(_05236_),
    .X(_05237_));
 sg13g2_buf_8 _21687_ (.A(_05237_),
    .X(_05238_));
 sg13g2_a22oi_1 _21688_ (.Y(_05239_),
    .B1(net576),
    .B2(\top_ihp.oisc.regs[30][11] ),
    .A2(net574),
    .A1(\top_ihp.oisc.regs[26][11] ));
 sg13g2_and2_1 _21689_ (.A(net725),
    .B(_04957_),
    .X(_05240_));
 sg13g2_buf_4 _21690_ (.X(_05241_),
    .A(_05240_));
 sg13g2_a22oi_1 _21691_ (.Y(_05242_),
    .B1(_05241_),
    .B2(\top_ihp.oisc.regs[19][11] ),
    .A2(net645),
    .A1(\top_ihp.oisc.regs[16][11] ));
 sg13g2_nand4_1 _21692_ (.B(_05235_),
    .C(_05239_),
    .A(_05234_),
    .Y(_05243_),
    .D(_05242_));
 sg13g2_nor2b_1 _21693_ (.A(net725),
    .B_N(_04957_),
    .Y(_05244_));
 sg13g2_buf_2 _21694_ (.A(_05244_),
    .X(_05245_));
 sg13g2_nor2_1 _21695_ (.A(_07570_),
    .B(_03679_),
    .Y(_05246_));
 sg13g2_a221oi_1 _21696_ (.B2(\top_ihp.oisc.regs[3][11] ),
    .C1(_05246_),
    .B1(_05245_),
    .A1(\top_ihp.oisc.regs[29][11] ),
    .Y(_05247_),
    .A2(_04892_));
 sg13g2_a22oi_1 _21697_ (.Y(_05248_),
    .B1(net587),
    .B2(\top_ihp.oisc.regs[23][11] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][11] ));
 sg13g2_a22oi_1 _21698_ (.Y(_05249_),
    .B1(net477),
    .B2(\top_ihp.oisc.regs[14][11] ),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][11] ));
 sg13g2_buf_1 _21699_ (.A(_04939_),
    .X(_05250_));
 sg13g2_a22oi_1 _21700_ (.Y(_05251_),
    .B1(net573),
    .B2(\top_ihp.oisc.regs[31][11] ),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][11] ));
 sg13g2_nand4_1 _21701_ (.B(_05248_),
    .C(_05249_),
    .A(_05247_),
    .Y(_05252_),
    .D(_05251_));
 sg13g2_nor3_1 _21702_ (.A(net699),
    .B(net694),
    .C(net679),
    .Y(_05253_));
 sg13g2_buf_2 _21703_ (.A(_05253_),
    .X(_05254_));
 sg13g2_buf_1 _21704_ (.A(_05254_),
    .X(_05255_));
 sg13g2_a22oi_1 _21705_ (.Y(_05256_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][11] ),
    .A2(_05154_),
    .A1(\top_ihp.oisc.regs[27][11] ));
 sg13g2_a22oi_1 _21706_ (.Y(_05257_),
    .B1(net608),
    .B2(\top_ihp.oisc.regs[1][11] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][11] ));
 sg13g2_mux2_1 _21707_ (.A0(\top_ihp.oisc.regs[22][11] ),
    .A1(\top_ihp.oisc.regs[18][11] ),
    .S(_04910_),
    .X(_05258_));
 sg13g2_a22oi_1 _21708_ (.Y(_05259_),
    .B1(net695),
    .B2(_05258_),
    .A2(_04898_),
    .A1(\top_ihp.oisc.regs[10][11] ));
 sg13g2_a22oi_1 _21709_ (.Y(_05260_),
    .B1(net577),
    .B2(\top_ihp.oisc.regs[4][11] ),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][11] ));
 sg13g2_nand4_1 _21710_ (.B(_05257_),
    .C(_05259_),
    .A(_05256_),
    .Y(_05261_),
    .D(_05260_));
 sg13g2_or4_1 _21711_ (.A(_05233_),
    .B(_05243_),
    .C(_05252_),
    .D(_05261_),
    .X(_05262_));
 sg13g2_nor3_1 _21712_ (.A(_05223_),
    .B(_05230_),
    .C(_05262_),
    .Y(_05263_));
 sg13g2_buf_1 _21713_ (.A(_04865_),
    .X(_05264_));
 sg13g2_a22oi_1 _21714_ (.Y(_05265_),
    .B1(net447),
    .B2(\top_ihp.oisc.regs[35][11] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][11] ));
 sg13g2_buf_1 _21715_ (.A(_05030_),
    .X(_05266_));
 sg13g2_a22oi_1 _21716_ (.Y(_05267_),
    .B1(net571),
    .B2(\top_ihp.oisc.regs[63][11] ),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[5][11] ));
 sg13g2_buf_8 _21717_ (.A(_05061_),
    .X(_05268_));
 sg13g2_a22oi_1 _21718_ (.Y(_05269_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][11] ),
    .A2(net570),
    .A1(\top_ihp.oisc.regs[57][11] ));
 sg13g2_a22oi_1 _21719_ (.Y(_05270_),
    .B1(net450),
    .B2(\top_ihp.oisc.regs[37][11] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[58][11] ));
 sg13g2_nand4_1 _21720_ (.B(_05267_),
    .C(_05269_),
    .A(_05265_),
    .Y(_05271_),
    .D(_05270_));
 sg13g2_buf_1 _21721_ (.A(net719),
    .X(_05272_));
 sg13g2_nor2_2 _21722_ (.A(net677),
    .B(_04947_),
    .Y(_05273_));
 sg13g2_a22oi_1 _21723_ (.Y(_05274_),
    .B1(_05273_),
    .B2(\top_ihp.oisc.regs[12][11] ),
    .A2(_05007_),
    .A1(\top_ihp.oisc.regs[2][11] ));
 sg13g2_a22oi_1 _21724_ (.Y(_05275_),
    .B1(_05019_),
    .B2(\top_ihp.oisc.regs[11][11] ),
    .A2(net609),
    .A1(\top_ihp.oisc.regs[15][11] ));
 sg13g2_buf_1 _21725_ (.A(_05021_),
    .X(_05276_));
 sg13g2_a22oi_1 _21726_ (.Y(_05277_),
    .B1(net569),
    .B2(\top_ihp.oisc.regs[9][11] ),
    .A2(net610),
    .A1(\top_ihp.oisc.regs[6][11] ));
 sg13g2_and2_1 _21727_ (.A(_05275_),
    .B(_05277_),
    .X(_05278_));
 sg13g2_o21ai_1 _21728_ (.B1(_05278_),
    .Y(_05279_),
    .A1(net688),
    .A2(_05274_));
 sg13g2_buf_1 _21729_ (.A(net689),
    .X(_05280_));
 sg13g2_buf_1 _21730_ (.A(_04829_),
    .X(_05281_));
 sg13g2_buf_1 _21731_ (.A(net667),
    .X(_05282_));
 sg13g2_mux2_1 _21732_ (.A0(\top_ihp.oisc.regs[28][11] ),
    .A1(\top_ihp.oisc.regs[20][11] ),
    .S(net644),
    .X(_05283_));
 sg13g2_a22oi_1 _21733_ (.Y(_05284_),
    .B1(_05283_),
    .B2(net650),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[24][11] ));
 sg13g2_a22oi_1 _21734_ (.Y(_05285_),
    .B1(net268),
    .B2(\top_ihp.oisc.regs[44][11] ),
    .A2(_05004_),
    .A1(\top_ihp.oisc.regs[48][11] ));
 sg13g2_o21ai_1 _21735_ (.B1(_05285_),
    .Y(_05286_),
    .A1(net668),
    .A2(_05284_));
 sg13g2_nor4_1 _21736_ (.A(net80),
    .B(_05271_),
    .C(_05279_),
    .D(_05286_),
    .Y(_05287_));
 sg13g2_a21oi_1 _21737_ (.A1(_00118_),
    .A2(net78),
    .Y(_05288_),
    .B1(net154));
 sg13g2_nor2_1 _21738_ (.A(_05246_),
    .B(_05288_),
    .Y(_05289_));
 sg13g2_a21oi_1 _21739_ (.A1(_05263_),
    .A2(_05287_),
    .Y(_00296_),
    .B1(_05289_));
 sg13g2_buf_1 _21740_ (.A(_04965_),
    .X(_05290_));
 sg13g2_a22oi_1 _21741_ (.Y(_05291_),
    .B1(net581),
    .B2(\top_ihp.oisc.regs[51][12] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[32][12] ));
 sg13g2_a22oi_1 _21742_ (.Y(_05292_),
    .B1(net579),
    .B2(\top_ihp.oisc.regs[48][12] ),
    .A2(net604),
    .A1(\top_ihp.oisc.regs[49][12] ));
 sg13g2_a22oi_1 _21743_ (.Y(_05293_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][12] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][12] ));
 sg13g2_buf_8 _21744_ (.A(_05044_),
    .X(_05294_));
 sg13g2_a22oi_1 _21745_ (.Y(_05295_),
    .B1(net261),
    .B2(\top_ihp.oisc.regs[44][12] ),
    .A2(net600),
    .A1(\top_ihp.oisc.regs[2][12] ));
 sg13g2_nand4_1 _21746_ (.B(_05292_),
    .C(_05293_),
    .A(_05291_),
    .Y(_05296_),
    .D(_05295_));
 sg13g2_buf_8 _21747_ (.A(_04998_),
    .X(_05297_));
 sg13g2_a22oi_1 _21748_ (.Y(_05298_),
    .B1(net594),
    .B2(\top_ihp.oisc.regs[62][12] ),
    .A2(net568),
    .A1(\top_ihp.oisc.regs[59][12] ));
 sg13g2_buf_1 _21749_ (.A(_05051_),
    .X(_05299_));
 sg13g2_buf_8 _21750_ (.A(_05094_),
    .X(_05300_));
 sg13g2_a22oi_1 _21751_ (.Y(_05301_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][12] ),
    .A2(net567),
    .A1(\top_ihp.oisc.regs[61][12] ));
 sg13g2_buf_2 _21752_ (.A(_04988_),
    .X(_05302_));
 sg13g2_a22oi_1 _21753_ (.Y(_05303_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[36][12] ),
    .A2(net474),
    .A1(\top_ihp.oisc.regs[33][12] ));
 sg13g2_a22oi_1 _21754_ (.Y(_05304_),
    .B1(net450),
    .B2(\top_ihp.oisc.regs[37][12] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][12] ));
 sg13g2_nand4_1 _21755_ (.B(_05301_),
    .C(_05303_),
    .A(_05298_),
    .Y(_05305_),
    .D(_05304_));
 sg13g2_a22oi_1 _21756_ (.Y(_05306_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][12] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[35][12] ));
 sg13g2_buf_8 _21757_ (.A(net451),
    .X(_05307_));
 sg13g2_a22oi_1 _21758_ (.Y(_05308_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][12] ),
    .A2(net273),
    .A1(\top_ihp.oisc.regs[56][12] ));
 sg13g2_buf_2 _21759_ (.A(_04983_),
    .X(_05309_));
 sg13g2_buf_2 _21760_ (.A(_05058_),
    .X(_05310_));
 sg13g2_a22oi_1 _21761_ (.Y(_05311_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[46][12] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][12] ));
 sg13g2_a22oi_1 _21762_ (.Y(_05312_),
    .B1(_04972_),
    .B2(\top_ihp.oisc.regs[15][12] ),
    .A2(_04722_),
    .A1(\top_ihp.oisc.regs[5][12] ));
 sg13g2_nor3_1 _21763_ (.A(net652),
    .B(_05017_),
    .C(_05312_),
    .Y(_05313_));
 sg13g2_a21oi_1 _21764_ (.A1(\top_ihp.oisc.regs[63][12] ),
    .A2(net596),
    .Y(_05314_),
    .B1(_05313_));
 sg13g2_nand4_1 _21765_ (.B(_05308_),
    .C(_05311_),
    .A(_05306_),
    .Y(_05315_),
    .D(_05314_));
 sg13g2_a22oi_1 _21766_ (.Y(_05316_),
    .B1(net645),
    .B2(\top_ihp.oisc.regs[16][12] ),
    .A2(net576),
    .A1(\top_ihp.oisc.regs[30][12] ));
 sg13g2_a22oi_1 _21767_ (.Y(_05317_),
    .B1(net574),
    .B2(\top_ihp.oisc.regs[26][12] ),
    .A2(net772),
    .A1(_07528_));
 sg13g2_nand2_1 _21768_ (.Y(_05318_),
    .A(_05316_),
    .B(_05317_));
 sg13g2_a21oi_1 _21769_ (.A1(\top_ihp.oisc.regs[50][12] ),
    .A2(net595),
    .Y(_05319_),
    .B1(_05318_));
 sg13g2_buf_1 _21770_ (.A(net477),
    .X(_05320_));
 sg13g2_buf_8 _21771_ (.A(net471),
    .X(_05321_));
 sg13g2_a22oi_1 _21772_ (.Y(_05322_),
    .B1(net257),
    .B2(\top_ihp.oisc.regs[10][12] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][12] ));
 sg13g2_a22oi_1 _21773_ (.Y(_05323_),
    .B1(_04894_),
    .B2(\top_ihp.oisc.regs[29][12] ),
    .A2(net617),
    .A1(\top_ihp.oisc.regs[7][12] ));
 sg13g2_a22oi_1 _21774_ (.Y(_05324_),
    .B1(net587),
    .B2(\top_ihp.oisc.regs[23][12] ),
    .A2(net573),
    .A1(\top_ihp.oisc.regs[31][12] ));
 sg13g2_a22oi_1 _21775_ (.Y(_05325_),
    .B1(net647),
    .B2(\top_ihp.oisc.regs[11][12] ),
    .A2(net597),
    .A1(\top_ihp.oisc.regs[9][12] ));
 sg13g2_buf_2 _21776_ (.A(_04792_),
    .X(_05326_));
 sg13g2_mux2_1 _21777_ (.A0(\top_ihp.oisc.regs[22][12] ),
    .A1(\top_ihp.oisc.regs[18][12] ),
    .S(net666),
    .X(_05327_));
 sg13g2_a22oi_1 _21778_ (.Y(_05328_),
    .B1(net695),
    .B2(_05327_),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][12] ));
 sg13g2_buf_1 _21779_ (.A(_04935_),
    .X(_05329_));
 sg13g2_a22oi_1 _21780_ (.Y(_05330_),
    .B1(net585),
    .B2(\top_ihp.oisc.regs[12][12] ),
    .A2(net565),
    .A1(\top_ihp.oisc.regs[1][12] ));
 sg13g2_and4_1 _21781_ (.A(_05324_),
    .B(_05325_),
    .C(_05328_),
    .D(_05330_),
    .X(_05331_));
 sg13g2_nand4_1 _21782_ (.B(_05322_),
    .C(_05323_),
    .A(_05319_),
    .Y(_05332_),
    .D(_05331_));
 sg13g2_nor4_1 _21783_ (.A(_05296_),
    .B(_05305_),
    .C(_05315_),
    .D(_05332_),
    .Y(_05333_));
 sg13g2_buf_8 _21784_ (.A(net454),
    .X(_05334_));
 sg13g2_nand2_1 _21785_ (.Y(_05335_),
    .A(\top_ihp.oisc.regs[34][12] ),
    .B(net256));
 sg13g2_a22oi_1 _21786_ (.Y(_05336_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][12] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][12] ));
 sg13g2_a22oi_1 _21787_ (.Y(_05337_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][12] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][12] ));
 sg13g2_a22oi_1 _21788_ (.Y(_05338_),
    .B1(net580),
    .B2(\top_ihp.oisc.regs[42][12] ),
    .A2(_04844_),
    .A1(\top_ihp.oisc.regs[47][12] ));
 sg13g2_nand4_1 _21789_ (.B(_05336_),
    .C(_05337_),
    .A(_05335_),
    .Y(_05339_),
    .D(_05338_));
 sg13g2_mux2_1 _21790_ (.A0(\top_ihp.oisc.regs[3][12] ),
    .A1(\top_ihp.oisc.regs[19][12] ),
    .S(net676),
    .X(_05340_));
 sg13g2_a22oi_1 _21791_ (.Y(_05341_),
    .B1(_04959_),
    .B2(_05340_),
    .A2(net468),
    .A1(\top_ihp.oisc.regs[6][12] ));
 sg13g2_buf_1 _21792_ (.A(net618),
    .X(_05342_));
 sg13g2_a22oi_1 _21793_ (.Y(_05343_),
    .B1(net598),
    .B2(\top_ihp.oisc.regs[4][12] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[17][12] ));
 sg13g2_buf_2 _21794_ (.A(_04816_),
    .X(_05344_));
 sg13g2_buf_1 _21795_ (.A(net584),
    .X(_05345_));
 sg13g2_a22oi_1 _21796_ (.Y(_05346_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][12] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][12] ));
 sg13g2_a22oi_1 _21797_ (.Y(_05347_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][12] ),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][12] ));
 sg13g2_nand4_1 _21798_ (.B(_05343_),
    .C(_05346_),
    .A(_05341_),
    .Y(_05348_),
    .D(_05347_));
 sg13g2_mux2_1 _21799_ (.A0(\top_ihp.oisc.regs[28][12] ),
    .A1(\top_ihp.oisc.regs[20][12] ),
    .S(_05282_),
    .X(_05349_));
 sg13g2_a22oi_1 _21800_ (.Y(_05350_),
    .B1(_05349_),
    .B2(net650),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[24][12] ));
 sg13g2_a22oi_1 _21801_ (.Y(_05351_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[52][12] ),
    .A2(net269),
    .A1(\top_ihp.oisc.regs[43][12] ));
 sg13g2_o21ai_1 _21802_ (.B1(_05351_),
    .Y(_05352_),
    .A1(net668),
    .A2(_05350_));
 sg13g2_nor4_1 _21803_ (.A(net80),
    .B(_05339_),
    .C(_05348_),
    .D(_05352_),
    .Y(_05353_));
 sg13g2_buf_8 _21804_ (.A(_04810_),
    .X(_05354_));
 sg13g2_a21oi_1 _21805_ (.A1(_00119_),
    .A2(net77),
    .Y(_05355_),
    .B1(net153));
 sg13g2_a21oi_1 _21806_ (.A1(_07528_),
    .A2(net709),
    .Y(_05356_),
    .B1(_05355_));
 sg13g2_a21oi_1 _21807_ (.A1(_05333_),
    .A2(_05353_),
    .Y(_00297_),
    .B1(_05356_));
 sg13g2_a22oi_1 _21808_ (.Y(_05357_),
    .B1(net447),
    .B2(\top_ihp.oisc.regs[35][13] ),
    .A2(net273),
    .A1(\top_ihp.oisc.regs[56][13] ));
 sg13g2_a22oi_1 _21809_ (.Y(_05358_),
    .B1(net452),
    .B2(\top_ihp.oisc.regs[39][13] ),
    .A2(net602),
    .A1(\top_ihp.oisc.regs[59][13] ));
 sg13g2_buf_8 _21810_ (.A(_04978_),
    .X(_05359_));
 sg13g2_a22oi_1 _21811_ (.Y(_05360_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][13] ),
    .A2(net563),
    .A1(\top_ihp.oisc.regs[49][13] ));
 sg13g2_buf_1 _21812_ (.A(_05039_),
    .X(_05361_));
 sg13g2_a22oi_1 _21813_ (.Y(_05362_),
    .B1(net562),
    .B2(\top_ihp.oisc.regs[50][13] ),
    .A2(net596),
    .A1(\top_ihp.oisc.regs[63][13] ));
 sg13g2_nand4_1 _21814_ (.B(_05358_),
    .C(_05360_),
    .A(_05357_),
    .Y(_05363_),
    .D(_05362_));
 sg13g2_a22oi_1 _21815_ (.Y(_05364_),
    .B1(net594),
    .B2(\top_ihp.oisc.regs[62][13] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][13] ));
 sg13g2_a22oi_1 _21816_ (.Y(_05365_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][13] ),
    .A2(net458),
    .A1(\top_ihp.oisc.regs[44][13] ));
 sg13g2_a22oi_1 _21817_ (.Y(_05366_),
    .B1(net453),
    .B2(\top_ihp.oisc.regs[45][13] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][13] ));
 sg13g2_buf_2 _21818_ (.A(_05027_),
    .X(_05367_));
 sg13g2_a22oi_1 _21819_ (.Y(_05368_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[43][13] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[58][13] ));
 sg13g2_nand4_1 _21820_ (.B(_05365_),
    .C(_05366_),
    .A(_05364_),
    .Y(_05369_),
    .D(_05368_));
 sg13g2_mux2_1 _21821_ (.A0(\top_ihp.oisc.regs[3][13] ),
    .A1(\top_ihp.oisc.regs[19][13] ),
    .S(net693),
    .X(_05370_));
 sg13g2_a22oi_1 _21822_ (.Y(_05371_),
    .B1(net692),
    .B2(_05370_),
    .A2(_05250_),
    .A1(\top_ihp.oisc.regs[31][13] ));
 sg13g2_a22oi_1 _21823_ (.Y(_05372_),
    .B1(_04893_),
    .B2(\top_ihp.oisc.regs[29][13] ),
    .A2(_04826_),
    .A1(\top_ihp.oisc.regs[14][13] ));
 sg13g2_a22oi_1 _21824_ (.Y(_05373_),
    .B1(net651),
    .B2(\top_ihp.oisc.regs[11][13] ),
    .A2(_05196_),
    .A1(\top_ihp.oisc.regs[4][13] ));
 sg13g2_a22oi_1 _21825_ (.Y(_05374_),
    .B1(net565),
    .B2(\top_ihp.oisc.regs[1][13] ),
    .A2(net653),
    .A1(\top_ihp.oisc.regs[15][13] ));
 sg13g2_and4_1 _21826_ (.A(_05371_),
    .B(_05372_),
    .C(_05373_),
    .D(_05374_),
    .X(_05375_));
 sg13g2_nand2_1 _21827_ (.Y(_05376_),
    .A(\top_ihp.oisc.regs[52][13] ),
    .B(net444));
 sg13g2_buf_1 _21828_ (.A(_04994_),
    .X(_05377_));
 sg13g2_a22oi_1 _21829_ (.Y(_05378_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][13] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[38][13] ));
 sg13g2_nand3_1 _21830_ (.B(_05376_),
    .C(_05378_),
    .A(_05375_),
    .Y(_05379_));
 sg13g2_buf_8 _21831_ (.A(net605),
    .X(_05380_));
 sg13g2_a22oi_1 _21832_ (.Y(_05381_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][13] ),
    .A2(net425),
    .A1(\top_ihp.oisc.regs[42][13] ));
 sg13g2_a22oi_1 _21833_ (.Y(_05382_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][13] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][13] ));
 sg13g2_buf_8 _21834_ (.A(_05052_),
    .X(_05383_));
 sg13g2_a22oi_1 _21835_ (.Y(_05384_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][13] ),
    .A2(net599),
    .A1(\top_ihp.oisc.regs[51][13] ));
 sg13g2_a22oi_1 _21836_ (.Y(_05385_),
    .B1(net262),
    .B2(\top_ihp.oisc.regs[36][13] ),
    .A2(net606),
    .A1(\top_ihp.oisc.regs[54][13] ));
 sg13g2_nand4_1 _21837_ (.B(_05382_),
    .C(_05384_),
    .A(_05381_),
    .Y(_05386_),
    .D(_05385_));
 sg13g2_nor4_1 _21838_ (.A(_05363_),
    .B(_05369_),
    .C(_05379_),
    .D(_05386_),
    .Y(_05387_));
 sg13g2_nand2_1 _21839_ (.Y(_05388_),
    .A(net699),
    .B(net670));
 sg13g2_a22oi_1 _21840_ (.Y(_05389_),
    .B1(net690),
    .B2(\top_ihp.oisc.regs[22][13] ),
    .A2(net797),
    .A1(\top_ihp.oisc.regs[20][13] ));
 sg13g2_a22oi_1 _21841_ (.Y(_05390_),
    .B1(_05204_),
    .B2(\top_ihp.oisc.regs[16][13] ),
    .A2(net764),
    .A1(net1034));
 sg13g2_o21ai_1 _21842_ (.B1(_05390_),
    .Y(_05391_),
    .A1(_05388_),
    .A2(_05389_));
 sg13g2_a21oi_1 _21843_ (.A1(\top_ihp.oisc.regs[33][13] ),
    .A2(net441),
    .Y(_05392_),
    .B1(_05391_));
 sg13g2_buf_1 _21844_ (.A(_05153_),
    .X(_05393_));
 sg13g2_a22oi_1 _21845_ (.Y(_05394_),
    .B1(_05255_),
    .B2(\top_ihp.oisc.regs[8][13] ),
    .A2(net561),
    .A1(\top_ihp.oisc.regs[27][13] ));
 sg13g2_a22oi_1 _21846_ (.Y(_05395_),
    .B1(_05276_),
    .B2(\top_ihp.oisc.regs[9][13] ),
    .A2(_04889_),
    .A1(\top_ihp.oisc.regs[13][13] ));
 sg13g2_and2_1 _21847_ (.A(_05394_),
    .B(_05395_),
    .X(_05396_));
 sg13g2_a22oi_1 _21848_ (.Y(_05397_),
    .B1(net456),
    .B2(\top_ihp.oisc.regs[46][13] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][13] ));
 sg13g2_buf_1 _21849_ (.A(_05003_),
    .X(_05398_));
 sg13g2_a22oi_1 _21850_ (.Y(_05399_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][13] ),
    .A2(net560),
    .A1(\top_ihp.oisc.regs[48][13] ));
 sg13g2_nand4_1 _21851_ (.B(_05396_),
    .C(_05397_),
    .A(_05392_),
    .Y(_05400_),
    .D(_05399_));
 sg13g2_buf_1 _21852_ (.A(net587),
    .X(_05401_));
 sg13g2_a22oi_1 _21853_ (.Y(_05402_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][13] ),
    .A2(_04921_),
    .A1(\top_ihp.oisc.regs[6][13] ));
 sg13g2_a22oi_1 _21854_ (.Y(_05403_),
    .B1(net257),
    .B2(\top_ihp.oisc.regs[10][13] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[17][13] ));
 sg13g2_mux2_1 _21855_ (.A0(\top_ihp.oisc.regs[30][13] ),
    .A1(\top_ihp.oisc.regs[26][13] ),
    .S(net654),
    .X(_05404_));
 sg13g2_a22oi_1 _21856_ (.Y(_05405_),
    .B1(net720),
    .B2(_05404_),
    .A2(net617),
    .A1(\top_ihp.oisc.regs[7][13] ));
 sg13g2_a22oi_1 _21857_ (.Y(_05406_),
    .B1(net464),
    .B2(\top_ihp.oisc.regs[28][13] ),
    .A2(net469),
    .A1(\top_ihp.oisc.regs[5][13] ));
 sg13g2_nand4_1 _21858_ (.B(_05403_),
    .C(_05405_),
    .A(_05402_),
    .Y(_05407_),
    .D(_05406_));
 sg13g2_a22oi_1 _21859_ (.Y(_05408_),
    .B1(_05273_),
    .B2(\top_ihp.oisc.regs[12][13] ),
    .A2(_05007_),
    .A1(\top_ihp.oisc.regs[2][13] ));
 sg13g2_buf_2 _21860_ (.A(net680),
    .X(_05409_));
 sg13g2_buf_1 _21861_ (.A(net797),
    .X(_05410_));
 sg13g2_nand3_1 _21862_ (.B(net643),
    .C(_05410_),
    .A(\top_ihp.oisc.regs[24][13] ),
    .Y(_05411_));
 sg13g2_buf_1 _21863_ (.A(net670),
    .X(_05412_));
 sg13g2_nand3_1 _21864_ (.B(net642),
    .C(_05126_),
    .A(\top_ihp.oisc.regs[18][13] ),
    .Y(_05413_));
 sg13g2_a21oi_1 _21865_ (.A1(_05411_),
    .A2(_05413_),
    .Y(_05414_),
    .B1(net650));
 sg13g2_a221oi_1 _21866_ (.B2(\top_ihp.oisc.regs[21][13] ),
    .C1(_05414_),
    .B1(_04903_),
    .A1(\top_ihp.oisc.regs[25][13] ),
    .Y(_05415_),
    .A2(_05344_));
 sg13g2_o21ai_1 _21867_ (.B1(_05415_),
    .Y(_05416_),
    .A1(_05272_),
    .A2(_05408_));
 sg13g2_nor4_1 _21868_ (.A(net80),
    .B(_05400_),
    .C(_05407_),
    .D(_05416_),
    .Y(_05417_));
 sg13g2_buf_1 _21869_ (.A(net735),
    .X(_05418_));
 sg13g2_a21oi_1 _21870_ (.A1(_00120_),
    .A2(net77),
    .Y(_05419_),
    .B1(net153));
 sg13g2_a21oi_1 _21871_ (.A1(_07525_),
    .A2(net687),
    .Y(_05420_),
    .B1(_05419_));
 sg13g2_a21oi_1 _21872_ (.A1(_05387_),
    .A2(_05417_),
    .Y(_00298_),
    .B1(_05420_));
 sg13g2_a22oi_1 _21873_ (.Y(_05421_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][14] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[38][14] ));
 sg13g2_a22oi_1 _21874_ (.Y(_05422_),
    .B1(net454),
    .B2(\top_ihp.oisc.regs[34][14] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][14] ));
 sg13g2_a22oi_1 _21875_ (.Y(_05423_),
    .B1(net591),
    .B2(\top_ihp.oisc.regs[52][14] ),
    .A2(net460),
    .A1(\top_ihp.oisc.regs[43][14] ));
 sg13g2_buf_2 _21876_ (.A(_05011_),
    .X(_05424_));
 sg13g2_nor2_1 _21877_ (.A(net694),
    .B(net670),
    .Y(_05425_));
 sg13g2_a22oi_1 _21878_ (.Y(_05426_),
    .B1(_05069_),
    .B2(\top_ihp.oisc.regs[2][14] ),
    .A2(_05425_),
    .A1(\top_ihp.oisc.regs[8][14] ));
 sg13g2_nor3_1 _21879_ (.A(net650),
    .B(net719),
    .C(_05426_),
    .Y(_05427_));
 sg13g2_a21oi_1 _21880_ (.A1(\top_ihp.oisc.regs[51][14] ),
    .A2(net559),
    .Y(_05428_),
    .B1(_05427_));
 sg13g2_nand4_1 _21881_ (.B(_05422_),
    .C(_05423_),
    .A(_05421_),
    .Y(_05429_),
    .D(_05428_));
 sg13g2_a22oi_1 _21882_ (.Y(_05430_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[15][14] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][14] ));
 sg13g2_a22oi_1 _21883_ (.Y(_05431_),
    .B1(net577),
    .B2(\top_ihp.oisc.regs[4][14] ),
    .A2(net655),
    .A1(\top_ihp.oisc.regs[13][14] ));
 sg13g2_a22oi_1 _21884_ (.Y(_05432_),
    .B1(net565),
    .B2(\top_ihp.oisc.regs[1][14] ),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][14] ));
 sg13g2_a22oi_1 _21885_ (.Y(_05433_),
    .B1(net613),
    .B2(\top_ihp.oisc.regs[29][14] ),
    .A2(net657),
    .A1(\top_ihp.oisc.regs[7][14] ));
 sg13g2_nand4_1 _21886_ (.B(_05431_),
    .C(_05432_),
    .A(_05430_),
    .Y(_05434_),
    .D(_05433_));
 sg13g2_and2_1 _21887_ (.A(_07521_),
    .B(net803),
    .X(_05435_));
 sg13g2_a221oi_1 _21888_ (.B2(\top_ihp.oisc.regs[3][14] ),
    .C1(_05435_),
    .B1(_05245_),
    .A1(\top_ihp.oisc.regs[31][14] ),
    .Y(_05436_),
    .A2(_04939_));
 sg13g2_a22oi_1 _21889_ (.Y(_05437_),
    .B1(net584),
    .B2(\top_ihp.oisc.regs[27][14] ),
    .A2(net648),
    .A1(\top_ihp.oisc.regs[23][14] ));
 sg13g2_nand2_1 _21890_ (.Y(_05438_),
    .A(\top_ihp.oisc.regs[46][14] ),
    .B(_05058_));
 sg13g2_and2_1 _21891_ (.A(\top_ihp.oisc.regs[16][14] ),
    .B(net645),
    .X(_05439_));
 sg13g2_a221oi_1 _21892_ (.B2(\top_ihp.oisc.regs[19][14] ),
    .C1(_05439_),
    .B1(_05241_),
    .A1(\top_ihp.oisc.regs[30][14] ),
    .Y(_05440_),
    .A2(net646));
 sg13g2_nand4_1 _21893_ (.B(_05437_),
    .C(_05438_),
    .A(_05436_),
    .Y(_05441_),
    .D(_05440_));
 sg13g2_or2_1 _21894_ (.X(_05442_),
    .B(_05441_),
    .A(_05434_));
 sg13g2_a22oi_1 _21895_ (.Y(_05443_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][14] ),
    .A2(net453),
    .A1(\top_ihp.oisc.regs[45][14] ));
 sg13g2_a22oi_1 _21896_ (.Y(_05444_),
    .B1(net568),
    .B2(\top_ihp.oisc.regs[59][14] ),
    .A2(net604),
    .A1(\top_ihp.oisc.regs[49][14] ));
 sg13g2_a22oi_1 _21897_ (.Y(_05445_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][14] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[36][14] ));
 sg13g2_a22oi_1 _21898_ (.Y(_05446_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][14] ),
    .A2(net459),
    .A1(\top_ihp.oisc.regs[56][14] ));
 sg13g2_nand4_1 _21899_ (.B(_05444_),
    .C(_05445_),
    .A(_05443_),
    .Y(_05447_),
    .D(_05446_));
 sg13g2_a22oi_1 _21900_ (.Y(_05448_),
    .B1(net434),
    .B2(\top_ihp.oisc.regs[32][14] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][14] ));
 sg13g2_a22oi_1 _21901_ (.Y(_05449_),
    .B1(net595),
    .B2(\top_ihp.oisc.regs[50][14] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[33][14] ));
 sg13g2_a22oi_1 _21902_ (.Y(_05450_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[63][14] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[54][14] ));
 sg13g2_a22oi_1 _21903_ (.Y(_05451_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][14] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][14] ));
 sg13g2_nand4_1 _21904_ (.B(_05449_),
    .C(_05450_),
    .A(_05448_),
    .Y(_05452_),
    .D(_05451_));
 sg13g2_nor4_1 _21905_ (.A(_05429_),
    .B(_05442_),
    .C(_05447_),
    .D(_05452_),
    .Y(_05453_));
 sg13g2_and3_1 _21906_ (.X(_05454_),
    .A(_04775_),
    .B(_04791_),
    .C(_04807_));
 sg13g2_a22oi_1 _21907_ (.Y(_05455_),
    .B1(net452),
    .B2(\top_ihp.oisc.regs[39][14] ),
    .A2(net457),
    .A1(\top_ihp.oisc.regs[35][14] ));
 sg13g2_a22oi_1 _21908_ (.Y(_05456_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][14] ),
    .A2(net458),
    .A1(\top_ihp.oisc.regs[44][14] ));
 sg13g2_a22oi_1 _21909_ (.Y(_05457_),
    .B1(net582),
    .B2(\top_ihp.oisc.regs[62][14] ),
    .A2(net615),
    .A1(\top_ihp.oisc.regs[55][14] ));
 sg13g2_a22oi_1 _21910_ (.Y(_05458_),
    .B1(net560),
    .B2(\top_ihp.oisc.regs[48][14] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][14] ));
 sg13g2_nand4_1 _21911_ (.B(_05456_),
    .C(_05457_),
    .A(_05455_),
    .Y(_05459_),
    .D(_05458_));
 sg13g2_buf_1 _21912_ (.A(net651),
    .X(_05460_));
 sg13g2_a22oi_1 _21913_ (.Y(_05461_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][14] ),
    .A2(net470),
    .A1(\top_ihp.oisc.regs[21][14] ));
 sg13g2_buf_8 _21914_ (.A(net569),
    .X(_05462_));
 sg13g2_a22oi_1 _21915_ (.Y(_05463_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[9][14] ),
    .A2(net469),
    .A1(\top_ihp.oisc.regs[5][14] ));
 sg13g2_buf_1 _21916_ (.A(net666),
    .X(_05464_));
 sg13g2_mux2_1 _21917_ (.A0(\top_ihp.oisc.regs[14][14] ),
    .A1(\top_ihp.oisc.regs[10][14] ),
    .S(net641),
    .X(_05465_));
 sg13g2_nand3_1 _21918_ (.B(_04778_),
    .C(_05465_),
    .A(net677),
    .Y(_05466_));
 sg13g2_buf_1 _21919_ (.A(net585),
    .X(_05467_));
 sg13g2_a22oi_1 _21920_ (.Y(_05468_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][14] ),
    .A2(net610),
    .A1(\top_ihp.oisc.regs[6][14] ));
 sg13g2_nand4_1 _21921_ (.B(_05463_),
    .C(_05466_),
    .A(_05461_),
    .Y(_05469_),
    .D(_05468_));
 sg13g2_mux2_1 _21922_ (.A0(\top_ihp.oisc.regs[28][14] ),
    .A1(\top_ihp.oisc.regs[20][14] ),
    .S(net642),
    .X(_05470_));
 sg13g2_a22oi_1 _21923_ (.Y(_05471_),
    .B1(_05470_),
    .B2(_05135_),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[24][14] ));
 sg13g2_buf_1 _21924_ (.A(_04882_),
    .X(_05472_));
 sg13g2_mux2_1 _21925_ (.A0(\top_ihp.oisc.regs[26][14] ),
    .A1(\top_ihp.oisc.regs[18][14] ),
    .S(net667),
    .X(_05473_));
 sg13g2_buf_1 _21926_ (.A(net641),
    .X(_05474_));
 sg13g2_a22oi_1 _21927_ (.Y(_05475_),
    .B1(_05473_),
    .B2(net556),
    .A2(net557),
    .A1(\top_ihp.oisc.regs[22][14] ));
 sg13g2_nand2b_1 _21928_ (.Y(_05476_),
    .B(net671),
    .A_N(_05475_));
 sg13g2_o21ai_1 _21929_ (.B1(_05476_),
    .Y(_05477_),
    .A1(net668),
    .A2(_05471_));
 sg13g2_nor4_1 _21930_ (.A(_05454_),
    .B(_05459_),
    .C(_05469_),
    .D(_05477_),
    .Y(_05478_));
 sg13g2_a21oi_1 _21931_ (.A1(_00121_),
    .A2(net78),
    .Y(_05479_),
    .B1(net154));
 sg13g2_nor2_1 _21932_ (.A(_05435_),
    .B(_05479_),
    .Y(_05480_));
 sg13g2_a21oi_1 _21933_ (.A1(_05453_),
    .A2(_05478_),
    .Y(_00299_),
    .B1(_05480_));
 sg13g2_buf_2 _21934_ (.A(_05054_),
    .X(_05481_));
 sg13g2_nand2_1 _21935_ (.Y(_05482_),
    .A(\top_ihp.oisc.regs[35][15] ),
    .B(net420));
 sg13g2_a22oi_1 _21936_ (.Y(_05483_),
    .B1(net262),
    .B2(\top_ihp.oisc.regs[36][15] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[54][15] ));
 sg13g2_a22oi_1 _21937_ (.Y(_05484_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][15] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[32][15] ));
 sg13g2_buf_8 _21938_ (.A(_04908_),
    .X(_05485_));
 sg13g2_a22oi_1 _21939_ (.Y(_05486_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[63][15] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[5][15] ));
 sg13g2_and4_1 _21940_ (.A(_05482_),
    .B(_05483_),
    .C(_05484_),
    .D(_05486_),
    .X(_05487_));
 sg13g2_mux2_1 _21941_ (.A0(\top_ihp.oisc.regs[3][15] ),
    .A1(\top_ihp.oisc.regs[19][15] ),
    .S(_04952_),
    .X(_05488_));
 sg13g2_a22oi_1 _21942_ (.Y(_05489_),
    .B1(net692),
    .B2(_05488_),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][15] ));
 sg13g2_a22oi_1 _21943_ (.Y(_05490_),
    .B1(net597),
    .B2(\top_ihp.oisc.regs[9][15] ),
    .A2(net464),
    .A1(\top_ihp.oisc.regs[28][15] ));
 sg13g2_a22oi_1 _21944_ (.Y(_05491_),
    .B1(net561),
    .B2(\top_ihp.oisc.regs[27][15] ),
    .A2(_05015_),
    .A1(\top_ihp.oisc.regs[4][15] ));
 sg13g2_a22oi_1 _21945_ (.Y(_05492_),
    .B1(net647),
    .B2(\top_ihp.oisc.regs[11][15] ),
    .A2(_04925_),
    .A1(\top_ihp.oisc.regs[15][15] ));
 sg13g2_nand4_1 _21946_ (.B(_05490_),
    .C(_05491_),
    .A(_05489_),
    .Y(_05493_),
    .D(_05492_));
 sg13g2_a22oi_1 _21947_ (.Y(_05494_),
    .B1(net471),
    .B2(\top_ihp.oisc.regs[10][15] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][15] ));
 sg13g2_a22oi_1 _21948_ (.Y(_05495_),
    .B1(net608),
    .B2(\top_ihp.oisc.regs[1][15] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][15] ));
 sg13g2_and2_1 _21949_ (.A(\top_ihp.oisc.regs[23][15] ),
    .B(_05140_),
    .X(_05496_));
 sg13g2_a221oi_1 _21950_ (.B2(\top_ihp.oisc.regs[21][15] ),
    .C1(_05496_),
    .B1(net583),
    .A1(\top_ihp.oisc.regs[17][15] ),
    .Y(_05497_),
    .A2(net586));
 sg13g2_nand3_1 _21951_ (.B(_05495_),
    .C(_05497_),
    .A(_05494_),
    .Y(_05498_));
 sg13g2_mux2_1 _21952_ (.A0(\top_ihp.oisc.regs[24][15] ),
    .A1(\top_ihp.oisc.regs[16][15] ),
    .S(net667),
    .X(_05499_));
 sg13g2_a22oi_1 _21953_ (.Y(_05500_),
    .B1(_05499_),
    .B2(net652),
    .A2(net557),
    .A1(\top_ihp.oisc.regs[20][15] ));
 sg13g2_nor2_1 _21954_ (.A(net689),
    .B(_05500_),
    .Y(_05501_));
 sg13g2_a22oi_1 _21955_ (.Y(_05502_),
    .B1(net673),
    .B2(\top_ihp.oisc.regs[8][15] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[6][15] ));
 sg13g2_a22oi_1 _21956_ (.Y(_05503_),
    .B1(net459),
    .B2(\top_ihp.oisc.regs[56][15] ),
    .A2(net563),
    .A1(\top_ihp.oisc.regs[49][15] ));
 sg13g2_o21ai_1 _21957_ (.B1(_05503_),
    .Y(_05504_),
    .A1(net688),
    .A2(_05502_));
 sg13g2_nor4_1 _21958_ (.A(_05493_),
    .B(_05498_),
    .C(_05501_),
    .D(_05504_),
    .Y(_05505_));
 sg13g2_a22oi_1 _21959_ (.Y(_05506_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][15] ),
    .A2(_05088_),
    .A1(\top_ihp.oisc.regs[37][15] ));
 sg13g2_a22oi_1 _21960_ (.Y(_05507_),
    .B1(net570),
    .B2(\top_ihp.oisc.regs[57][15] ),
    .A2(_05046_),
    .A1(\top_ihp.oisc.regs[62][15] ));
 sg13g2_a22oi_1 _21961_ (.Y(_05508_),
    .B1(net458),
    .B2(\top_ihp.oisc.regs[44][15] ),
    .A2(_05027_),
    .A1(\top_ihp.oisc.regs[43][15] ));
 sg13g2_a22oi_1 _21962_ (.Y(_05509_),
    .B1(_04994_),
    .B2(\top_ihp.oisc.regs[38][15] ),
    .A2(net615),
    .A1(\top_ihp.oisc.regs[55][15] ));
 sg13g2_nand4_1 _21963_ (.B(_05507_),
    .C(_05508_),
    .A(_05506_),
    .Y(_05510_),
    .D(_05509_));
 sg13g2_a22oi_1 _21964_ (.Y(_05511_),
    .B1(net474),
    .B2(\top_ihp.oisc.regs[33][15] ),
    .A2(net476),
    .A1(\top_ihp.oisc.regs[47][15] ));
 sg13g2_a22oi_1 _21965_ (.Y(_05512_),
    .B1(net591),
    .B2(\top_ihp.oisc.regs[52][15] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][15] ));
 sg13g2_nand2_1 _21966_ (.Y(_05513_),
    .A(_05511_),
    .B(_05512_));
 sg13g2_buf_2 _21967_ (.A(_04892_),
    .X(_05514_));
 sg13g2_a22oi_1 _21968_ (.Y(_05515_),
    .B1(net585),
    .B2(\top_ihp.oisc.regs[12][15] ),
    .A2(net555),
    .A1(\top_ihp.oisc.regs[29][15] ));
 sg13g2_a22oi_1 _21969_ (.Y(_05516_),
    .B1(net607),
    .B2(\top_ihp.oisc.regs[31][15] ),
    .A2(net477),
    .A1(\top_ihp.oisc.regs[14][15] ));
 sg13g2_nand2_1 _21970_ (.Y(_05517_),
    .A(\top_ihp.oisc.regs[40][15] ),
    .B(net451));
 sg13g2_and2_1 _21971_ (.A(net697),
    .B(net721),
    .X(_05518_));
 sg13g2_buf_1 _21972_ (.A(_05518_),
    .X(_05519_));
 sg13g2_buf_2 _21973_ (.A(_05519_),
    .X(_05520_));
 sg13g2_a22oi_1 _21974_ (.Y(_05521_),
    .B1(net720),
    .B2(\top_ihp.oisc.regs[30][15] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[22][15] ));
 sg13g2_nand2_1 _21975_ (.Y(_05522_),
    .A(net1036),
    .B(net803));
 sg13g2_o21ai_1 _21976_ (.B1(_05522_),
    .Y(_05523_),
    .A1(net672),
    .A2(_05521_));
 sg13g2_a221oi_1 _21977_ (.B2(\top_ihp.oisc.regs[18][15] ),
    .C1(_05523_),
    .B1(net554),
    .A1(\top_ihp.oisc.regs[26][15] ),
    .Y(_05524_),
    .A2(net574));
 sg13g2_nand4_1 _21978_ (.B(_05516_),
    .C(_05517_),
    .A(_05515_),
    .Y(_05525_),
    .D(_05524_));
 sg13g2_nor3_1 _21979_ (.A(_05510_),
    .B(_05513_),
    .C(_05525_),
    .Y(_05526_));
 sg13g2_a22oi_1 _21980_ (.Y(_05527_),
    .B1(net603),
    .B2(\top_ihp.oisc.regs[58][15] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][15] ));
 sg13g2_a22oi_1 _21981_ (.Y(_05528_),
    .B1(net456),
    .B2(\top_ihp.oisc.regs[46][15] ),
    .A2(_05011_),
    .A1(\top_ihp.oisc.regs[51][15] ));
 sg13g2_a22oi_1 _21982_ (.Y(_05529_),
    .B1(net593),
    .B2(\top_ihp.oisc.regs[61][15] ),
    .A2(net600),
    .A1(\top_ihp.oisc.regs[2][15] ));
 sg13g2_a22oi_1 _21983_ (.Y(_05530_),
    .B1(net454),
    .B2(\top_ihp.oisc.regs[34][15] ),
    .A2(_04998_),
    .A1(\top_ihp.oisc.regs[59][15] ));
 sg13g2_nand4_1 _21984_ (.B(_05528_),
    .C(_05529_),
    .A(_05527_),
    .Y(_05531_),
    .D(_05530_));
 sg13g2_a22oi_1 _21985_ (.Y(_05532_),
    .B1(_05039_),
    .B2(\top_ihp.oisc.regs[50][15] ),
    .A2(net560),
    .A1(\top_ihp.oisc.regs[48][15] ));
 sg13g2_a22oi_1 _21986_ (.Y(_05533_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][15] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[45][15] ));
 sg13g2_nand2_1 _21987_ (.Y(_05534_),
    .A(_05532_),
    .B(_05533_));
 sg13g2_nor3_1 _21988_ (.A(_04810_),
    .B(_05531_),
    .C(_05534_),
    .Y(_05535_));
 sg13g2_and3_1 _21989_ (.X(_05536_),
    .A(_05505_),
    .B(_05526_),
    .C(_05535_));
 sg13g2_a21o_1 _21990_ (.A2(net79),
    .A1(_00122_),
    .B1(net154),
    .X(_05537_));
 sg13g2_a22oi_1 _21991_ (.Y(_00300_),
    .B1(_05537_),
    .B2(_05522_),
    .A2(_05536_),
    .A1(_05487_));
 sg13g2_buf_8 _21992_ (.A(_04810_),
    .X(_05538_));
 sg13g2_a22oi_1 _21993_ (.Y(_05539_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][16] ),
    .A2(net456),
    .A1(\top_ihp.oisc.regs[46][16] ));
 sg13g2_a22oi_1 _21994_ (.Y(_05540_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[54][16] ),
    .A2(_04921_),
    .A1(\top_ihp.oisc.regs[6][16] ));
 sg13g2_a22oi_1 _21995_ (.Y(_05541_),
    .B1(net599),
    .B2(\top_ihp.oisc.regs[51][16] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][16] ));
 sg13g2_a22oi_1 _21996_ (.Y(_05542_),
    .B1(net591),
    .B2(\top_ihp.oisc.regs[52][16] ),
    .A2(net462),
    .A1(\top_ihp.oisc.regs[36][16] ));
 sg13g2_nand4_1 _21997_ (.B(_05540_),
    .C(_05541_),
    .A(_05539_),
    .Y(_05543_),
    .D(_05542_));
 sg13g2_a22oi_1 _21998_ (.Y(_05544_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][16] ),
    .A2(_04890_),
    .A1(\top_ihp.oisc.regs[13][16] ));
 sg13g2_mux2_1 _21999_ (.A0(\top_ihp.oisc.regs[3][16] ),
    .A1(\top_ihp.oisc.regs[19][16] ),
    .S(net693),
    .X(_05545_));
 sg13g2_a22oi_1 _22000_ (.Y(_05546_),
    .B1(_05545_),
    .B2(net675),
    .A2(_05016_),
    .A1(\top_ihp.oisc.regs[4][16] ));
 sg13g2_buf_1 _22001_ (.A(net564),
    .X(_05547_));
 sg13g2_a22oi_1 _22002_ (.Y(_05548_),
    .B1(_05462_),
    .B2(\top_ihp.oisc.regs[9][16] ),
    .A2(_05547_),
    .A1(\top_ihp.oisc.regs[25][16] ));
 sg13g2_a22oi_1 _22003_ (.Y(_05549_),
    .B1(net257),
    .B2(\top_ihp.oisc.regs[10][16] ),
    .A2(net555),
    .A1(\top_ihp.oisc.regs[29][16] ));
 sg13g2_nand4_1 _22004_ (.B(_05546_),
    .C(_05548_),
    .A(_05544_),
    .Y(_05550_),
    .D(_05549_));
 sg13g2_a22oi_1 _22005_ (.Y(_05551_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][16] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[5][16] ));
 sg13g2_a22oi_1 _22006_ (.Y(_05552_),
    .B1(_05460_),
    .B2(\top_ihp.oisc.regs[11][16] ),
    .A2(net470),
    .A1(\top_ihp.oisc.regs[21][16] ));
 sg13g2_nor2_2 _22007_ (.A(net699),
    .B(net694),
    .Y(_05553_));
 sg13g2_mux2_1 _22008_ (.A0(\top_ihp.oisc.regs[14][16] ),
    .A1(\top_ihp.oisc.regs[12][16] ),
    .S(net656),
    .X(_05554_));
 sg13g2_a22oi_1 _22009_ (.Y(_05555_),
    .B1(_05554_),
    .B2(net650),
    .A2(_05553_),
    .A1(\top_ihp.oisc.regs[8][16] ));
 sg13g2_nand2b_1 _22010_ (.Y(_05556_),
    .B(_04778_),
    .A_N(_05555_));
 sg13g2_nand3_1 _22011_ (.B(_05552_),
    .C(_05556_),
    .A(_05551_),
    .Y(_05557_));
 sg13g2_nor4_1 _22012_ (.A(net76),
    .B(_05543_),
    .C(_05550_),
    .D(_05557_),
    .Y(_05558_));
 sg13g2_a22oi_1 _22013_ (.Y(_05559_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][16] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][16] ));
 sg13g2_a22oi_1 _22014_ (.Y(_05560_),
    .B1(net451),
    .B2(\top_ihp.oisc.regs[40][16] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][16] ));
 sg13g2_a22oi_1 _22015_ (.Y(_05561_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][16] ),
    .A2(_05009_),
    .A1(\top_ihp.oisc.regs[2][16] ));
 sg13g2_a22oi_1 _22016_ (.Y(_05562_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[32][16] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][16] ));
 sg13g2_nand4_1 _22017_ (.B(_05560_),
    .C(_05561_),
    .A(_05559_),
    .Y(_05563_),
    .D(_05562_));
 sg13g2_nand2_1 _22018_ (.Y(_05564_),
    .A(\top_ihp.oisc.regs[48][16] ),
    .B(net601));
 sg13g2_a22oi_1 _22019_ (.Y(_05565_),
    .B1(net273),
    .B2(\top_ihp.oisc.regs[56][16] ),
    .A2(net474),
    .A1(\top_ihp.oisc.regs[33][16] ));
 sg13g2_a22oi_1 _22020_ (.Y(_05566_),
    .B1(net571),
    .B2(\top_ihp.oisc.regs[63][16] ),
    .A2(net460),
    .A1(\top_ihp.oisc.regs[43][16] ));
 sg13g2_a22oi_1 _22021_ (.Y(_05567_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][16] ),
    .A2(net582),
    .A1(\top_ihp.oisc.regs[62][16] ));
 sg13g2_nand4_1 _22022_ (.B(_05565_),
    .C(_05566_),
    .A(_05564_),
    .Y(_05568_),
    .D(_05567_));
 sg13g2_a22oi_1 _22023_ (.Y(_05569_),
    .B1(net608),
    .B2(\top_ihp.oisc.regs[1][16] ),
    .A2(net609),
    .A1(\top_ihp.oisc.regs[15][16] ));
 sg13g2_a22oi_1 _22024_ (.Y(_05570_),
    .B1(_04834_),
    .B2(\top_ihp.oisc.regs[24][16] ),
    .A2(net618),
    .A1(\top_ihp.oisc.regs[17][16] ));
 sg13g2_nand2_1 _22025_ (.Y(_05571_),
    .A(\top_ihp.oisc.regs[26][16] ),
    .B(_04873_));
 sg13g2_nand2_1 _22026_ (.Y(_05572_),
    .A(\top_ihp.oisc.regs[18][16] ),
    .B(net670));
 sg13g2_nand2_1 _22027_ (.Y(_05573_),
    .A(net666),
    .B(net690));
 sg13g2_a21oi_1 _22028_ (.A1(_05571_),
    .A2(_05572_),
    .Y(_05574_),
    .B1(_05573_));
 sg13g2_a21oi_1 _22029_ (.A1(\top_ihp.oisc.regs[31][16] ),
    .A2(_05250_),
    .Y(_05575_),
    .B1(_05574_));
 sg13g2_mux2_1 _22030_ (.A0(\top_ihp.oisc.regs[28][16] ),
    .A1(\top_ihp.oisc.regs[20][16] ),
    .S(_05132_),
    .X(_05576_));
 sg13g2_nor2_1 _22031_ (.A(net672),
    .B(net689),
    .Y(_05577_));
 sg13g2_a22oi_1 _22032_ (.Y(_05578_),
    .B1(_05576_),
    .B2(_05577_),
    .A2(_04846_),
    .A1(\top_ihp.oisc.regs[7][16] ));
 sg13g2_and4_1 _22033_ (.A(_05569_),
    .B(_05570_),
    .C(_05575_),
    .D(_05578_),
    .X(_05579_));
 sg13g2_a22oi_1 _22034_ (.Y(_05580_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][16] ),
    .A2(net568),
    .A1(\top_ihp.oisc.regs[59][16] ));
 sg13g2_nand3_1 _22035_ (.B(net669),
    .C(net695),
    .A(\top_ihp.oisc.regs[22][16] ),
    .Y(_05581_));
 sg13g2_nand3_1 _22036_ (.B(net641),
    .C(net722),
    .A(\top_ihp.oisc.regs[16][16] ),
    .Y(_05582_));
 sg13g2_a22oi_1 _22037_ (.Y(_05583_),
    .B1(net646),
    .B2(\top_ihp.oisc.regs[30][16] ),
    .A2(net764),
    .A1(_07507_));
 sg13g2_nand3_1 _22038_ (.B(_05582_),
    .C(_05583_),
    .A(_05581_),
    .Y(_05584_));
 sg13g2_a21oi_1 _22039_ (.A1(\top_ihp.oisc.regs[38][16] ),
    .A2(net426),
    .Y(_05585_),
    .B1(_05584_));
 sg13g2_nand3_1 _22040_ (.B(_05580_),
    .C(_05585_),
    .A(_05579_),
    .Y(_05586_));
 sg13g2_a22oi_1 _22041_ (.Y(_05587_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][16] ),
    .A2(net595),
    .A1(\top_ihp.oisc.regs[50][16] ));
 sg13g2_a22oi_1 _22042_ (.Y(_05588_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[35][16] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][16] ));
 sg13g2_a22oi_1 _22043_ (.Y(_05589_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][16] ),
    .A2(net261),
    .A1(\top_ihp.oisc.regs[44][16] ));
 sg13g2_buf_8 _22044_ (.A(net563),
    .X(_05590_));
 sg13g2_buf_2 _22045_ (.A(_05088_),
    .X(_05591_));
 sg13g2_a22oi_1 _22046_ (.Y(_05592_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][16] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[49][16] ));
 sg13g2_nand4_1 _22047_ (.B(_05588_),
    .C(_05589_),
    .A(_05587_),
    .Y(_05593_),
    .D(_05592_));
 sg13g2_nor4_1 _22048_ (.A(_05563_),
    .B(_05568_),
    .C(_05586_),
    .D(_05593_),
    .Y(_05594_));
 sg13g2_a21oi_1 _22049_ (.A1(_00123_),
    .A2(_05354_),
    .Y(_05595_),
    .B1(_05211_));
 sg13g2_a21oi_1 _22050_ (.A1(_07507_),
    .A2(net687),
    .Y(_05596_),
    .B1(_05595_));
 sg13g2_a21oi_1 _22051_ (.A1(_05558_),
    .A2(_05594_),
    .Y(_00301_),
    .B1(_05596_));
 sg13g2_buf_1 _22052_ (.A(_04843_),
    .X(_05597_));
 sg13g2_a22oi_1 _22053_ (.Y(_05598_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][17] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][17] ));
 sg13g2_a22oi_1 _22054_ (.Y(_05599_),
    .B1(net599),
    .B2(\top_ihp.oisc.regs[51][17] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][17] ));
 sg13g2_a22oi_1 _22055_ (.Y(_05600_),
    .B1(net273),
    .B2(\top_ihp.oisc.regs[56][17] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][17] ));
 sg13g2_a22oi_1 _22056_ (.Y(_05601_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][17] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][17] ));
 sg13g2_nand4_1 _22057_ (.B(_05599_),
    .C(_05600_),
    .A(_05598_),
    .Y(_05602_),
    .D(_05601_));
 sg13g2_nand2_1 _22058_ (.Y(_05603_),
    .A(\top_ihp.oisc.regs[43][17] ),
    .B(net269));
 sg13g2_a22oi_1 _22059_ (.Y(_05604_),
    .B1(net578),
    .B2(\top_ihp.oisc.regs[50][17] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][17] ));
 sg13g2_a22oi_1 _22060_ (.Y(_05605_),
    .B1(net567),
    .B2(\top_ihp.oisc.regs[61][17] ),
    .A2(net563),
    .A1(\top_ihp.oisc.regs[49][17] ));
 sg13g2_a22oi_1 _22061_ (.Y(_05606_),
    .B1(net571),
    .B2(\top_ihp.oisc.regs[63][17] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[58][17] ));
 sg13g2_nand4_1 _22062_ (.B(_05604_),
    .C(_05605_),
    .A(_05603_),
    .Y(_05607_),
    .D(_05606_));
 sg13g2_a221oi_1 _22063_ (.B2(_04690_),
    .C1(net997),
    .B1(_04718_),
    .A1(_04687_),
    .Y(_05608_),
    .A2(_04742_));
 sg13g2_buf_2 _22064_ (.A(_05608_),
    .X(_05609_));
 sg13g2_a22oi_1 _22065_ (.Y(_05610_),
    .B1(net690),
    .B2(\top_ihp.oisc.regs[30][17] ),
    .A2(net797),
    .A1(\top_ihp.oisc.regs[28][17] ));
 sg13g2_inv_1 _22066_ (.Y(_05611_),
    .A(_05610_));
 sg13g2_a22oi_1 _22067_ (.Y(_05612_),
    .B1(_04916_),
    .B2(\top_ihp.oisc.regs[18][17] ),
    .A2(net722),
    .A1(\top_ihp.oisc.regs[16][17] ));
 sg13g2_nand3_1 _22068_ (.B(net699),
    .C(net722),
    .A(\top_ihp.oisc.regs[20][17] ),
    .Y(_05613_));
 sg13g2_o21ai_1 _22069_ (.B1(_05613_),
    .Y(_05614_),
    .A1(net669),
    .A2(_05612_));
 sg13g2_a221oi_1 _22070_ (.B2(_05611_),
    .C1(_05614_),
    .B1(net718),
    .A1(net1035),
    .Y(_05615_),
    .A2(net772));
 sg13g2_a22oi_1 _22071_ (.Y(_05616_),
    .B1(net612),
    .B2(\top_ihp.oisc.regs[21][17] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][17] ));
 sg13g2_a22oi_1 _22072_ (.Y(_05617_),
    .B1(net561),
    .B2(\top_ihp.oisc.regs[27][17] ),
    .A2(net648),
    .A1(\top_ihp.oisc.regs[23][17] ));
 sg13g2_a22oi_1 _22073_ (.Y(_05618_),
    .B1(net597),
    .B2(\top_ihp.oisc.regs[9][17] ),
    .A2(net565),
    .A1(\top_ihp.oisc.regs[1][17] ));
 sg13g2_and4_1 _22074_ (.A(_05615_),
    .B(_05616_),
    .C(_05617_),
    .D(_05618_),
    .X(_05619_));
 sg13g2_buf_2 _22075_ (.A(_05046_),
    .X(_05620_));
 sg13g2_a22oi_1 _22076_ (.Y(_05621_),
    .B1(net553),
    .B2(\top_ihp.oisc.regs[62][17] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[54][17] ));
 sg13g2_a22oi_1 _22077_ (.Y(_05622_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][17] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[2][17] ));
 sg13g2_nand3_1 _22078_ (.B(_05621_),
    .C(_05622_),
    .A(_05619_),
    .Y(_05623_));
 sg13g2_a22oi_1 _22079_ (.Y(_05624_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][17] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][17] ));
 sg13g2_a22oi_1 _22080_ (.Y(_05625_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][17] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[36][17] ));
 sg13g2_a22oi_1 _22081_ (.Y(_05626_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[52][17] ),
    .A2(net579),
    .A1(\top_ihp.oisc.regs[48][17] ));
 sg13g2_a22oi_1 _22082_ (.Y(_05627_),
    .B1(net453),
    .B2(\top_ihp.oisc.regs[45][17] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][17] ));
 sg13g2_nand4_1 _22083_ (.B(_05625_),
    .C(_05626_),
    .A(_05624_),
    .Y(_05628_),
    .D(_05627_));
 sg13g2_nor4_1 _22084_ (.A(_05602_),
    .B(_05607_),
    .C(_05623_),
    .D(_05628_),
    .Y(_05629_));
 sg13g2_a22oi_1 _22085_ (.Y(_05630_),
    .B1(net261),
    .B2(\top_ihp.oisc.regs[44][17] ),
    .A2(net602),
    .A1(\top_ihp.oisc.regs[59][17] ));
 sg13g2_a22oi_1 _22086_ (.Y(_05631_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[46][17] ),
    .A2(net457),
    .A1(\top_ihp.oisc.regs[35][17] ));
 sg13g2_a22oi_1 _22087_ (.Y(_05632_),
    .B1(_04882_),
    .B2(\top_ihp.oisc.regs[22][17] ),
    .A2(_04880_),
    .A1(\top_ihp.oisc.regs[26][17] ));
 sg13g2_inv_1 _22088_ (.Y(_05633_),
    .A(_05632_));
 sg13g2_a22oi_1 _22089_ (.Y(_05634_),
    .B1(_04972_),
    .B2(\top_ihp.oisc.regs[14][17] ),
    .A2(_04722_),
    .A1(\top_ihp.oisc.regs[4][17] ));
 sg13g2_nor3_1 _22090_ (.A(net652),
    .B(net719),
    .C(_05634_),
    .Y(_05635_));
 sg13g2_a21oi_1 _22091_ (.A1(net671),
    .A2(_05633_),
    .Y(_05636_),
    .B1(_05635_));
 sg13g2_a22oi_1 _22092_ (.Y(_05637_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[41][17] ),
    .A2(net570),
    .A1(\top_ihp.oisc.regs[57][17] ));
 sg13g2_nand4_1 _22093_ (.B(_05631_),
    .C(_05636_),
    .A(_05630_),
    .Y(_05638_),
    .D(_05637_));
 sg13g2_mux2_1 _22094_ (.A0(\top_ihp.oisc.regs[3][17] ),
    .A1(\top_ihp.oisc.regs[19][17] ),
    .S(net676),
    .X(_05639_));
 sg13g2_a22oi_1 _22095_ (.Y(_05640_),
    .B1(net675),
    .B2(_05639_),
    .A2(net555),
    .A1(\top_ihp.oisc.regs[29][17] ));
 sg13g2_a22oi_1 _22096_ (.Y(_05641_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][17] ),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][17] ));
 sg13g2_a22oi_1 _22097_ (.Y(_05642_),
    .B1(net467),
    .B2(\top_ihp.oisc.regs[15][17] ),
    .A2(net471),
    .A1(\top_ihp.oisc.regs[10][17] ));
 sg13g2_a22oi_1 _22098_ (.Y(_05643_),
    .B1(net465),
    .B2(\top_ihp.oisc.regs[31][17] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[17][17] ));
 sg13g2_nand4_1 _22099_ (.B(_05641_),
    .C(_05642_),
    .A(_05640_),
    .Y(_05644_),
    .D(_05643_));
 sg13g2_a22oi_1 _22100_ (.Y(_05645_),
    .B1(net673),
    .B2(\top_ihp.oisc.regs[8][17] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[6][17] ));
 sg13g2_or2_1 _22101_ (.X(_05646_),
    .B(_05645_),
    .A(net688));
 sg13g2_a22oi_1 _22102_ (.Y(_05647_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][17] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[5][17] ));
 sg13g2_a22oi_1 _22103_ (.Y(_05648_),
    .B1(net473),
    .B2(\top_ihp.oisc.regs[13][17] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][17] ));
 sg13g2_nand3_1 _22104_ (.B(_05647_),
    .C(_05648_),
    .A(_05646_),
    .Y(_05649_));
 sg13g2_nor4_1 _22105_ (.A(net80),
    .B(_05638_),
    .C(_05644_),
    .D(_05649_),
    .Y(_05650_));
 sg13g2_a21oi_1 _22106_ (.A1(_00124_),
    .A2(net77),
    .Y(_05651_),
    .B1(net153));
 sg13g2_a21oi_1 _22107_ (.A1(_07517_),
    .A2(net687),
    .Y(_05652_),
    .B1(_05651_));
 sg13g2_a21oi_1 _22108_ (.A1(_05629_),
    .A2(_05650_),
    .Y(_00302_),
    .B1(_05652_));
 sg13g2_buf_1 _22109_ (.A(net718),
    .X(_05653_));
 sg13g2_mux2_1 _22110_ (.A0(\top_ihp.oisc.regs[20][18] ),
    .A1(\top_ihp.oisc.regs[16][18] ),
    .S(net652),
    .X(_05654_));
 sg13g2_buf_1 _22111_ (.A(net667),
    .X(_05655_));
 sg13g2_a22oi_1 _22112_ (.Y(_05656_),
    .B1(_05654_),
    .B2(net640),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][18] ));
 sg13g2_nor2_1 _22113_ (.A(_05280_),
    .B(_05656_),
    .Y(_05657_));
 sg13g2_a22oi_1 _22114_ (.Y(_05658_),
    .B1(net467),
    .B2(\top_ihp.oisc.regs[15][18] ),
    .A2(net472),
    .A1(\top_ihp.oisc.regs[29][18] ));
 sg13g2_a22oi_1 _22115_ (.Y(_05659_),
    .B1(_05467_),
    .B2(\top_ihp.oisc.regs[12][18] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[9][18] ));
 sg13g2_a22oi_1 _22116_ (.Y(_05660_),
    .B1(net257),
    .B2(\top_ihp.oisc.regs[10][18] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][18] ));
 sg13g2_mux2_1 _22117_ (.A0(\top_ihp.oisc.regs[3][18] ),
    .A1(\top_ihp.oisc.regs[19][18] ),
    .S(net676),
    .X(_05661_));
 sg13g2_nand2_1 _22118_ (.Y(_05662_),
    .A(net675),
    .B(_05661_));
 sg13g2_nand4_1 _22119_ (.B(_05659_),
    .C(_05660_),
    .A(_05658_),
    .Y(_05663_),
    .D(_05662_));
 sg13g2_nor3_1 _22120_ (.A(net79),
    .B(_05657_),
    .C(_05663_),
    .Y(_05664_));
 sg13g2_a22oi_1 _22121_ (.Y(_05665_),
    .B1(_05071_),
    .B2(\top_ihp.oisc.regs[34][18] ),
    .A2(_04869_),
    .A1(\top_ihp.oisc.regs[55][18] ));
 sg13g2_a22oi_1 _22122_ (.Y(_05666_),
    .B1(_05066_),
    .B2(\top_ihp.oisc.regs[52][18] ),
    .A2(_05046_),
    .A1(\top_ihp.oisc.regs[62][18] ));
 sg13g2_a22oi_1 _22123_ (.Y(_05667_),
    .B1(_05003_),
    .B2(\top_ihp.oisc.regs[48][18] ),
    .A2(_04974_),
    .A1(\top_ihp.oisc.regs[42][18] ));
 sg13g2_a22oi_1 _22124_ (.Y(_05668_),
    .B1(_05125_),
    .B2(\top_ihp.oisc.regs[26][18] ),
    .A2(net797),
    .A1(\top_ihp.oisc.regs[24][18] ));
 sg13g2_nand3_1 _22125_ (.B(net698),
    .C(_05125_),
    .A(\top_ihp.oisc.regs[18][18] ),
    .Y(_05669_));
 sg13g2_o21ai_1 _22126_ (.B1(_05669_),
    .Y(_05670_),
    .A1(_05132_),
    .A2(_05668_));
 sg13g2_a22oi_1 _22127_ (.Y(_05671_),
    .B1(_05670_),
    .B2(net641),
    .A2(_04988_),
    .A1(\top_ihp.oisc.regs[36][18] ));
 sg13g2_nand4_1 _22128_ (.B(_05666_),
    .C(_05667_),
    .A(_05665_),
    .Y(_05672_),
    .D(_05671_));
 sg13g2_a22oi_1 _22129_ (.Y(_05673_),
    .B1(_05030_),
    .B2(\top_ihp.oisc.regs[63][18] ),
    .A2(_04969_),
    .A1(\top_ihp.oisc.regs[54][18] ));
 sg13g2_a22oi_1 _22130_ (.Y(_05674_),
    .B1(_05088_),
    .B2(\top_ihp.oisc.regs[37][18] ),
    .A2(_05035_),
    .A1(\top_ihp.oisc.regs[56][18] ));
 sg13g2_a22oi_1 _22131_ (.Y(_05675_),
    .B1(_05061_),
    .B2(\top_ihp.oisc.regs[57][18] ),
    .A2(_05054_),
    .A1(\top_ihp.oisc.regs[35][18] ));
 sg13g2_a22oi_1 _22132_ (.Y(_05676_),
    .B1(_05051_),
    .B2(\top_ihp.oisc.regs[61][18] ),
    .A2(_04983_),
    .A1(\top_ihp.oisc.regs[58][18] ));
 sg13g2_nand4_1 _22133_ (.B(_05674_),
    .C(_05675_),
    .A(_05673_),
    .Y(_05677_),
    .D(_05676_));
 sg13g2_a22oi_1 _22134_ (.Y(_05678_),
    .B1(_04972_),
    .B2(\top_ihp.oisc.regs[14][18] ),
    .A2(_04722_),
    .A1(\top_ihp.oisc.regs[4][18] ));
 sg13g2_a22oi_1 _22135_ (.Y(_05679_),
    .B1(net673),
    .B2(\top_ihp.oisc.regs[8][18] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[6][18] ));
 sg13g2_o21ai_1 _22136_ (.B1(_05679_),
    .Y(_05680_),
    .A1(net641),
    .A2(_05678_));
 sg13g2_nor2b_1 _22137_ (.A(net688),
    .B_N(_05680_),
    .Y(_05681_));
 sg13g2_a22oi_1 _22138_ (.Y(_05682_),
    .B1(_05085_),
    .B2(\top_ihp.oisc.regs[40][18] ),
    .A2(_05043_),
    .A1(\top_ihp.oisc.regs[44][18] ));
 sg13g2_a22oi_1 _22139_ (.Y(_05683_),
    .B1(_05096_),
    .B2(\top_ihp.oisc.regs[60][18] ),
    .A2(_05093_),
    .A1(\top_ihp.oisc.regs[41][18] ));
 sg13g2_a22oi_1 _22140_ (.Y(_05684_),
    .B1(_04865_),
    .B2(\top_ihp.oisc.regs[53][18] ),
    .A2(_04843_),
    .A1(\top_ihp.oisc.regs[47][18] ));
 sg13g2_a22oi_1 _22141_ (.Y(_05685_),
    .B1(_04994_),
    .B2(\top_ihp.oisc.regs[38][18] ),
    .A2(_04875_),
    .A1(\top_ihp.oisc.regs[33][18] ));
 sg13g2_nand4_1 _22142_ (.B(_05683_),
    .C(_05684_),
    .A(_05682_),
    .Y(_05686_),
    .D(_05685_));
 sg13g2_or4_1 _22143_ (.A(_05672_),
    .B(_05677_),
    .C(_05681_),
    .D(_05686_),
    .X(_05687_));
 sg13g2_a22oi_1 _22144_ (.Y(_05688_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[43][18] ),
    .A2(net604),
    .A1(\top_ihp.oisc.regs[49][18] ));
 sg13g2_a22oi_1 _22145_ (.Y(_05689_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][18] ),
    .A2(net456),
    .A1(\top_ihp.oisc.regs[46][18] ));
 sg13g2_a22oi_1 _22146_ (.Y(_05690_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[45][18] ),
    .A2(net562),
    .A1(\top_ihp.oisc.regs[50][18] ));
 sg13g2_nand3_1 _22147_ (.B(net677),
    .C(net718),
    .A(\top_ihp.oisc.regs[31][18] ),
    .Y(_05691_));
 sg13g2_nand3_1 _22148_ (.B(net672),
    .C(_04722_),
    .A(\top_ihp.oisc.regs[17][18] ),
    .Y(_05692_));
 sg13g2_a21oi_1 _22149_ (.A1(_05691_),
    .A2(_05692_),
    .Y(_05693_),
    .B1(net696));
 sg13g2_a21oi_1 _22150_ (.A1(\top_ihp.oisc.regs[2][18] ),
    .A2(net600),
    .Y(_05694_),
    .B1(_05693_));
 sg13g2_nand4_1 _22151_ (.B(_05689_),
    .C(_05690_),
    .A(_05688_),
    .Y(_05695_),
    .D(_05694_));
 sg13g2_a22oi_1 _22152_ (.Y(_05696_),
    .B1(net419),
    .B2(\top_ihp.oisc.regs[5][18] ),
    .A2(_04902_),
    .A1(\top_ihp.oisc.regs[21][18] ));
 sg13g2_a22oi_1 _22153_ (.Y(_05697_),
    .B1(net466),
    .B2(\top_ihp.oisc.regs[1][18] ),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][18] ));
 sg13g2_a22oi_1 _22154_ (.Y(_05698_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][18] ),
    .A2(net617),
    .A1(\top_ihp.oisc.regs[7][18] ));
 sg13g2_a22oi_1 _22155_ (.Y(_05699_),
    .B1(_05154_),
    .B2(\top_ihp.oisc.regs[27][18] ),
    .A2(_05019_),
    .A1(\top_ihp.oisc.regs[11][18] ));
 sg13g2_nand4_1 _22156_ (.B(_05697_),
    .C(_05698_),
    .A(_05696_),
    .Y(_05700_),
    .D(_05699_));
 sg13g2_a22oi_1 _22157_ (.Y(_05701_),
    .B1(net581),
    .B2(\top_ihp.oisc.regs[51][18] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[32][18] ));
 sg13g2_nand2_1 _22158_ (.Y(_05702_),
    .A(\top_ihp.oisc.regs[30][18] ),
    .B(_05201_));
 sg13g2_and2_1 _22159_ (.A(net703),
    .B(net721),
    .X(_05703_));
 sg13g2_buf_1 _22160_ (.A(_05703_),
    .X(_05704_));
 sg13g2_buf_2 _22161_ (.A(_05704_),
    .X(_05705_));
 sg13g2_a22oi_1 _22162_ (.Y(_05706_),
    .B1(_05705_),
    .B2(\top_ihp.oisc.regs[22][18] ),
    .A2(net735),
    .A1(_07455_));
 sg13g2_buf_8 _22163_ (.A(_04999_),
    .X(_05707_));
 sg13g2_nand2_1 _22164_ (.Y(_05708_),
    .A(\top_ihp.oisc.regs[59][18] ),
    .B(net414));
 sg13g2_nand4_1 _22165_ (.B(_05702_),
    .C(_05706_),
    .A(_05701_),
    .Y(_05709_),
    .D(_05708_));
 sg13g2_nor4_1 _22166_ (.A(_05687_),
    .B(_05695_),
    .C(_05700_),
    .D(_05709_),
    .Y(_05710_));
 sg13g2_a21oi_1 _22167_ (.A1(_00125_),
    .A2(net77),
    .Y(_05711_),
    .B1(net153));
 sg13g2_a21oi_1 _22168_ (.A1(_07455_),
    .A2(net687),
    .Y(_05712_),
    .B1(_05711_));
 sg13g2_a21oi_1 _22169_ (.A1(_05664_),
    .A2(_05710_),
    .Y(_00303_),
    .B1(_05712_));
 sg13g2_a22oi_1 _22170_ (.Y(_05713_),
    .B1(net453),
    .B2(\top_ihp.oisc.regs[45][19] ),
    .A2(net261),
    .A1(\top_ihp.oisc.regs[44][19] ));
 sg13g2_a22oi_1 _22171_ (.Y(_05714_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[42][19] ),
    .A2(net469),
    .A1(\top_ihp.oisc.regs[5][19] ));
 sg13g2_a22oi_1 _22172_ (.Y(_05715_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[41][19] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[37][19] ));
 sg13g2_a22oi_1 _22173_ (.Y(_05716_),
    .B1(net591),
    .B2(\top_ihp.oisc.regs[52][19] ),
    .A2(net593),
    .A1(\top_ihp.oisc.regs[61][19] ));
 sg13g2_nand4_1 _22174_ (.B(_05714_),
    .C(_05715_),
    .A(_05713_),
    .Y(_05717_),
    .D(_05716_));
 sg13g2_a22oi_1 _22175_ (.Y(_05718_),
    .B1(_05467_),
    .B2(\top_ihp.oisc.regs[12][19] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][19] ));
 sg13g2_a22oi_1 _22176_ (.Y(_05719_),
    .B1(net466),
    .B2(\top_ihp.oisc.regs[1][19] ),
    .A2(_04902_),
    .A1(\top_ihp.oisc.regs[21][19] ));
 sg13g2_nor3_1 _22177_ (.A(_05025_),
    .B(net644),
    .C(net691),
    .Y(_05720_));
 sg13g2_a22oi_1 _22178_ (.Y(_05721_),
    .B1(_05720_),
    .B2(\top_ihp.oisc.regs[11][19] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][19] ));
 sg13g2_a22oi_1 _22179_ (.Y(_05722_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[9][19] ),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][19] ));
 sg13g2_nand4_1 _22180_ (.B(_05719_),
    .C(_05721_),
    .A(_05718_),
    .Y(_05723_),
    .D(_05722_));
 sg13g2_mux2_1 _22181_ (.A0(\top_ihp.oisc.regs[20][19] ),
    .A1(\top_ihp.oisc.regs[16][19] ),
    .S(net672),
    .X(_05724_));
 sg13g2_a22oi_1 _22182_ (.Y(_05725_),
    .B1(_05724_),
    .B2(net640),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][19] ));
 sg13g2_nand2b_1 _22183_ (.Y(_05726_),
    .B(net763),
    .A_N(_05725_));
 sg13g2_nor3_2 _22184_ (.A(net681),
    .B(net680),
    .C(net765),
    .Y(_05727_));
 sg13g2_mux2_1 _22185_ (.A0(\top_ihp.oisc.regs[6][19] ),
    .A1(\top_ihp.oisc.regs[2][19] ),
    .S(net652),
    .X(_05728_));
 sg13g2_a22oi_1 _22186_ (.Y(_05729_),
    .B1(_05727_),
    .B2(_05728_),
    .A2(_05345_),
    .A1(\top_ihp.oisc.regs[27][19] ));
 sg13g2_a22oi_1 _22187_ (.Y(_05730_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][19] ),
    .A2(_05342_),
    .A1(\top_ihp.oisc.regs[17][19] ));
 sg13g2_nand3_1 _22188_ (.B(_05729_),
    .C(_05730_),
    .A(_05726_),
    .Y(_05731_));
 sg13g2_nor4_1 _22189_ (.A(net76),
    .B(_05717_),
    .C(_05723_),
    .D(_05731_),
    .Y(_05732_));
 sg13g2_a22oi_1 _22190_ (.Y(_05733_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[43][19] ),
    .A2(net560),
    .A1(\top_ihp.oisc.regs[48][19] ));
 sg13g2_a22oi_1 _22191_ (.Y(_05734_),
    .B1(net454),
    .B2(\top_ihp.oisc.regs[34][19] ),
    .A2(net559),
    .A1(\top_ihp.oisc.regs[51][19] ));
 sg13g2_a22oi_1 _22192_ (.Y(_05735_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][19] ),
    .A2(net476),
    .A1(\top_ihp.oisc.regs[47][19] ));
 sg13g2_a22oi_1 _22193_ (.Y(_05736_),
    .B1(_04882_),
    .B2(\top_ihp.oisc.regs[4][19] ),
    .A2(_04880_),
    .A1(\top_ihp.oisc.regs[8][19] ));
 sg13g2_nor3_1 _22194_ (.A(net677),
    .B(net719),
    .C(_05736_),
    .Y(_05737_));
 sg13g2_a21oi_1 _22195_ (.A1(\top_ihp.oisc.regs[46][19] ),
    .A2(net456),
    .Y(_05738_),
    .B1(_05737_));
 sg13g2_nand4_1 _22196_ (.B(_05734_),
    .C(_05735_),
    .A(_05733_),
    .Y(_05739_),
    .D(_05738_));
 sg13g2_a22oi_1 _22197_ (.Y(_05740_),
    .B1(net436),
    .B2(\top_ihp.oisc.regs[33][19] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][19] ));
 sg13g2_a22oi_1 _22198_ (.Y(_05741_),
    .B1(net554),
    .B2(\top_ihp.oisc.regs[18][19] ),
    .A2(_05202_),
    .A1(net1042));
 sg13g2_inv_1 _22199_ (.Y(_05742_),
    .A(_05741_));
 sg13g2_a221oi_1 _22200_ (.B2(\top_ihp.oisc.regs[22][19] ),
    .C1(_05742_),
    .B1(net552),
    .A1(\top_ihp.oisc.regs[36][19] ),
    .Y(_05743_),
    .A2(net462));
 sg13g2_a22oi_1 _22201_ (.Y(_05744_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[15][19] ),
    .A2(net657),
    .A1(\top_ihp.oisc.regs[7][19] ));
 sg13g2_a22oi_1 _22202_ (.Y(_05745_),
    .B1(net573),
    .B2(\top_ihp.oisc.regs[31][19] ),
    .A2(_04898_),
    .A1(\top_ihp.oisc.regs[10][19] ));
 sg13g2_mux2_1 _22203_ (.A0(\top_ihp.oisc.regs[3][19] ),
    .A1(\top_ihp.oisc.regs[19][19] ),
    .S(net725),
    .X(_05746_));
 sg13g2_a22oi_1 _22204_ (.Y(_05747_),
    .B1(_04957_),
    .B2(_05746_),
    .A2(net613),
    .A1(\top_ihp.oisc.regs[29][19] ));
 sg13g2_mux2_1 _22205_ (.A0(\top_ihp.oisc.regs[30][19] ),
    .A1(\top_ihp.oisc.regs[26][19] ),
    .S(net666),
    .X(_05748_));
 sg13g2_a22oi_1 _22206_ (.Y(_05749_),
    .B1(_04930_),
    .B2(_05748_),
    .A2(net655),
    .A1(\top_ihp.oisc.regs[13][19] ));
 sg13g2_and4_1 _22207_ (.A(_05744_),
    .B(_05745_),
    .C(_05747_),
    .D(_05749_),
    .X(_05750_));
 sg13g2_nand3_1 _22208_ (.B(_05743_),
    .C(_05750_),
    .A(_05740_),
    .Y(_05751_));
 sg13g2_a22oi_1 _22209_ (.Y(_05752_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[59][19] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][19] ));
 sg13g2_a22oi_1 _22210_ (.Y(_05753_),
    .B1(net452),
    .B2(\top_ihp.oisc.regs[39][19] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][19] ));
 sg13g2_a22oi_1 _22211_ (.Y(_05754_),
    .B1(net457),
    .B2(\top_ihp.oisc.regs[35][19] ),
    .A2(net582),
    .A1(\top_ihp.oisc.regs[62][19] ));
 sg13g2_a22oi_1 _22212_ (.Y(_05755_),
    .B1(net578),
    .B2(\top_ihp.oisc.regs[50][19] ),
    .A2(net596),
    .A1(\top_ihp.oisc.regs[63][19] ));
 sg13g2_nand4_1 _22213_ (.B(_05753_),
    .C(_05754_),
    .A(_05752_),
    .Y(_05756_),
    .D(_05755_));
 sg13g2_nand2_1 _22214_ (.Y(_05757_),
    .A(\top_ihp.oisc.regs[58][19] ),
    .B(net442));
 sg13g2_buf_8 _22215_ (.A(net459),
    .X(_05758_));
 sg13g2_a22oi_1 _22216_ (.Y(_05759_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][19] ),
    .A2(net255),
    .A1(\top_ihp.oisc.regs[56][19] ));
 sg13g2_buf_8 _22217_ (.A(net570),
    .X(_05760_));
 sg13g2_a22oi_1 _22218_ (.Y(_05761_),
    .B1(net413),
    .B2(\top_ihp.oisc.regs[57][19] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[49][19] ));
 sg13g2_a22oi_1 _22219_ (.Y(_05762_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[54][19] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[32][19] ));
 sg13g2_nand4_1 _22220_ (.B(_05759_),
    .C(_05761_),
    .A(_05757_),
    .Y(_05763_),
    .D(_05762_));
 sg13g2_nor4_1 _22221_ (.A(_05739_),
    .B(_05751_),
    .C(_05756_),
    .D(_05763_),
    .Y(_05764_));
 sg13g2_a21oi_1 _22222_ (.A1(_00126_),
    .A2(net77),
    .Y(_05765_),
    .B1(net153));
 sg13g2_a21oi_1 _22223_ (.A1(_07459_),
    .A2(net687),
    .Y(_05766_),
    .B1(_05765_));
 sg13g2_a21oi_1 _22224_ (.A1(_05732_),
    .A2(_05764_),
    .Y(_00304_),
    .B1(_05766_));
 sg13g2_nand2_1 _22225_ (.Y(_05767_),
    .A(net1041),
    .B(_03688_));
 sg13g2_a21o_1 _22226_ (.A2(net76),
    .A1(_00108_),
    .B1(net154),
    .X(_05768_));
 sg13g2_a22oi_1 _22227_ (.Y(_05769_),
    .B1(net581),
    .B2(\top_ihp.oisc.regs[51][1] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][1] ));
 sg13g2_a22oi_1 _22228_ (.Y(_05770_),
    .B1(net579),
    .B2(\top_ihp.oisc.regs[48][1] ),
    .A2(_04909_),
    .A1(\top_ihp.oisc.regs[5][1] ));
 sg13g2_a22oi_1 _22229_ (.Y(_05771_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][1] ),
    .A2(net567),
    .A1(\top_ihp.oisc.regs[61][1] ));
 sg13g2_a22oi_1 _22230_ (.Y(_05772_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][1] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][1] ));
 sg13g2_nand4_1 _22231_ (.B(_05770_),
    .C(_05771_),
    .A(_05769_),
    .Y(_05773_),
    .D(_05772_));
 sg13g2_a22oi_1 _22232_ (.Y(_05774_),
    .B1(_05273_),
    .B2(\top_ihp.oisc.regs[12][1] ),
    .A2(_05007_),
    .A1(\top_ihp.oisc.regs[2][1] ));
 sg13g2_mux2_1 _22233_ (.A0(\top_ihp.oisc.regs[24][1] ),
    .A1(\top_ihp.oisc.regs[16][1] ),
    .S(net667),
    .X(_05775_));
 sg13g2_a22oi_1 _22234_ (.Y(_05776_),
    .B1(_05775_),
    .B2(net556),
    .A2(net557),
    .A1(\top_ihp.oisc.regs[20][1] ));
 sg13g2_nand2b_1 _22235_ (.Y(_05777_),
    .B(net763),
    .A_N(_05776_));
 sg13g2_o21ai_1 _22236_ (.B1(_05777_),
    .Y(_05778_),
    .A1(_05272_),
    .A2(_05774_));
 sg13g2_a22oi_1 _22237_ (.Y(_05779_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][1] ),
    .A2(net468),
    .A1(\top_ihp.oisc.regs[6][1] ));
 sg13g2_a22oi_1 _22238_ (.Y(_05780_),
    .B1(net465),
    .B2(\top_ihp.oisc.regs[31][1] ),
    .A2(net472),
    .A1(\top_ihp.oisc.regs[29][1] ));
 sg13g2_a22oi_1 _22239_ (.Y(_05781_),
    .B1(net464),
    .B2(\top_ihp.oisc.regs[28][1] ),
    .A2(net473),
    .A1(\top_ihp.oisc.regs[13][1] ));
 sg13g2_a22oi_1 _22240_ (.Y(_05782_),
    .B1(net467),
    .B2(\top_ihp.oisc.regs[15][1] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][1] ));
 sg13g2_nand4_1 _22241_ (.B(_05780_),
    .C(_05781_),
    .A(_05779_),
    .Y(_05783_),
    .D(_05782_));
 sg13g2_nor4_1 _22242_ (.A(net79),
    .B(_05773_),
    .C(_05778_),
    .D(_05783_),
    .Y(_05784_));
 sg13g2_a22oi_1 _22243_ (.Y(_05785_),
    .B1(_05760_),
    .B2(\top_ihp.oisc.regs[57][1] ),
    .A2(net255),
    .A1(\top_ihp.oisc.regs[56][1] ));
 sg13g2_a22oi_1 _22244_ (.Y(_05786_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[58][1] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][1] ));
 sg13g2_a22oi_1 _22245_ (.Y(_05787_),
    .B1(net455),
    .B2(\top_ihp.oisc.regs[52][1] ),
    .A2(net562),
    .A1(\top_ihp.oisc.regs[50][1] ));
 sg13g2_a22oi_1 _22246_ (.Y(_05788_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][1] ),
    .A2(net582),
    .A1(\top_ihp.oisc.regs[62][1] ));
 sg13g2_nand4_1 _22247_ (.B(_05786_),
    .C(_05787_),
    .A(_05785_),
    .Y(_05789_),
    .D(_05788_));
 sg13g2_a22oi_1 _22248_ (.Y(_05790_),
    .B1(net577),
    .B2(\top_ihp.oisc.regs[4][1] ),
    .A2(_05329_),
    .A1(\top_ihp.oisc.regs[1][1] ));
 sg13g2_a22oi_1 _22249_ (.Y(_05791_),
    .B1(_05255_),
    .B2(\top_ihp.oisc.regs[8][1] ),
    .A2(_05022_),
    .A1(\top_ihp.oisc.regs[9][1] ));
 sg13g2_mux2_1 _22250_ (.A0(\top_ihp.oisc.regs[3][1] ),
    .A1(\top_ihp.oisc.regs[19][1] ),
    .S(net693),
    .X(_05792_));
 sg13g2_a22oi_1 _22251_ (.Y(_05793_),
    .B1(net692),
    .B2(_05792_),
    .A2(_05158_),
    .A1(\top_ihp.oisc.regs[21][1] ));
 sg13g2_a22oi_1 _22252_ (.Y(_05794_),
    .B1(net561),
    .B2(\top_ihp.oisc.regs[27][1] ),
    .A2(net618),
    .A1(\top_ihp.oisc.regs[17][1] ));
 sg13g2_nand4_1 _22253_ (.B(_05791_),
    .C(_05793_),
    .A(_05790_),
    .Y(_05795_),
    .D(_05794_));
 sg13g2_a22oi_1 _22254_ (.Y(_05796_),
    .B1(_05142_),
    .B2(\top_ihp.oisc.regs[23][1] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][1] ));
 sg13g2_a22oi_1 _22255_ (.Y(_05797_),
    .B1(net471),
    .B2(\top_ihp.oisc.regs[10][1] ),
    .A2(net477),
    .A1(\top_ihp.oisc.regs[14][1] ));
 sg13g2_nand2_1 _22256_ (.Y(_05798_),
    .A(\top_ihp.oisc.regs[40][1] ),
    .B(net451));
 sg13g2_a22oi_1 _22257_ (.Y(_05799_),
    .B1(net720),
    .B2(\top_ihp.oisc.regs[26][1] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[18][1] ));
 sg13g2_o21ai_1 _22258_ (.B1(_05767_),
    .Y(_05800_),
    .A1(net669),
    .A2(_05799_));
 sg13g2_a221oi_1 _22259_ (.B2(\top_ihp.oisc.regs[22][1] ),
    .C1(_05800_),
    .B1(net552),
    .A1(\top_ihp.oisc.regs[30][1] ),
    .Y(_05801_),
    .A2(net646));
 sg13g2_nand4_1 _22260_ (.B(_05797_),
    .C(_05798_),
    .A(_05796_),
    .Y(_05802_),
    .D(_05801_));
 sg13g2_or2_1 _22261_ (.X(_05803_),
    .B(_05802_),
    .A(_05795_));
 sg13g2_a22oi_1 _22262_ (.Y(_05804_),
    .B1(net268),
    .B2(\top_ihp.oisc.regs[44][1] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][1] ));
 sg13g2_a22oi_1 _22263_ (.Y(_05805_),
    .B1(net270),
    .B2(\top_ihp.oisc.regs[46][1] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[35][1] ));
 sg13g2_a22oi_1 _22264_ (.Y(_05806_),
    .B1(net417),
    .B2(\top_ihp.oisc.regs[49][1] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[32][1] ));
 sg13g2_a22oi_1 _22265_ (.Y(_05807_),
    .B1(net436),
    .B2(\top_ihp.oisc.regs[33][1] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][1] ));
 sg13g2_nand4_1 _22266_ (.B(_05805_),
    .C(_05806_),
    .A(_05804_),
    .Y(_05808_),
    .D(_05807_));
 sg13g2_a22oi_1 _22267_ (.Y(_05809_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][1] ),
    .A2(net272),
    .A1(\top_ihp.oisc.regs[34][1] ));
 sg13g2_a22oi_1 _22268_ (.Y(_05810_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][1] ),
    .A2(net262),
    .A1(\top_ihp.oisc.regs[36][1] ));
 sg13g2_a22oi_1 _22269_ (.Y(_05811_),
    .B1(_05110_),
    .B2(\top_ihp.oisc.regs[43][1] ),
    .A2(net267),
    .A1(\top_ihp.oisc.regs[38][1] ));
 sg13g2_a22oi_1 _22270_ (.Y(_05812_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[63][1] ),
    .A2(net568),
    .A1(\top_ihp.oisc.regs[59][1] ));
 sg13g2_nand4_1 _22271_ (.B(_05810_),
    .C(_05811_),
    .A(_05809_),
    .Y(_05813_),
    .D(_05812_));
 sg13g2_nor4_2 _22272_ (.A(_05789_),
    .B(_05803_),
    .C(_05808_),
    .Y(_05814_),
    .D(_05813_));
 sg13g2_a22oi_1 _22273_ (.Y(_00305_),
    .B1(_05784_),
    .B2(_05814_),
    .A2(_05768_),
    .A1(_05767_));
 sg13g2_mux2_1 _22274_ (.A0(\top_ihp.oisc.regs[28][20] ),
    .A1(\top_ihp.oisc.regs[20][20] ),
    .S(net670),
    .X(_05815_));
 sg13g2_a22oi_1 _22275_ (.Y(_05816_),
    .B1(_05815_),
    .B2(net669),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[24][20] ));
 sg13g2_a22oi_1 _22276_ (.Y(_05817_),
    .B1(_05076_),
    .B2(\top_ihp.oisc.regs[45][20] ),
    .A2(_05011_),
    .A1(\top_ihp.oisc.regs[51][20] ));
 sg13g2_o21ai_1 _22277_ (.B1(_05817_),
    .Y(_05818_),
    .A1(net689),
    .A2(_05816_));
 sg13g2_a22oi_1 _22278_ (.Y(_05819_),
    .B1(_04826_),
    .B2(\top_ihp.oisc.regs[14][20] ),
    .A2(_05144_),
    .A1(\top_ihp.oisc.regs[17][20] ));
 sg13g2_a22oi_1 _22279_ (.Y(_05820_),
    .B1(net655),
    .B2(\top_ihp.oisc.regs[13][20] ),
    .A2(net657),
    .A1(\top_ihp.oisc.regs[7][20] ));
 sg13g2_a22oi_1 _22280_ (.Y(_05821_),
    .B1(_05254_),
    .B2(\top_ihp.oisc.regs[8][20] ),
    .A2(_04951_),
    .A1(\top_ihp.oisc.regs[16][20] ));
 sg13g2_a22oi_1 _22281_ (.Y(_05822_),
    .B1(_05150_),
    .B2(\top_ihp.oisc.regs[12][20] ),
    .A2(net647),
    .A1(\top_ihp.oisc.regs[11][20] ));
 sg13g2_nand4_1 _22282_ (.B(_05820_),
    .C(_05821_),
    .A(_05819_),
    .Y(_05823_),
    .D(_05822_));
 sg13g2_mux2_1 _22283_ (.A0(\top_ihp.oisc.regs[3][20] ),
    .A1(\top_ihp.oisc.regs[19][20] ),
    .S(net725),
    .X(_05824_));
 sg13g2_a22oi_1 _22284_ (.Y(_05825_),
    .B1(_05824_),
    .B2(_04957_),
    .A2(net648),
    .A1(\top_ihp.oisc.regs[23][20] ));
 sg13g2_a22oi_1 _22285_ (.Y(_05826_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[15][20] ),
    .A2(_04817_),
    .A1(\top_ihp.oisc.regs[25][20] ));
 sg13g2_mux2_1 _22286_ (.A0(\top_ihp.oisc.regs[22][20] ),
    .A1(\top_ihp.oisc.regs[18][20] ),
    .S(net666),
    .X(_05827_));
 sg13g2_a22oi_1 _22287_ (.Y(_05828_),
    .B1(_05827_),
    .B2(net695),
    .A2(net561),
    .A1(\top_ihp.oisc.regs[27][20] ));
 sg13g2_mux2_1 _22288_ (.A0(\top_ihp.oisc.regs[30][20] ),
    .A1(\top_ihp.oisc.regs[26][20] ),
    .S(net666),
    .X(_05829_));
 sg13g2_a22oi_1 _22289_ (.Y(_05830_),
    .B1(net720),
    .B2(_05829_),
    .A2(_04907_),
    .A1(\top_ihp.oisc.regs[5][20] ));
 sg13g2_nand4_1 _22290_ (.B(_05826_),
    .C(_05828_),
    .A(_05825_),
    .Y(_05831_),
    .D(_05830_));
 sg13g2_nand2_1 _22291_ (.Y(_05832_),
    .A(\top_ihp.oisc.regs[58][20] ),
    .B(net603));
 sg13g2_a22oi_1 _22292_ (.Y(_05833_),
    .B1(_05329_),
    .B2(\top_ihp.oisc.regs[1][20] ),
    .A2(net772),
    .A1(_07450_));
 sg13g2_a22oi_1 _22293_ (.Y(_05834_),
    .B1(net573),
    .B2(\top_ihp.oisc.regs[31][20] ),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][20] ));
 sg13g2_a22oi_1 _22294_ (.Y(_05835_),
    .B1(net597),
    .B2(\top_ihp.oisc.regs[9][20] ),
    .A2(_04893_),
    .A1(\top_ihp.oisc.regs[29][20] ));
 sg13g2_nand4_1 _22295_ (.B(_05833_),
    .C(_05834_),
    .A(_05832_),
    .Y(_05836_),
    .D(_05835_));
 sg13g2_or4_1 _22296_ (.A(_05818_),
    .B(_05823_),
    .C(_05831_),
    .D(_05836_),
    .X(_05837_));
 sg13g2_a22oi_1 _22297_ (.Y(_05838_),
    .B1(_05114_),
    .B2(\top_ihp.oisc.regs[44][20] ),
    .A2(_05040_),
    .A1(\top_ihp.oisc.regs[50][20] ));
 sg13g2_a22oi_1 _22298_ (.Y(_05839_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][20] ),
    .A2(net262),
    .A1(\top_ihp.oisc.regs[36][20] ));
 sg13g2_a22oi_1 _22299_ (.Y(_05840_),
    .B1(net601),
    .B2(\top_ihp.oisc.regs[48][20] ),
    .A2(net425),
    .A1(\top_ihp.oisc.regs[42][20] ));
 sg13g2_a22oi_1 _22300_ (.Y(_05841_),
    .B1(net436),
    .B2(\top_ihp.oisc.regs[33][20] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][20] ));
 sg13g2_nand4_1 _22301_ (.B(_05839_),
    .C(_05840_),
    .A(_05838_),
    .Y(_05842_),
    .D(_05841_));
 sg13g2_a22oi_1 _22302_ (.Y(_05843_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[52][20] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[57][20] ));
 sg13g2_a22oi_1 _22303_ (.Y(_05844_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][20] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[62][20] ));
 sg13g2_a22oi_1 _22304_ (.Y(_05845_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][20] ),
    .A2(net255),
    .A1(\top_ihp.oisc.regs[56][20] ));
 sg13g2_a22oi_1 _22305_ (.Y(_05846_),
    .B1(net557),
    .B2(\top_ihp.oisc.regs[6][20] ),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[10][20] ));
 sg13g2_nor2_1 _22306_ (.A(_04799_),
    .B(_05846_),
    .Y(_05847_));
 sg13g2_a21oi_1 _22307_ (.A1(\top_ihp.oisc.regs[63][20] ),
    .A2(net439),
    .Y(_05848_),
    .B1(_05847_));
 sg13g2_nand4_1 _22308_ (.B(_05844_),
    .C(_05845_),
    .A(_05843_),
    .Y(_05849_),
    .D(_05848_));
 sg13g2_nor3_1 _22309_ (.A(_05837_),
    .B(_05842_),
    .C(_05849_),
    .Y(_05850_));
 sg13g2_a22oi_1 _22310_ (.Y(_05851_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][20] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[39][20] ));
 sg13g2_a22oi_1 _22311_ (.Y(_05852_),
    .B1(net270),
    .B2(\top_ihp.oisc.regs[46][20] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[32][20] ));
 sg13g2_a22oi_1 _22312_ (.Y(_05853_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][20] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][20] ));
 sg13g2_a22oi_1 _22313_ (.Y(_05854_),
    .B1(_05110_),
    .B2(\top_ihp.oisc.regs[43][20] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[49][20] ));
 sg13g2_nand4_1 _22314_ (.B(_05852_),
    .C(_05853_),
    .A(_05851_),
    .Y(_05855_),
    .D(_05854_));
 sg13g2_a22oi_1 _22315_ (.Y(_05856_),
    .B1(_04765_),
    .B2(\top_ihp.oisc.regs[4][20] ),
    .A2(_04763_),
    .A1(\top_ihp.oisc.regs[2][20] ));
 sg13g2_nor3_1 _22316_ (.A(net643),
    .B(net719),
    .C(_05856_),
    .Y(_05857_));
 sg13g2_a221oi_1 _22317_ (.B2(\top_ihp.oisc.regs[35][20] ),
    .C1(_05857_),
    .B1(net420),
    .A1(\top_ihp.oisc.regs[54][20] ),
    .Y(_05858_),
    .A2(net606));
 sg13g2_a22oi_1 _22318_ (.Y(_05859_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][20] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][20] ));
 sg13g2_a22oi_1 _22319_ (.Y(_05860_),
    .B1(_05707_),
    .B2(\top_ihp.oisc.regs[59][20] ),
    .A2(_05170_),
    .A1(\top_ihp.oisc.regs[38][20] ));
 sg13g2_nand3_1 _22320_ (.B(_05859_),
    .C(_05860_),
    .A(_05858_),
    .Y(_05861_));
 sg13g2_nor3_1 _22321_ (.A(_05101_),
    .B(_05855_),
    .C(_05861_),
    .Y(_05862_));
 sg13g2_a21oi_1 _22322_ (.A1(_00127_),
    .A2(net77),
    .Y(_05863_),
    .B1(net153));
 sg13g2_a21oi_1 _22323_ (.A1(_07450_),
    .A2(net687),
    .Y(_05864_),
    .B1(_05863_));
 sg13g2_a21oi_1 _22324_ (.A1(_05850_),
    .A2(_05862_),
    .Y(_00306_),
    .B1(_05864_));
 sg13g2_a22oi_1 _22325_ (.Y(_05865_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][21] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][21] ));
 sg13g2_a22oi_1 _22326_ (.Y(_05866_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][21] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][21] ));
 sg13g2_a22oi_1 _22327_ (.Y(_05867_),
    .B1(net578),
    .B2(\top_ihp.oisc.regs[50][21] ),
    .A2(net563),
    .A1(\top_ihp.oisc.regs[49][21] ));
 sg13g2_a22oi_1 _22328_ (.Y(_05868_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[38][21] ),
    .A2(net615),
    .A1(\top_ihp.oisc.regs[55][21] ));
 sg13g2_nand4_1 _22329_ (.B(_05866_),
    .C(_05867_),
    .A(_05865_),
    .Y(_05869_),
    .D(_05868_));
 sg13g2_and2_1 _22330_ (.A(\top_ihp.oisc.regs[45][21] ),
    .B(_05076_),
    .X(_05870_));
 sg13g2_a221oi_1 _22331_ (.B2(\top_ihp.oisc.regs[39][21] ),
    .C1(_05870_),
    .B1(net445),
    .A1(\top_ihp.oisc.regs[61][21] ),
    .Y(_05871_),
    .A2(net593));
 sg13g2_a22oi_1 _22332_ (.Y(_05872_),
    .B1(net579),
    .B2(\top_ihp.oisc.regs[48][21] ),
    .A2(net606),
    .A1(\top_ihp.oisc.regs[54][21] ));
 sg13g2_a22oi_1 _22333_ (.Y(_05873_),
    .B1(net608),
    .B2(\top_ihp.oisc.regs[1][21] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][21] ));
 sg13g2_a22oi_1 _22334_ (.Y(_05874_),
    .B1(_04940_),
    .B2(\top_ihp.oisc.regs[31][21] ),
    .A2(net612),
    .A1(\top_ihp.oisc.regs[21][21] ));
 sg13g2_nand4_1 _22335_ (.B(_05872_),
    .C(_05873_),
    .A(_05871_),
    .Y(_05875_),
    .D(_05874_));
 sg13g2_a22oi_1 _22336_ (.Y(_05876_),
    .B1(_05760_),
    .B2(\top_ihp.oisc.regs[57][21] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[2][21] ));
 sg13g2_a22oi_1 _22337_ (.Y(_05877_),
    .B1(net594),
    .B2(\top_ihp.oisc.regs[62][21] ),
    .A2(net261),
    .A1(\top_ihp.oisc.regs[44][21] ));
 sg13g2_a22oi_1 _22338_ (.Y(_05878_),
    .B1(net455),
    .B2(\top_ihp.oisc.regs[52][21] ),
    .A2(_05264_),
    .A1(\top_ihp.oisc.regs[53][21] ));
 sg13g2_a22oi_1 _22339_ (.Y(_05879_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][21] ),
    .A2(_04999_),
    .A1(\top_ihp.oisc.regs[59][21] ));
 sg13g2_nand4_1 _22340_ (.B(_05877_),
    .C(_05878_),
    .A(_05876_),
    .Y(_05880_),
    .D(_05879_));
 sg13g2_a22oi_1 _22341_ (.Y(_05881_),
    .B1(net269),
    .B2(\top_ihp.oisc.regs[43][21] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[33][21] ));
 sg13g2_a22oi_1 _22342_ (.Y(_05882_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[35][21] ),
    .A2(net442),
    .A1(\top_ihp.oisc.regs[58][21] ));
 sg13g2_a22oi_1 _22343_ (.Y(_05883_),
    .B1(net581),
    .B2(\top_ihp.oisc.regs[51][21] ),
    .A2(net425),
    .A1(\top_ihp.oisc.regs[42][21] ));
 sg13g2_a22oi_1 _22344_ (.Y(_05884_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][21] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[46][21] ));
 sg13g2_nand4_1 _22345_ (.B(_05882_),
    .C(_05883_),
    .A(_05881_),
    .Y(_05885_),
    .D(_05884_));
 sg13g2_nor4_2 _22346_ (.A(_05869_),
    .B(_05875_),
    .C(_05880_),
    .Y(_05886_),
    .D(_05885_));
 sg13g2_and2_1 _22347_ (.A(_07461_),
    .B(_03689_),
    .X(_05887_));
 sg13g2_a221oi_1 _22348_ (.B2(\top_ihp.oisc.regs[3][21] ),
    .C1(_05887_),
    .B1(_05245_),
    .A1(\top_ihp.oisc.regs[19][21] ),
    .Y(_05888_),
    .A2(_05241_));
 sg13g2_a22oi_1 _22349_ (.Y(_05889_),
    .B1(_05254_),
    .B2(\top_ihp.oisc.regs[8][21] ),
    .A2(_04888_),
    .A1(\top_ihp.oisc.regs[13][21] ));
 sg13g2_mux2_1 _22350_ (.A0(\top_ihp.oisc.regs[30][21] ),
    .A1(\top_ihp.oisc.regs[26][21] ),
    .S(_05326_),
    .X(_05890_));
 sg13g2_a22oi_1 _22351_ (.Y(_05891_),
    .B1(net720),
    .B2(_05890_),
    .A2(net653),
    .A1(\top_ihp.oisc.regs[15][21] ));
 sg13g2_a22oi_1 _22352_ (.Y(_05892_),
    .B1(_05146_),
    .B2(\top_ihp.oisc.regs[11][21] ),
    .A2(_04833_),
    .A1(\top_ihp.oisc.regs[24][21] ));
 sg13g2_and4_1 _22353_ (.A(_05888_),
    .B(_05889_),
    .C(_05891_),
    .D(_05892_),
    .X(_05893_));
 sg13g2_a22oi_1 _22354_ (.Y(_05894_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[63][21] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[36][21] ));
 sg13g2_a22oi_1 _22355_ (.Y(_05895_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][21] ),
    .A2(net459),
    .A1(\top_ihp.oisc.regs[56][21] ));
 sg13g2_nand3_1 _22356_ (.B(_05894_),
    .C(_05895_),
    .A(_05893_),
    .Y(_05896_));
 sg13g2_mux2_1 _22357_ (.A0(\top_ihp.oisc.regs[20][21] ),
    .A1(\top_ihp.oisc.regs[16][21] ),
    .S(net654),
    .X(_05897_));
 sg13g2_a22oi_1 _22358_ (.Y(_05898_),
    .B1(_05897_),
    .B2(_04853_),
    .A2(net617),
    .A1(\top_ihp.oisc.regs[7][21] ));
 sg13g2_a22oi_1 _22359_ (.Y(_05899_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][21] ),
    .A2(net569),
    .A1(\top_ihp.oisc.regs[9][21] ));
 sg13g2_a22oi_1 _22360_ (.Y(_05900_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][21] ),
    .A2(_05016_),
    .A1(\top_ihp.oisc.regs[4][21] ));
 sg13g2_a22oi_1 _22361_ (.Y(_05901_),
    .B1(net555),
    .B2(\top_ihp.oisc.regs[29][21] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[17][21] ));
 sg13g2_nand4_1 _22362_ (.B(_05899_),
    .C(_05900_),
    .A(_05898_),
    .Y(_05902_),
    .D(_05901_));
 sg13g2_a22oi_1 _22363_ (.Y(_05903_),
    .B1(net468),
    .B2(\top_ihp.oisc.regs[6][21] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[5][21] ));
 sg13g2_mux2_1 _22364_ (.A0(\top_ihp.oisc.regs[22][21] ),
    .A1(\top_ihp.oisc.regs[18][21] ),
    .S(net652),
    .X(_05904_));
 sg13g2_nand2_1 _22365_ (.Y(_05905_),
    .A(net695),
    .B(_05904_));
 sg13g2_a22oi_1 _22366_ (.Y(_05906_),
    .B1(net464),
    .B2(\top_ihp.oisc.regs[28][21] ),
    .A2(net257),
    .A1(\top_ihp.oisc.regs[10][21] ));
 sg13g2_a22oi_1 _22367_ (.Y(_05907_),
    .B1(_05345_),
    .B2(\top_ihp.oisc.regs[27][21] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][21] ));
 sg13g2_nand4_1 _22368_ (.B(_05905_),
    .C(_05906_),
    .A(_05903_),
    .Y(_05908_),
    .D(_05907_));
 sg13g2_nor4_1 _22369_ (.A(net80),
    .B(_05896_),
    .C(_05902_),
    .D(_05908_),
    .Y(_05909_));
 sg13g2_a21oi_1 _22370_ (.A1(_00128_),
    .A2(net78),
    .Y(_05910_),
    .B1(_05105_));
 sg13g2_nor2_1 _22371_ (.A(_05887_),
    .B(_05910_),
    .Y(_05911_));
 sg13g2_a21oi_1 _22372_ (.A1(_05886_),
    .A2(_05909_),
    .Y(_00307_),
    .B1(_05911_));
 sg13g2_a22oi_1 _22373_ (.Y(_05912_),
    .B1(_05183_),
    .B2(\top_ihp.oisc.regs[48][22] ),
    .A2(net606),
    .A1(\top_ihp.oisc.regs[54][22] ));
 sg13g2_a22oi_1 _22374_ (.Y(_05913_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][22] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[37][22] ));
 sg13g2_a22oi_1 _22375_ (.Y(_05914_),
    .B1(net591),
    .B2(\top_ihp.oisc.regs[52][22] ),
    .A2(_05052_),
    .A1(\top_ihp.oisc.regs[61][22] ));
 sg13g2_a22oi_1 _22376_ (.Y(_05915_),
    .B1(_05055_),
    .B2(\top_ihp.oisc.regs[35][22] ),
    .A2(net562),
    .A1(\top_ihp.oisc.regs[50][22] ));
 sg13g2_nand4_1 _22377_ (.B(_05913_),
    .C(_05914_),
    .A(_05912_),
    .Y(_05916_),
    .D(_05915_));
 sg13g2_inv_1 _22378_ (.Y(_05917_),
    .A(\top_ihp.oisc.regs[6][22] ));
 sg13g2_nor2_1 _22379_ (.A(_05917_),
    .B(_04772_),
    .Y(_05918_));
 sg13g2_a22oi_1 _22380_ (.Y(_05919_),
    .B1(net674),
    .B2(_05918_),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][22] ));
 sg13g2_a22oi_1 _22381_ (.Y(_05920_),
    .B1(_05150_),
    .B2(\top_ihp.oisc.regs[12][22] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][22] ));
 sg13g2_mux2_1 _22382_ (.A0(\top_ihp.oisc.regs[3][22] ),
    .A1(\top_ihp.oisc.regs[19][22] ),
    .S(net725),
    .X(_05921_));
 sg13g2_a22oi_1 _22383_ (.Y(_05922_),
    .B1(_04957_),
    .B2(_05921_),
    .A2(net655),
    .A1(\top_ihp.oisc.regs[13][22] ));
 sg13g2_a22oi_1 _22384_ (.Y(_05923_),
    .B1(net561),
    .B2(\top_ihp.oisc.regs[27][22] ),
    .A2(_05146_),
    .A1(\top_ihp.oisc.regs[11][22] ));
 sg13g2_and4_1 _22385_ (.A(_05919_),
    .B(_05920_),
    .C(_05922_),
    .D(_05923_),
    .X(_05924_));
 sg13g2_a22oi_1 _22386_ (.Y(_05925_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][22] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[46][22] ));
 sg13g2_a22oi_1 _22387_ (.Y(_05926_),
    .B1(_05224_),
    .B2(\top_ihp.oisc.regs[36][22] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][22] ));
 sg13g2_nand3_1 _22388_ (.B(_05925_),
    .C(_05926_),
    .A(_05924_),
    .Y(_05927_));
 sg13g2_a22oi_1 _22389_ (.Y(_05928_),
    .B1(net553),
    .B2(\top_ihp.oisc.regs[62][22] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][22] ));
 sg13g2_a22oi_1 _22390_ (.Y(_05929_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[42][22] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[32][22] ));
 sg13g2_a22oi_1 _22391_ (.Y(_05930_),
    .B1(net453),
    .B2(\top_ihp.oisc.regs[45][22] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][22] ));
 sg13g2_a22oi_1 _22392_ (.Y(_05931_),
    .B1(net261),
    .B2(\top_ihp.oisc.regs[44][22] ),
    .A2(net459),
    .A1(\top_ihp.oisc.regs[56][22] ));
 sg13g2_nand4_1 _22393_ (.B(_05929_),
    .C(_05930_),
    .A(_05928_),
    .Y(_05932_),
    .D(_05931_));
 sg13g2_a22oi_1 _22394_ (.Y(_05933_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][22] ),
    .A2(net439),
    .A1(\top_ihp.oisc.regs[63][22] ));
 sg13g2_a22oi_1 _22395_ (.Y(_05934_),
    .B1(_05707_),
    .B2(\top_ihp.oisc.regs[59][22] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][22] ));
 sg13g2_a22oi_1 _22396_ (.Y(_05935_),
    .B1(_05170_),
    .B2(\top_ihp.oisc.regs[38][22] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][22] ));
 sg13g2_a22oi_1 _22397_ (.Y(_05936_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][22] ),
    .A2(_05590_),
    .A1(\top_ihp.oisc.regs[49][22] ));
 sg13g2_nand4_1 _22398_ (.B(_05934_),
    .C(_05935_),
    .A(_05933_),
    .Y(_05937_),
    .D(_05936_));
 sg13g2_nor4_1 _22399_ (.A(_05916_),
    .B(_05927_),
    .C(_05932_),
    .D(_05937_),
    .Y(_05938_));
 sg13g2_mux2_1 _22400_ (.A0(\top_ihp.oisc.regs[22][22] ),
    .A1(\top_ihp.oisc.regs[18][22] ),
    .S(net654),
    .X(_05939_));
 sg13g2_a22oi_1 _22401_ (.Y(_05940_),
    .B1(_05939_),
    .B2(net695),
    .A2(net433),
    .A1(\top_ihp.oisc.regs[8][22] ));
 sg13g2_a22oi_1 _22402_ (.Y(_05941_),
    .B1(_04899_),
    .B2(\top_ihp.oisc.regs[10][22] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][22] ));
 sg13g2_a22oi_1 _22403_ (.Y(_05942_),
    .B1(net598),
    .B2(\top_ihp.oisc.regs[4][22] ),
    .A2(_04936_),
    .A1(\top_ihp.oisc.regs[1][22] ));
 sg13g2_a22oi_1 _22404_ (.Y(_05943_),
    .B1(net607),
    .B2(\top_ihp.oisc.regs[31][22] ),
    .A2(_04821_),
    .A1(\top_ihp.oisc.regs[17][22] ));
 sg13g2_nand4_1 _22405_ (.B(_05941_),
    .C(_05942_),
    .A(_05940_),
    .Y(_05944_),
    .D(_05943_));
 sg13g2_mux2_1 _22406_ (.A0(\top_ihp.oisc.regs[20][22] ),
    .A1(\top_ihp.oisc.regs[16][22] ),
    .S(net654),
    .X(_05945_));
 sg13g2_a22oi_1 _22407_ (.Y(_05946_),
    .B1(_05945_),
    .B2(net640),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][22] ));
 sg13g2_mux2_1 _22408_ (.A0(\top_ihp.oisc.regs[30][22] ),
    .A1(\top_ihp.oisc.regs[26][22] ),
    .S(net678),
    .X(_05947_));
 sg13g2_and2_1 _22409_ (.A(_04930_),
    .B(_05947_),
    .X(_05948_));
 sg13g2_a221oi_1 _22410_ (.B2(\top_ihp.oisc.regs[5][22] ),
    .C1(_05948_),
    .B1(net469),
    .A1(\top_ihp.oisc.regs[29][22] ),
    .Y(_05949_),
    .A2(_05514_));
 sg13g2_o21ai_1 _22411_ (.B1(_05949_),
    .Y(_05950_),
    .A1(net668),
    .A2(_05946_));
 sg13g2_nand2_1 _22412_ (.Y(_05951_),
    .A(\top_ihp.oisc.regs[51][22] ),
    .B(net559));
 sg13g2_a22oi_1 _22413_ (.Y(_05952_),
    .B1(_04827_),
    .B2(\top_ihp.oisc.regs[14][22] ),
    .A2(_03690_),
    .A1(_07444_));
 sg13g2_a22oi_1 _22414_ (.Y(_05953_),
    .B1(net587),
    .B2(\top_ihp.oisc.regs[23][22] ),
    .A2(_04926_),
    .A1(\top_ihp.oisc.regs[15][22] ));
 sg13g2_a22oi_1 _22415_ (.Y(_05954_),
    .B1(net569),
    .B2(\top_ihp.oisc.regs[9][22] ),
    .A2(_05158_),
    .A1(\top_ihp.oisc.regs[21][22] ));
 sg13g2_and4_1 _22416_ (.A(_05951_),
    .B(_05952_),
    .C(_05953_),
    .D(_05954_),
    .X(_05955_));
 sg13g2_a22oi_1 _22417_ (.Y(_05956_),
    .B1(net413),
    .B2(\top_ihp.oisc.regs[57][22] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[2][22] ));
 sg13g2_a22oi_1 _22418_ (.Y(_05957_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][22] ),
    .A2(net269),
    .A1(\top_ihp.oisc.regs[43][22] ));
 sg13g2_nand3_1 _22419_ (.B(_05956_),
    .C(_05957_),
    .A(_05955_),
    .Y(_05958_));
 sg13g2_nor4_1 _22420_ (.A(_04811_),
    .B(_05944_),
    .C(_05950_),
    .D(_05958_),
    .Y(_05959_));
 sg13g2_a21oi_1 _22421_ (.A1(_00129_),
    .A2(net77),
    .Y(_05960_),
    .B1(_05211_));
 sg13g2_a21oi_1 _22422_ (.A1(_07444_),
    .A2(net687),
    .Y(_05961_),
    .B1(_05960_));
 sg13g2_a21oi_1 _22423_ (.A1(_05938_),
    .A2(_05959_),
    .Y(_00308_),
    .B1(_05961_));
 sg13g2_a22oi_1 _22424_ (.Y(_05962_),
    .B1(net594),
    .B2(\top_ihp.oisc.regs[62][23] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[32][23] ));
 sg13g2_a22oi_1 _22425_ (.Y(_05963_),
    .B1(net451),
    .B2(\top_ihp.oisc.regs[40][23] ),
    .A2(net562),
    .A1(\top_ihp.oisc.regs[50][23] ));
 sg13g2_a22oi_1 _22426_ (.Y(_05964_),
    .B1(net273),
    .B2(\top_ihp.oisc.regs[56][23] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][23] ));
 sg13g2_a22oi_1 _22427_ (.Y(_05965_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][23] ),
    .A2(net570),
    .A1(\top_ihp.oisc.regs[57][23] ));
 sg13g2_nand4_1 _22428_ (.B(_05963_),
    .C(_05964_),
    .A(_05962_),
    .Y(_05966_),
    .D(_05965_));
 sg13g2_a22oi_1 _22429_ (.Y(_05967_),
    .B1(net262),
    .B2(\top_ihp.oisc.regs[36][23] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][23] ));
 sg13g2_a22oi_1 _22430_ (.Y(_05968_),
    .B1(net453),
    .B2(\top_ihp.oisc.regs[45][23] ),
    .A2(net604),
    .A1(\top_ihp.oisc.regs[49][23] ));
 sg13g2_a22oi_1 _22431_ (.Y(_05969_),
    .B1(net579),
    .B2(\top_ihp.oisc.regs[48][23] ),
    .A2(net602),
    .A1(\top_ihp.oisc.regs[59][23] ));
 sg13g2_nor2_1 _22432_ (.A(net703),
    .B(_04818_),
    .Y(_05970_));
 sg13g2_buf_2 _22433_ (.A(_05970_),
    .X(_05971_));
 sg13g2_a22oi_1 _22434_ (.Y(_05972_),
    .B1(_05971_),
    .B2(\top_ihp.oisc.regs[16][23] ),
    .A2(net718),
    .A1(\top_ihp.oisc.regs[28][23] ));
 sg13g2_nor2_1 _22435_ (.A(_05130_),
    .B(_05972_),
    .Y(_05973_));
 sg13g2_a21oi_1 _22436_ (.A1(\top_ihp.oisc.regs[44][23] ),
    .A2(net458),
    .Y(_05974_),
    .B1(_05973_));
 sg13g2_nand4_1 _22437_ (.B(_05968_),
    .C(_05969_),
    .A(_05967_),
    .Y(_05975_),
    .D(_05974_));
 sg13g2_a22oi_1 _22438_ (.Y(_05976_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][23] ),
    .A2(net599),
    .A1(\top_ihp.oisc.regs[51][23] ));
 sg13g2_a22oi_1 _22439_ (.Y(_05977_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][23] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][23] ));
 sg13g2_a22oi_1 _22440_ (.Y(_05978_),
    .B1(net447),
    .B2(\top_ihp.oisc.regs[35][23] ),
    .A2(net567),
    .A1(\top_ihp.oisc.regs[61][23] ));
 sg13g2_a22oi_1 _22441_ (.Y(_05979_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[58][23] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][23] ));
 sg13g2_nand4_1 _22442_ (.B(_05977_),
    .C(_05978_),
    .A(_05976_),
    .Y(_05980_),
    .D(_05979_));
 sg13g2_mux2_1 _22443_ (.A0(\top_ihp.oisc.regs[6][23] ),
    .A1(\top_ihp.oisc.regs[2][23] ),
    .S(net678),
    .X(_05981_));
 sg13g2_a22oi_1 _22444_ (.Y(_05982_),
    .B1(_05981_),
    .B2(net644),
    .A2(_05653_),
    .A1(\top_ihp.oisc.regs[14][23] ));
 sg13g2_or2_1 _22445_ (.X(_05983_),
    .B(_05982_),
    .A(_04799_));
 sg13g2_a22oi_1 _22446_ (.Y(_05984_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][23] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[54][23] ));
 sg13g2_nand2_1 _22447_ (.Y(_05985_),
    .A(\top_ihp.oisc.regs[41][23] ),
    .B(net266));
 sg13g2_a22oi_1 _22448_ (.Y(_05986_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[52][23] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[46][23] ));
 sg13g2_nand4_1 _22449_ (.B(_05984_),
    .C(_05985_),
    .A(_05983_),
    .Y(_05987_),
    .D(_05986_));
 sg13g2_nor4_1 _22450_ (.A(_05966_),
    .B(_05975_),
    .C(_05980_),
    .D(_05987_),
    .Y(_05988_));
 sg13g2_a22oi_1 _22451_ (.Y(_05989_),
    .B1(_05519_),
    .B2(\top_ihp.oisc.regs[18][23] ),
    .A2(_04855_),
    .A1(\top_ihp.oisc.regs[20][23] ));
 sg13g2_a22oi_1 _22452_ (.Y(_05990_),
    .B1(_05200_),
    .B2(\top_ihp.oisc.regs[30][23] ),
    .A2(_05237_),
    .A1(\top_ihp.oisc.regs[26][23] ));
 sg13g2_nand2_1 _22453_ (.Y(_05991_),
    .A(_05989_),
    .B(_05990_));
 sg13g2_a221oi_1 _22454_ (.B2(\top_ihp.oisc.regs[12][23] ),
    .C1(_05991_),
    .B1(net421),
    .A1(\top_ihp.oisc.regs[21][23] ),
    .Y(_05992_),
    .A2(net612));
 sg13g2_a22oi_1 _22455_ (.Y(_05993_),
    .B1(_05704_),
    .B2(\top_ihp.oisc.regs[22][23] ),
    .A2(net803),
    .A1(_07442_));
 sg13g2_nand2_1 _22456_ (.Y(_05994_),
    .A(\top_ihp.oisc.regs[23][23] ),
    .B(net648));
 sg13g2_nand2_1 _22457_ (.Y(_05995_),
    .A(_05993_),
    .B(_05994_));
 sg13g2_a221oi_1 _22458_ (.B2(\top_ihp.oisc.regs[15][23] ),
    .C1(_05995_),
    .B1(_04926_),
    .A1(\top_ihp.oisc.regs[7][23] ),
    .Y(_05996_),
    .A2(net617));
 sg13g2_a22oi_1 _22459_ (.Y(_05997_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[43][23] ),
    .A2(net474),
    .A1(\top_ihp.oisc.regs[33][23] ));
 sg13g2_a22oi_1 _22460_ (.Y(_05998_),
    .B1(net596),
    .B2(\top_ihp.oisc.regs[63][23] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][23] ));
 sg13g2_nand4_1 _22461_ (.B(_05996_),
    .C(_05997_),
    .A(_05992_),
    .Y(_05999_),
    .D(_05998_));
 sg13g2_mux2_1 _22462_ (.A0(\top_ihp.oisc.regs[3][23] ),
    .A1(\top_ihp.oisc.regs[19][23] ),
    .S(net676),
    .X(_06000_));
 sg13g2_a22oi_1 _22463_ (.Y(_06001_),
    .B1(net675),
    .B2(_06000_),
    .A2(_05321_),
    .A1(\top_ihp.oisc.regs[10][23] ));
 sg13g2_a22oi_1 _22464_ (.Y(_06002_),
    .B1(net598),
    .B2(\top_ihp.oisc.regs[4][23] ),
    .A2(net469),
    .A1(\top_ihp.oisc.regs[5][23] ));
 sg13g2_a22oi_1 _22465_ (.Y(_06003_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][23] ),
    .A2(_05276_),
    .A1(\top_ihp.oisc.regs[9][23] ));
 sg13g2_a22oi_1 _22466_ (.Y(_06004_),
    .B1(net466),
    .B2(\top_ihp.oisc.regs[1][23] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][23] ));
 sg13g2_nand4_1 _22467_ (.B(_06002_),
    .C(_06003_),
    .A(_06001_),
    .Y(_06005_),
    .D(_06004_));
 sg13g2_a22oi_1 _22468_ (.Y(_06006_),
    .B1(net473),
    .B2(\top_ihp.oisc.regs[13][23] ),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][23] ));
 sg13g2_a22oi_1 _22469_ (.Y(_06007_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][23] ),
    .A2(net555),
    .A1(\top_ihp.oisc.regs[29][23] ));
 sg13g2_nand2_1 _22470_ (.Y(_06008_),
    .A(\top_ihp.oisc.regs[17][23] ),
    .B(net429));
 sg13g2_a22oi_1 _22471_ (.Y(_06009_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][23] ),
    .A2(net465),
    .A1(\top_ihp.oisc.regs[31][23] ));
 sg13g2_nand4_1 _22472_ (.B(_06007_),
    .C(_06008_),
    .A(_06006_),
    .Y(_06010_),
    .D(_06009_));
 sg13g2_nor4_1 _22473_ (.A(net80),
    .B(_05999_),
    .C(_06005_),
    .D(_06010_),
    .Y(_06011_));
 sg13g2_a21oi_1 _22474_ (.A1(_00130_),
    .A2(net77),
    .Y(_06012_),
    .B1(net153));
 sg13g2_a21oi_1 _22475_ (.A1(_07442_),
    .A2(net687),
    .Y(_06013_),
    .B1(_06012_));
 sg13g2_a21oi_1 _22476_ (.A1(_05988_),
    .A2(_06011_),
    .Y(_00309_),
    .B1(_06013_));
 sg13g2_a22oi_1 _22477_ (.Y(_06014_),
    .B1(net268),
    .B2(\top_ihp.oisc.regs[44][24] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][24] ));
 sg13g2_a22oi_1 _22478_ (.Y(_06015_),
    .B1(_05591_),
    .B2(\top_ihp.oisc.regs[37][24] ),
    .A2(net460),
    .A1(\top_ihp.oisc.regs[43][24] ));
 sg13g2_a22oi_1 _22479_ (.Y(_06016_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][24] ),
    .A2(net560),
    .A1(\top_ihp.oisc.regs[48][24] ));
 sg13g2_a22oi_1 _22480_ (.Y(_06017_),
    .B1(net604),
    .B2(\top_ihp.oisc.regs[49][24] ),
    .A2(net476),
    .A1(\top_ihp.oisc.regs[47][24] ));
 sg13g2_nand4_1 _22481_ (.B(_06015_),
    .C(_06016_),
    .A(_06014_),
    .Y(_06018_),
    .D(_06017_));
 sg13g2_a22oi_1 _22482_ (.Y(_06019_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][24] ),
    .A2(net467),
    .A1(\top_ihp.oisc.regs[15][24] ));
 sg13g2_a22oi_1 _22483_ (.Y(_06020_),
    .B1(net470),
    .B2(\top_ihp.oisc.regs[21][24] ),
    .A2(net555),
    .A1(\top_ihp.oisc.regs[29][24] ));
 sg13g2_a22oi_1 _22484_ (.Y(_06021_),
    .B1(_05321_),
    .B2(\top_ihp.oisc.regs[10][24] ),
    .A2(_05547_),
    .A1(\top_ihp.oisc.regs[25][24] ));
 sg13g2_nor2_1 _22485_ (.A(net644),
    .B(net689),
    .Y(_06022_));
 sg13g2_mux2_1 _22486_ (.A0(\top_ihp.oisc.regs[28][24] ),
    .A1(\top_ihp.oisc.regs[24][24] ),
    .S(_04911_),
    .X(_06023_));
 sg13g2_a22oi_1 _22487_ (.Y(_06024_),
    .B1(_06022_),
    .B2(_06023_),
    .A2(net607),
    .A1(\top_ihp.oisc.regs[31][24] ));
 sg13g2_nand4_1 _22488_ (.B(_06020_),
    .C(_06021_),
    .A(_06019_),
    .Y(_06025_),
    .D(_06024_));
 sg13g2_mux2_1 _22489_ (.A0(\top_ihp.oisc.regs[14][24] ),
    .A1(\top_ihp.oisc.regs[12][24] ),
    .S(net656),
    .X(_06026_));
 sg13g2_a22oi_1 _22490_ (.Y(_06027_),
    .B1(_06026_),
    .B2(net650),
    .A2(_05553_),
    .A1(\top_ihp.oisc.regs[8][24] ));
 sg13g2_and2_1 _22491_ (.A(\top_ihp.oisc.regs[7][24] ),
    .B(_05139_),
    .X(_06028_));
 sg13g2_a221oi_1 _22492_ (.B2(\top_ihp.oisc.regs[6][24] ),
    .C1(_06028_),
    .B1(net468),
    .A1(\top_ihp.oisc.regs[5][24] ),
    .Y(_06029_),
    .A2(net469));
 sg13g2_o21ai_1 _22493_ (.B1(_06029_),
    .Y(_06030_),
    .A1(_04896_),
    .A2(_06027_));
 sg13g2_nor4_1 _22494_ (.A(_05538_),
    .B(_06018_),
    .C(_06025_),
    .D(_06030_),
    .Y(_06031_));
 sg13g2_a22oi_1 _22495_ (.Y(_06032_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[38][24] ),
    .A2(_04871_),
    .A1(\top_ihp.oisc.regs[55][24] ));
 sg13g2_a22oi_1 _22496_ (.Y(_06033_),
    .B1(net454),
    .B2(\top_ihp.oisc.regs[34][24] ),
    .A2(net462),
    .A1(\top_ihp.oisc.regs[36][24] ));
 sg13g2_nand2_1 _22497_ (.Y(_06034_),
    .A(\top_ihp.oisc.regs[2][24] ),
    .B(_05180_));
 sg13g2_a22oi_1 _22498_ (.Y(_06035_),
    .B1(_05166_),
    .B2(\top_ihp.oisc.regs[62][24] ),
    .A2(net474),
    .A1(\top_ihp.oisc.regs[33][24] ));
 sg13g2_nand4_1 _22499_ (.B(_06033_),
    .C(_06034_),
    .A(_06032_),
    .Y(_06036_),
    .D(_06035_));
 sg13g2_a22oi_1 _22500_ (.Y(_06037_),
    .B1(_05300_),
    .B2(\top_ihp.oisc.regs[41][24] ),
    .A2(net591),
    .A1(\top_ihp.oisc.regs[52][24] ));
 sg13g2_a22oi_1 _22501_ (.Y(_06038_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][24] ),
    .A2(net559),
    .A1(\top_ihp.oisc.regs[51][24] ));
 sg13g2_a22oi_1 _22502_ (.Y(_06039_),
    .B1(net562),
    .B2(\top_ihp.oisc.regs[50][24] ),
    .A2(_04975_),
    .A1(\top_ihp.oisc.regs[42][24] ));
 sg13g2_a22oi_1 _22503_ (.Y(_06040_),
    .B1(_05971_),
    .B2(\top_ihp.oisc.regs[18][24] ),
    .A2(net718),
    .A1(\top_ihp.oisc.regs[30][24] ));
 sg13g2_inv_1 _22504_ (.Y(_06041_),
    .A(_06040_));
 sg13g2_a22oi_1 _22505_ (.Y(_06042_),
    .B1(net671),
    .B2(_06041_),
    .A2(net596),
    .A1(\top_ihp.oisc.regs[63][24] ));
 sg13g2_nand4_1 _22506_ (.B(_06038_),
    .C(_06039_),
    .A(_06037_),
    .Y(_06043_),
    .D(_06042_));
 sg13g2_nand2_1 _22507_ (.Y(_06044_),
    .A(\top_ihp.oisc.regs[27][24] ),
    .B(net584));
 sg13g2_a22oi_1 _22508_ (.Y(_06045_),
    .B1(net574),
    .B2(\top_ihp.oisc.regs[26][24] ),
    .A2(net772),
    .A1(_07626_));
 sg13g2_a22oi_1 _22509_ (.Y(_06046_),
    .B1(_05241_),
    .B2(\top_ihp.oisc.regs[19][24] ),
    .A2(net645),
    .A1(\top_ihp.oisc.regs[16][24] ));
 sg13g2_a22oi_1 _22510_ (.Y(_06047_),
    .B1(net721),
    .B2(\top_ihp.oisc.regs[22][24] ),
    .A2(net722),
    .A1(\top_ihp.oisc.regs[20][24] ));
 sg13g2_nor2_1 _22511_ (.A(net672),
    .B(_06047_),
    .Y(_06048_));
 sg13g2_a21oi_1 _22512_ (.A1(\top_ihp.oisc.regs[3][24] ),
    .A2(_05245_),
    .Y(_06049_),
    .B1(_06048_));
 sg13g2_and4_1 _22513_ (.A(_06044_),
    .B(_06045_),
    .C(_06046_),
    .D(_06049_),
    .X(_06050_));
 sg13g2_a22oi_1 _22514_ (.Y(_06051_),
    .B1(net577),
    .B2(\top_ihp.oisc.regs[4][24] ),
    .A2(net597),
    .A1(\top_ihp.oisc.regs[9][24] ));
 sg13g2_a22oi_1 _22515_ (.Y(_06052_),
    .B1(_04936_),
    .B2(\top_ihp.oisc.regs[1][24] ),
    .A2(_04821_),
    .A1(\top_ihp.oisc.regs[17][24] ));
 sg13g2_and2_1 _22516_ (.A(_06051_),
    .B(_06052_),
    .X(_06053_));
 sg13g2_a22oi_1 _22517_ (.Y(_06054_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][24] ),
    .A2(net432),
    .A1(\top_ihp.oisc.regs[32][24] ));
 sg13g2_a22oi_1 _22518_ (.Y(_06055_),
    .B1(net273),
    .B2(\top_ihp.oisc.regs[56][24] ),
    .A2(net602),
    .A1(\top_ihp.oisc.regs[59][24] ));
 sg13g2_nand4_1 _22519_ (.B(_06053_),
    .C(_06054_),
    .A(_06050_),
    .Y(_06056_),
    .D(_06055_));
 sg13g2_a22oi_1 _22520_ (.Y(_06057_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][24] ),
    .A2(_05215_),
    .A1(\top_ihp.oisc.regs[54][24] ));
 sg13g2_a22oi_1 _22521_ (.Y(_06058_),
    .B1(_05219_),
    .B2(\top_ihp.oisc.regs[40][24] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[39][24] ));
 sg13g2_a22oi_1 _22522_ (.Y(_06059_),
    .B1(_05310_),
    .B2(\top_ihp.oisc.regs[46][24] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][24] ));
 sg13g2_a22oi_1 _22523_ (.Y(_06060_),
    .B1(_04765_),
    .B2(\top_ihp.oisc.regs[13][24] ),
    .A2(_04763_),
    .A1(\top_ihp.oisc.regs[11][24] ));
 sg13g2_nor3_1 _22524_ (.A(net644),
    .B(_05017_),
    .C(_06060_),
    .Y(_06061_));
 sg13g2_a21oi_1 _22525_ (.A1(\top_ihp.oisc.regs[35][24] ),
    .A2(net457),
    .Y(_06062_),
    .B1(_06061_));
 sg13g2_nand4_1 _22526_ (.B(_06058_),
    .C(_06059_),
    .A(_06057_),
    .Y(_06063_),
    .D(_06062_));
 sg13g2_nor4_2 _22527_ (.A(_06036_),
    .B(_06043_),
    .C(_06056_),
    .Y(_06064_),
    .D(_06063_));
 sg13g2_buf_1 _22528_ (.A(_05104_),
    .X(_06065_));
 sg13g2_a21oi_1 _22529_ (.A1(_00131_),
    .A2(_05354_),
    .Y(_06066_),
    .B1(_06065_));
 sg13g2_a21oi_1 _22530_ (.A1(_07626_),
    .A2(_05418_),
    .Y(_06067_),
    .B1(_06066_));
 sg13g2_a21oi_1 _22531_ (.A1(_06031_),
    .A2(_06064_),
    .Y(_00310_),
    .B1(_06067_));
 sg13g2_a22oi_1 _22532_ (.Y(_06068_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][25] ),
    .A2(_04899_),
    .A1(\top_ihp.oisc.regs[10][25] ));
 sg13g2_a22oi_1 _22533_ (.Y(_06069_),
    .B1(net419),
    .B2(\top_ihp.oisc.regs[5][25] ),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][25] ));
 sg13g2_a22oi_1 _22534_ (.Y(_06070_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][25] ),
    .A2(net618),
    .A1(\top_ihp.oisc.regs[17][25] ));
 sg13g2_a22oi_1 _22535_ (.Y(_06071_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][25] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][25] ));
 sg13g2_nand4_1 _22536_ (.B(_06069_),
    .C(_06070_),
    .A(_06068_),
    .Y(_06072_),
    .D(_06071_));
 sg13g2_mux2_1 _22537_ (.A0(\top_ihp.oisc.regs[20][25] ),
    .A1(\top_ihp.oisc.regs[16][25] ),
    .S(_04931_),
    .X(_06073_));
 sg13g2_a22oi_1 _22538_ (.Y(_06074_),
    .B1(_06073_),
    .B2(net640),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][25] ));
 sg13g2_nor2_2 _22539_ (.A(net668),
    .B(_06074_),
    .Y(_06075_));
 sg13g2_a22oi_1 _22540_ (.Y(_06076_),
    .B1(net468),
    .B2(\top_ihp.oisc.regs[6][25] ),
    .A2(net472),
    .A1(\top_ihp.oisc.regs[29][25] ));
 sg13g2_a22oi_1 _22541_ (.Y(_06077_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][25] ),
    .A2(net470),
    .A1(\top_ihp.oisc.regs[21][25] ));
 sg13g2_nand2_1 _22542_ (.Y(_06078_),
    .A(_06076_),
    .B(_06077_));
 sg13g2_a22oi_1 _22543_ (.Y(_06079_),
    .B1(_05035_),
    .B2(\top_ihp.oisc.regs[56][25] ),
    .A2(_04969_),
    .A1(\top_ihp.oisc.regs[54][25] ));
 sg13g2_a22oi_1 _22544_ (.Y(_06080_),
    .B1(_05093_),
    .B2(\top_ihp.oisc.regs[41][25] ),
    .A2(_04869_),
    .A1(\top_ihp.oisc.regs[55][25] ));
 sg13g2_a22oi_1 _22545_ (.Y(_06081_),
    .B1(_05051_),
    .B2(\top_ihp.oisc.regs[61][25] ),
    .A2(_04983_),
    .A1(\top_ihp.oisc.regs[58][25] ));
 sg13g2_a22oi_1 _22546_ (.Y(_06082_),
    .B1(_05085_),
    .B2(\top_ihp.oisc.regs[40][25] ),
    .A2(_05030_),
    .A1(\top_ihp.oisc.regs[63][25] ));
 sg13g2_nand4_1 _22547_ (.B(_06080_),
    .C(_06081_),
    .A(_06079_),
    .Y(_06083_),
    .D(_06082_));
 sg13g2_a22oi_1 _22548_ (.Y(_06084_),
    .B1(net573),
    .B2(\top_ihp.oisc.regs[31][25] ),
    .A2(net655),
    .A1(\top_ihp.oisc.regs[13][25] ));
 sg13g2_mux2_1 _22549_ (.A0(\top_ihp.oisc.regs[3][25] ),
    .A1(\top_ihp.oisc.regs[19][25] ),
    .S(net725),
    .X(_06085_));
 sg13g2_nor2_1 _22550_ (.A(_07811_),
    .B(_03679_),
    .Y(_06086_));
 sg13g2_a221oi_1 _22551_ (.B2(_04957_),
    .C1(_06086_),
    .B1(_06085_),
    .A1(\top_ihp.oisc.regs[22][25] ),
    .Y(_06087_),
    .A2(_05704_));
 sg13g2_a22oi_1 _22552_ (.Y(_06088_),
    .B1(net648),
    .B2(\top_ihp.oisc.regs[23][25] ),
    .A2(net565),
    .A1(\top_ihp.oisc.regs[1][25] ));
 sg13g2_a22oi_1 _22553_ (.Y(_06089_),
    .B1(_05015_),
    .B2(\top_ihp.oisc.regs[4][25] ),
    .A2(net657),
    .A1(\top_ihp.oisc.regs[7][25] ));
 sg13g2_nand4_1 _22554_ (.B(_06087_),
    .C(_06088_),
    .A(_06084_),
    .Y(_06090_),
    .D(_06089_));
 sg13g2_a22oi_1 _22555_ (.Y(_06091_),
    .B1(net563),
    .B2(\top_ihp.oisc.regs[49][25] ),
    .A2(_04843_),
    .A1(\top_ihp.oisc.regs[47][25] ));
 sg13g2_nand2_1 _22556_ (.Y(_06092_),
    .A(\top_ihp.oisc.regs[45][25] ),
    .B(_05076_));
 sg13g2_nand2_1 _22557_ (.Y(_06093_),
    .A(\top_ihp.oisc.regs[26][25] ),
    .B(net574));
 sg13g2_a22oi_1 _22558_ (.Y(_06094_),
    .B1(net554),
    .B2(\top_ihp.oisc.regs[18][25] ),
    .A2(_05200_),
    .A1(\top_ihp.oisc.regs[30][25] ));
 sg13g2_nand4_1 _22559_ (.B(_06092_),
    .C(_06093_),
    .A(_06091_),
    .Y(_06095_),
    .D(_06094_));
 sg13g2_or4_1 _22560_ (.A(_04809_),
    .B(_06083_),
    .C(_06090_),
    .D(_06095_),
    .X(_06096_));
 sg13g2_nor4_1 _22561_ (.A(_06072_),
    .B(_06075_),
    .C(_06078_),
    .D(_06096_),
    .Y(_06097_));
 sg13g2_a22oi_1 _22562_ (.Y(_06098_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[52][25] ),
    .A2(_05320_),
    .A1(\top_ihp.oisc.regs[14][25] ));
 sg13g2_and2_1 _22563_ (.A(\top_ihp.oisc.regs[2][25] ),
    .B(net600),
    .X(_06099_));
 sg13g2_a221oi_1 _22564_ (.B2(\top_ihp.oisc.regs[57][25] ),
    .C1(_06099_),
    .B1(net570),
    .A1(\top_ihp.oisc.regs[48][25] ),
    .Y(_06100_),
    .A2(net560));
 sg13g2_a22oi_1 _22565_ (.Y(_06101_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[59][25] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][25] ));
 sg13g2_a22oi_1 _22566_ (.Y(_06102_),
    .B1(net270),
    .B2(\top_ihp.oisc.regs[46][25] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[38][25] ));
 sg13g2_nand4_1 _22567_ (.B(_06100_),
    .C(_06101_),
    .A(_06098_),
    .Y(_06103_),
    .D(_06102_));
 sg13g2_a22oi_1 _22568_ (.Y(_06104_),
    .B1(_05073_),
    .B2(\top_ihp.oisc.regs[34][25] ),
    .A2(net553),
    .A1(\top_ihp.oisc.regs[62][25] ));
 sg13g2_a22oi_1 _22569_ (.Y(_06105_),
    .B1(net595),
    .B2(\top_ihp.oisc.regs[50][25] ),
    .A2(net581),
    .A1(\top_ihp.oisc.regs[51][25] ));
 sg13g2_a22oi_1 _22570_ (.Y(_06106_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[35][25] ),
    .A2(net434),
    .A1(\top_ihp.oisc.regs[32][25] ));
 sg13g2_a22oi_1 _22571_ (.Y(_06107_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][25] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][25] ));
 sg13g2_nand4_1 _22572_ (.B(_06105_),
    .C(_06106_),
    .A(_06104_),
    .Y(_06108_),
    .D(_06107_));
 sg13g2_a22oi_1 _22573_ (.Y(_06109_),
    .B1(_05114_),
    .B2(\top_ihp.oisc.regs[44][25] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][25] ));
 sg13g2_a22oi_1 _22574_ (.Y(_06110_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][25] ),
    .A2(net262),
    .A1(\top_ihp.oisc.regs[36][25] ));
 sg13g2_nor2_1 _22575_ (.A(net666),
    .B(net681),
    .Y(_06111_));
 sg13g2_a22oi_1 _22576_ (.Y(_06112_),
    .B1(_05553_),
    .B2(\top_ihp.oisc.regs[9][25] ),
    .A2(_06111_),
    .A1(\top_ihp.oisc.regs[15][25] ));
 sg13g2_nor3_1 _22577_ (.A(net640),
    .B(net691),
    .C(_06112_),
    .Y(_06113_));
 sg13g2_a221oi_1 _22578_ (.B2(\top_ihp.oisc.regs[39][25] ),
    .C1(_06113_),
    .B1(net452),
    .A1(\top_ihp.oisc.regs[43][25] ),
    .Y(_06114_),
    .A2(_05367_));
 sg13g2_nand3_1 _22579_ (.B(_06110_),
    .C(_06114_),
    .A(_06109_),
    .Y(_06115_));
 sg13g2_nor3_2 _22580_ (.A(_06103_),
    .B(_06108_),
    .C(_06115_),
    .Y(_06116_));
 sg13g2_a21oi_1 _22581_ (.A1(_00132_),
    .A2(net78),
    .Y(_06117_),
    .B1(net154));
 sg13g2_nor2_1 _22582_ (.A(_06086_),
    .B(_06117_),
    .Y(_06118_));
 sg13g2_a21oi_1 _22583_ (.A1(_06097_),
    .A2(_06116_),
    .Y(_00311_),
    .B1(_06118_));
 sg13g2_a22oi_1 _22584_ (.Y(_06119_),
    .B1(net581),
    .B2(\top_ihp.oisc.regs[51][26] ),
    .A2(net442),
    .A1(\top_ihp.oisc.regs[58][26] ));
 sg13g2_a22oi_1 _22585_ (.Y(_06120_),
    .B1(net264),
    .B2(\top_ihp.oisc.regs[45][26] ),
    .A2(net578),
    .A1(\top_ihp.oisc.regs[50][26] ));
 sg13g2_a22oi_1 _22586_ (.Y(_06121_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][26] ),
    .A2(_05109_),
    .A1(\top_ihp.oisc.regs[55][26] ));
 sg13g2_a22oi_1 _22587_ (.Y(_06122_),
    .B1(_05107_),
    .B2(\top_ihp.oisc.regs[46][26] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[35][26] ));
 sg13g2_nand4_1 _22588_ (.B(_06120_),
    .C(_06121_),
    .A(_06119_),
    .Y(_06123_),
    .D(_06122_));
 sg13g2_a22oi_1 _22589_ (.Y(_06124_),
    .B1(net601),
    .B2(\top_ihp.oisc.regs[48][26] ),
    .A2(net267),
    .A1(\top_ihp.oisc.regs[38][26] ));
 sg13g2_a22oi_1 _22590_ (.Y(_06125_),
    .B1(net553),
    .B2(\top_ihp.oisc.regs[62][26] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][26] ));
 sg13g2_a22oi_1 _22591_ (.Y(_06126_),
    .B1(_05073_),
    .B2(\top_ihp.oisc.regs[34][26] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[57][26] ));
 sg13g2_a22oi_1 _22592_ (.Y(_06127_),
    .B1(_05224_),
    .B2(\top_ihp.oisc.regs[36][26] ),
    .A2(_05226_),
    .A1(\top_ihp.oisc.regs[32][26] ));
 sg13g2_nand4_1 _22593_ (.B(_06125_),
    .C(_06126_),
    .A(_06124_),
    .Y(_06128_),
    .D(_06127_));
 sg13g2_a22oi_1 _22594_ (.Y(_06129_),
    .B1(net611),
    .B2(\top_ihp.oisc.regs[5][26] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][26] ));
 sg13g2_a22oi_1 _22595_ (.Y(_06130_),
    .B1(_05196_),
    .B2(\top_ihp.oisc.regs[4][26] ),
    .A2(net477),
    .A1(\top_ihp.oisc.regs[14][26] ));
 sg13g2_mux2_1 _22596_ (.A0(\top_ihp.oisc.regs[3][26] ),
    .A1(\top_ihp.oisc.regs[19][26] ),
    .S(net693),
    .X(_06131_));
 sg13g2_a22oi_1 _22597_ (.Y(_06132_),
    .B1(_06131_),
    .B2(_04958_),
    .A2(net585),
    .A1(\top_ihp.oisc.regs[12][26] ));
 sg13g2_a22oi_1 _22598_ (.Y(_06133_),
    .B1(net651),
    .B2(\top_ihp.oisc.regs[11][26] ),
    .A2(net607),
    .A1(\top_ihp.oisc.regs[31][26] ));
 sg13g2_and4_1 _22599_ (.A(_06129_),
    .B(_06130_),
    .C(_06132_),
    .D(_06133_),
    .X(_06134_));
 sg13g2_nand2_1 _22600_ (.Y(_06135_),
    .A(\top_ihp.oisc.regs[30][26] ),
    .B(net576));
 sg13g2_a22oi_1 _22601_ (.Y(_06136_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[22][26] ),
    .A2(_04855_),
    .A1(\top_ihp.oisc.regs[20][26] ));
 sg13g2_nand2_1 _22602_ (.Y(_06137_),
    .A(\top_ihp.oisc.regs[9][26] ),
    .B(_05022_));
 sg13g2_a22oi_1 _22603_ (.Y(_06138_),
    .B1(net574),
    .B2(\top_ihp.oisc.regs[26][26] ),
    .A2(net764),
    .A1(net1030));
 sg13g2_nand4_1 _22604_ (.B(_06136_),
    .C(_06137_),
    .A(_06135_),
    .Y(_06139_),
    .D(_06138_));
 sg13g2_a221oi_1 _22605_ (.B2(\top_ihp.oisc.regs[40][26] ),
    .C1(_06139_),
    .B1(net259),
    .A1(\top_ihp.oisc.regs[63][26] ),
    .Y(_06140_),
    .A2(net571));
 sg13g2_a22oi_1 _22606_ (.Y(_06141_),
    .B1(_04901_),
    .B2(\top_ihp.oisc.regs[21][26] ),
    .A2(_04892_),
    .A1(\top_ihp.oisc.regs[29][26] ));
 sg13g2_a22oi_1 _22607_ (.Y(_06142_),
    .B1(_05153_),
    .B2(\top_ihp.oisc.regs[27][26] ),
    .A2(net655),
    .A1(\top_ihp.oisc.regs[13][26] ));
 sg13g2_mux2_1 _22608_ (.A0(\top_ihp.oisc.regs[6][26] ),
    .A1(\top_ihp.oisc.regs[2][26] ),
    .S(net704),
    .X(_06143_));
 sg13g2_a22oi_1 _22609_ (.Y(_06144_),
    .B1(_05727_),
    .B2(_06143_),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][26] ));
 sg13g2_a22oi_1 _22610_ (.Y(_06145_),
    .B1(_04935_),
    .B2(\top_ihp.oisc.regs[1][26] ),
    .A2(net653),
    .A1(\top_ihp.oisc.regs[15][26] ));
 sg13g2_nand4_1 _22611_ (.B(_06142_),
    .C(_06144_),
    .A(_06141_),
    .Y(_06146_),
    .D(_06145_));
 sg13g2_a221oi_1 _22612_ (.B2(\top_ihp.oisc.regs[52][26] ),
    .C1(_06146_),
    .B1(net455),
    .A1(\top_ihp.oisc.regs[54][26] ),
    .Y(_06147_),
    .A2(net606));
 sg13g2_nand3_1 _22613_ (.B(_06140_),
    .C(_06147_),
    .A(_06134_),
    .Y(_06148_));
 sg13g2_nor3_1 _22614_ (.A(_06123_),
    .B(_06128_),
    .C(_06148_),
    .Y(_06149_));
 sg13g2_mux2_1 _22615_ (.A0(\top_ihp.oisc.regs[24][26] ),
    .A1(\top_ihp.oisc.regs[16][26] ),
    .S(_05282_),
    .X(_06150_));
 sg13g2_a22oi_1 _22616_ (.Y(_06151_),
    .B1(_06150_),
    .B2(net556),
    .A2(_05653_),
    .A1(\top_ihp.oisc.regs[28][26] ));
 sg13g2_nor2_1 _22617_ (.A(net668),
    .B(_06151_),
    .Y(_06152_));
 sg13g2_a22oi_1 _22618_ (.Y(_06153_),
    .B1(_05083_),
    .B2(\top_ihp.oisc.regs[25][26] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[23][26] ));
 sg13g2_and3_1 _22619_ (.X(_06154_),
    .A(\top_ihp.oisc.regs[18][26] ),
    .B(net644),
    .C(net671));
 sg13g2_nand2_1 _22620_ (.Y(_06155_),
    .A(\top_ihp.oisc.regs[10][26] ),
    .B(net677));
 sg13g2_nand2_1 _22621_ (.Y(_06156_),
    .A(\top_ihp.oisc.regs[8][26] ),
    .B(net656));
 sg13g2_a21oi_1 _22622_ (.A1(_06155_),
    .A2(_06156_),
    .Y(_06157_),
    .B1(net679));
 sg13g2_o21ai_1 _22623_ (.B1(net556),
    .Y(_06158_),
    .A1(_06154_),
    .A2(_06157_));
 sg13g2_o21ai_1 _22624_ (.B1(_06158_),
    .Y(_06159_),
    .A1(_04878_),
    .A2(_06153_));
 sg13g2_a22oi_1 _22625_ (.Y(_06160_),
    .B1(net602),
    .B2(\top_ihp.oisc.regs[59][26] ),
    .A2(net476),
    .A1(\top_ihp.oisc.regs[47][26] ));
 sg13g2_a22oi_1 _22626_ (.Y(_06161_),
    .B1(_05079_),
    .B2(\top_ihp.oisc.regs[39][26] ),
    .A2(net458),
    .A1(\top_ihp.oisc.regs[44][26] ));
 sg13g2_a22oi_1 _22627_ (.Y(_06162_),
    .B1(_05096_),
    .B2(\top_ihp.oisc.regs[60][26] ),
    .A2(_04974_),
    .A1(\top_ihp.oisc.regs[42][26] ));
 sg13g2_a22oi_1 _22628_ (.Y(_06163_),
    .B1(net460),
    .B2(\top_ihp.oisc.regs[43][26] ),
    .A2(_04978_),
    .A1(\top_ihp.oisc.regs[49][26] ));
 sg13g2_and4_1 _22629_ (.A(_06160_),
    .B(_06161_),
    .C(_06162_),
    .D(_06163_),
    .X(_06164_));
 sg13g2_a22oi_1 _22630_ (.Y(_06165_),
    .B1(net255),
    .B2(\top_ihp.oisc.regs[56][26] ),
    .A2(_05217_),
    .A1(\top_ihp.oisc.regs[33][26] ));
 sg13g2_a22oi_1 _22631_ (.Y(_06166_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][26] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[61][26] ));
 sg13g2_nand3_1 _22632_ (.B(_06165_),
    .C(_06166_),
    .A(_06164_),
    .Y(_06167_));
 sg13g2_nor4_1 _22633_ (.A(_05210_),
    .B(_06152_),
    .C(_06159_),
    .D(_06167_),
    .Y(_06168_));
 sg13g2_buf_8 _22634_ (.A(_04810_),
    .X(_06169_));
 sg13g2_a21oi_1 _22635_ (.A1(_00133_),
    .A2(net75),
    .Y(_06170_),
    .B1(net152));
 sg13g2_a21oi_1 _22636_ (.A1(_07614_),
    .A2(_05418_),
    .Y(_06171_),
    .B1(_06170_));
 sg13g2_a21oi_1 _22637_ (.A1(_06149_),
    .A2(_06168_),
    .Y(_00312_),
    .B1(_06171_));
 sg13g2_a22oi_1 _22638_ (.Y(_06172_),
    .B1(net610),
    .B2(\top_ihp.oisc.regs[6][27] ),
    .A2(_04816_),
    .A1(\top_ihp.oisc.regs[25][27] ));
 sg13g2_a22oi_1 _22639_ (.Y(_06173_),
    .B1(net646),
    .B2(\top_ihp.oisc.regs[30][27] ),
    .A2(net764),
    .A1(_07681_));
 sg13g2_nand2_1 _22640_ (.Y(_06174_),
    .A(\top_ihp.oisc.regs[11][27] ),
    .B(net647));
 sg13g2_nand3_1 _22641_ (.B(_06173_),
    .C(_06174_),
    .A(_06172_),
    .Y(_06175_));
 sg13g2_a221oi_1 _22642_ (.B2(\top_ihp.oisc.regs[45][27] ),
    .C1(_06175_),
    .B1(net438),
    .A1(\top_ihp.oisc.regs[33][27] ),
    .Y(_06176_),
    .A2(net474));
 sg13g2_a22oi_1 _22643_ (.Y(_06177_),
    .B1(net557),
    .B2(\top_ihp.oisc.regs[4][27] ),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[8][27] ));
 sg13g2_nor3_1 _22644_ (.A(net677),
    .B(_05119_),
    .C(_06177_),
    .Y(_06178_));
 sg13g2_a22oi_1 _22645_ (.Y(_06179_),
    .B1(net557),
    .B2(\top_ihp.oisc.regs[23][27] ),
    .A2(net588),
    .A1(\top_ihp.oisc.regs[27][27] ));
 sg13g2_nor3_1 _22646_ (.A(_04877_),
    .B(_04878_),
    .C(_06179_),
    .Y(_06180_));
 sg13g2_nor2_1 _22647_ (.A(_06178_),
    .B(_06180_),
    .Y(_06181_));
 sg13g2_a22oi_1 _22648_ (.Y(_06182_),
    .B1(_05080_),
    .B2(\top_ihp.oisc.regs[39][27] ),
    .A2(net568),
    .A1(\top_ihp.oisc.regs[59][27] ));
 sg13g2_nand3_1 _22649_ (.B(_06181_),
    .C(_06182_),
    .A(_06176_),
    .Y(_06183_));
 sg13g2_nor3_2 _22650_ (.A(net666),
    .B(net681),
    .C(net691),
    .Y(_06184_));
 sg13g2_mux2_1 _22651_ (.A0(\top_ihp.oisc.regs[15][27] ),
    .A1(\top_ihp.oisc.regs[7][27] ),
    .S(net644),
    .X(_06185_));
 sg13g2_a22oi_1 _22652_ (.Y(_06186_),
    .B1(_06184_),
    .B2(_06185_),
    .A2(net470),
    .A1(\top_ihp.oisc.regs[21][27] ));
 sg13g2_nand3_1 _22653_ (.B(net643),
    .C(net797),
    .A(\top_ihp.oisc.regs[24][27] ),
    .Y(_06187_));
 sg13g2_nand3_1 _22654_ (.B(_05281_),
    .C(net690),
    .A(\top_ihp.oisc.regs[18][27] ),
    .Y(_06188_));
 sg13g2_nand2_1 _22655_ (.Y(_06189_),
    .A(_06187_),
    .B(_06188_));
 sg13g2_mux2_1 _22656_ (.A0(\top_ihp.oisc.regs[3][27] ),
    .A1(\top_ihp.oisc.regs[19][27] ),
    .S(net693),
    .X(_06190_));
 sg13g2_a22oi_1 _22657_ (.Y(_06191_),
    .B1(_06190_),
    .B2(net675),
    .A2(_06189_),
    .A1(net556));
 sg13g2_a22oi_1 _22658_ (.Y(_06192_),
    .B1(_04941_),
    .B2(\top_ihp.oisc.regs[31][27] ),
    .A2(_04909_),
    .A1(\top_ihp.oisc.regs[5][27] ));
 sg13g2_a22oi_1 _22659_ (.Y(_06193_),
    .B1(net466),
    .B2(\top_ihp.oisc.regs[1][27] ),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][27] ));
 sg13g2_nand4_1 _22660_ (.B(_06191_),
    .C(_06192_),
    .A(_06186_),
    .Y(_06194_),
    .D(_06193_));
 sg13g2_mux2_1 _22661_ (.A0(\top_ihp.oisc.regs[20][27] ),
    .A1(\top_ihp.oisc.regs[16][27] ),
    .S(_04911_),
    .X(_06195_));
 sg13g2_a22oi_1 _22662_ (.Y(_06196_),
    .B1(_06195_),
    .B2(net640),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][27] ));
 sg13g2_and2_1 _22663_ (.A(\top_ihp.oisc.regs[17][27] ),
    .B(net618),
    .X(_06197_));
 sg13g2_a221oi_1 _22664_ (.B2(\top_ihp.oisc.regs[9][27] ),
    .C1(_06197_),
    .B1(net422),
    .A1(\top_ihp.oisc.regs[29][27] ),
    .Y(_06198_),
    .A2(net555));
 sg13g2_o21ai_1 _22665_ (.B1(_06198_),
    .Y(_06199_),
    .A1(net668),
    .A2(_06196_));
 sg13g2_nor4_1 _22666_ (.A(net76),
    .B(_06183_),
    .C(_06194_),
    .D(_06199_),
    .Y(_06200_));
 sg13g2_a22oi_1 _22667_ (.Y(_06201_),
    .B1(net255),
    .B2(\top_ihp.oisc.regs[56][27] ),
    .A2(_04989_),
    .A1(\top_ihp.oisc.regs[36][27] ));
 sg13g2_a22oi_1 _22668_ (.Y(_06202_),
    .B1(_05059_),
    .B2(\top_ihp.oisc.regs[46][27] ),
    .A2(_04871_),
    .A1(\top_ihp.oisc.regs[55][27] ));
 sg13g2_a22oi_1 _22669_ (.Y(_06203_),
    .B1(net450),
    .B2(\top_ihp.oisc.regs[37][27] ),
    .A2(_04975_),
    .A1(\top_ihp.oisc.regs[42][27] ));
 sg13g2_a22oi_1 _22670_ (.Y(_06204_),
    .B1(_05367_),
    .B2(\top_ihp.oisc.regs[43][27] ),
    .A2(_05359_),
    .A1(\top_ihp.oisc.regs[49][27] ));
 sg13g2_nand4_1 _22671_ (.B(_06202_),
    .C(_06203_),
    .A(_06201_),
    .Y(_06205_),
    .D(_06204_));
 sg13g2_a22oi_1 _22672_ (.Y(_06206_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][27] ),
    .A2(net570),
    .A1(\top_ihp.oisc.regs[57][27] ));
 sg13g2_nand2_1 _22673_ (.Y(_06207_),
    .A(\top_ihp.oisc.regs[60][27] ),
    .B(net590));
 sg13g2_a22oi_1 _22674_ (.Y(_06208_),
    .B1(_05971_),
    .B2(\top_ihp.oisc.regs[2][27] ),
    .A2(net718),
    .A1(\top_ihp.oisc.regs[14][27] ));
 sg13g2_nor2_1 _22675_ (.A(_04799_),
    .B(_06208_),
    .Y(_06209_));
 sg13g2_a21oi_1 _22676_ (.A1(\top_ihp.oisc.regs[38][27] ),
    .A2(net461),
    .Y(_06210_),
    .B1(_06209_));
 sg13g2_a22oi_1 _22677_ (.Y(_06211_),
    .B1(net566),
    .B2(\top_ihp.oisc.regs[58][27] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][27] ));
 sg13g2_nand4_1 _22678_ (.B(_06207_),
    .C(_06210_),
    .A(_06206_),
    .Y(_06212_),
    .D(_06211_));
 sg13g2_a22oi_1 _22679_ (.Y(_06213_),
    .B1(_05171_),
    .B2(\top_ihp.oisc.regs[52][27] ),
    .A2(net599),
    .A1(\top_ihp.oisc.regs[51][27] ));
 sg13g2_a22oi_1 _22680_ (.Y(_06214_),
    .B1(net571),
    .B2(\top_ihp.oisc.regs[63][27] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][27] ));
 sg13g2_a22oi_1 _22681_ (.Y(_06215_),
    .B1(net261),
    .B2(\top_ihp.oisc.regs[44][27] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][27] ));
 sg13g2_a22oi_1 _22682_ (.Y(_06216_),
    .B1(net557),
    .B2(\top_ihp.oisc.regs[22][27] ),
    .A2(_05131_),
    .A1(\top_ihp.oisc.regs[26][27] ));
 sg13g2_nor2b_1 _22683_ (.A(_06216_),
    .B_N(net671),
    .Y(_06217_));
 sg13g2_a21oi_1 _22684_ (.A1(\top_ihp.oisc.regs[50][27] ),
    .A2(_05361_),
    .Y(_06218_),
    .B1(_06217_));
 sg13g2_nand4_1 _22685_ (.B(_06214_),
    .C(_06215_),
    .A(_06213_),
    .Y(_06219_),
    .D(_06218_));
 sg13g2_a22oi_1 _22686_ (.Y(_06220_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[35][27] ),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[48][27] ));
 sg13g2_a22oi_1 _22687_ (.Y(_06221_),
    .B1(_05300_),
    .B2(\top_ihp.oisc.regs[41][27] ),
    .A2(_05383_),
    .A1(\top_ihp.oisc.regs[61][27] ));
 sg13g2_a22oi_1 _22688_ (.Y(_06222_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][27] ),
    .A2(net594),
    .A1(\top_ihp.oisc.regs[62][27] ));
 sg13g2_a22oi_1 _22689_ (.Y(_06223_),
    .B1(_04765_),
    .B2(\top_ihp.oisc.regs[12][27] ),
    .A2(_04763_),
    .A1(\top_ihp.oisc.regs[10][27] ));
 sg13g2_nor2_1 _22690_ (.A(net679),
    .B(_06223_),
    .Y(_06224_));
 sg13g2_a21oi_1 _22691_ (.A1(\top_ihp.oisc.regs[32][27] ),
    .A2(net432),
    .Y(_06225_),
    .B1(_06224_));
 sg13g2_nand4_1 _22692_ (.B(_06221_),
    .C(_06222_),
    .A(_06220_),
    .Y(_06226_),
    .D(_06225_));
 sg13g2_nor4_2 _22693_ (.A(_06205_),
    .B(_06212_),
    .C(_06219_),
    .Y(_06227_),
    .D(_06226_));
 sg13g2_buf_1 _22694_ (.A(net735),
    .X(_06228_));
 sg13g2_a21oi_1 _22695_ (.A1(_00134_),
    .A2(net75),
    .Y(_06229_),
    .B1(net152));
 sg13g2_a21oi_1 _22696_ (.A1(_07681_),
    .A2(net685),
    .Y(_06230_),
    .B1(_06229_));
 sg13g2_a21oi_1 _22697_ (.A1(_06200_),
    .A2(_06227_),
    .Y(_00313_),
    .B1(_06230_));
 sg13g2_and2_1 _22698_ (.A(\top_ihp.oisc.regs[25][28] ),
    .B(net619),
    .X(_06231_));
 sg13g2_a221oi_1 _22699_ (.B2(\top_ihp.oisc.regs[30][28] ),
    .C1(_06231_),
    .B1(net576),
    .A1(\top_ihp.oisc.regs[26][28] ),
    .Y(_06232_),
    .A2(net574));
 sg13g2_a22oi_1 _22700_ (.Y(_06233_),
    .B1(_04847_),
    .B2(\top_ihp.oisc.regs[7][28] ),
    .A2(_05342_),
    .A1(\top_ihp.oisc.regs[17][28] ));
 sg13g2_mux2_1 _22701_ (.A0(\top_ihp.oisc.regs[6][28] ),
    .A1(\top_ihp.oisc.regs[2][28] ),
    .S(net654),
    .X(_06234_));
 sg13g2_a22oi_1 _22702_ (.Y(_06235_),
    .B1(_05727_),
    .B2(_06234_),
    .A2(net651),
    .A1(\top_ihp.oisc.regs[11][28] ));
 sg13g2_a22oi_1 _22703_ (.Y(_06236_),
    .B1(net469),
    .B2(\top_ihp.oisc.regs[5][28] ),
    .A2(net477),
    .A1(\top_ihp.oisc.regs[14][28] ));
 sg13g2_nand4_1 _22704_ (.B(_06233_),
    .C(_06235_),
    .A(_06232_),
    .Y(_06237_),
    .D(_06236_));
 sg13g2_a22oi_1 _22705_ (.Y(_06238_),
    .B1(net598),
    .B2(\top_ihp.oisc.regs[4][28] ),
    .A2(net465),
    .A1(\top_ihp.oisc.regs[31][28] ));
 sg13g2_a22oi_1 _22706_ (.Y(_06239_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][28] ),
    .A2(net555),
    .A1(\top_ihp.oisc.regs[29][28] ));
 sg13g2_mux2_1 _22707_ (.A0(\top_ihp.oisc.regs[3][28] ),
    .A1(\top_ihp.oisc.regs[19][28] ),
    .S(_04953_),
    .X(_06240_));
 sg13g2_a22oi_1 _22708_ (.Y(_06241_),
    .B1(_04958_),
    .B2(_06240_),
    .A2(net612),
    .A1(\top_ihp.oisc.regs[21][28] ));
 sg13g2_nand3_1 _22709_ (.B(net643),
    .C(net763),
    .A(\top_ihp.oisc.regs[24][28] ),
    .Y(_06242_));
 sg13g2_nand3_1 _22710_ (.B(net667),
    .C(net690),
    .A(\top_ihp.oisc.regs[18][28] ),
    .Y(_06243_));
 sg13g2_nand2_1 _22711_ (.Y(_06244_),
    .A(_06242_),
    .B(_06243_));
 sg13g2_a22oi_1 _22712_ (.Y(_06245_),
    .B1(_06244_),
    .B2(net556),
    .A2(net584),
    .A1(\top_ihp.oisc.regs[27][28] ));
 sg13g2_nand4_1 _22713_ (.B(_06239_),
    .C(_06241_),
    .A(_06238_),
    .Y(_06246_),
    .D(_06245_));
 sg13g2_mux2_1 _22714_ (.A0(\top_ihp.oisc.regs[20][28] ),
    .A1(\top_ihp.oisc.regs[16][28] ),
    .S(_05122_),
    .X(_06247_));
 sg13g2_a22oi_1 _22715_ (.Y(_06248_),
    .B1(_06247_),
    .B2(_05655_),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][28] ));
 sg13g2_nand2b_1 _22716_ (.Y(_06249_),
    .B(net763),
    .A_N(_06248_));
 sg13g2_a22oi_1 _22717_ (.Y(_06250_),
    .B1(_05189_),
    .B2(\top_ihp.oisc.regs[41][28] ),
    .A2(net579),
    .A1(\top_ihp.oisc.regs[48][28] ));
 sg13g2_a22oi_1 _22718_ (.Y(_06251_),
    .B1(_05401_),
    .B2(\top_ihp.oisc.regs[23][28] ),
    .A2(_04937_),
    .A1(\top_ihp.oisc.regs[1][28] ));
 sg13g2_nand2_1 _22719_ (.Y(_06252_),
    .A(\top_ihp.oisc.regs[9][28] ),
    .B(net422));
 sg13g2_nand4_1 _22720_ (.B(_06250_),
    .C(_06251_),
    .A(_06249_),
    .Y(_06253_),
    .D(_06252_));
 sg13g2_nor4_1 _22721_ (.A(net76),
    .B(_06237_),
    .C(_06246_),
    .D(_06253_),
    .Y(_06254_));
 sg13g2_a22oi_1 _22722_ (.Y(_06255_),
    .B1(_05758_),
    .B2(\top_ihp.oisc.regs[56][28] ),
    .A2(_04995_),
    .A1(\top_ihp.oisc.regs[38][28] ));
 sg13g2_a22oi_1 _22723_ (.Y(_06256_),
    .B1(_05097_),
    .B2(\top_ihp.oisc.regs[60][28] ),
    .A2(net559),
    .A1(\top_ihp.oisc.regs[51][28] ));
 sg13g2_a22oi_1 _22724_ (.Y(_06257_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[45][28] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][28] ));
 sg13g2_a22oi_1 _22725_ (.Y(_06258_),
    .B1(net457),
    .B2(\top_ihp.oisc.regs[35][28] ),
    .A2(net615),
    .A1(\top_ihp.oisc.regs[55][28] ));
 sg13g2_nand4_1 _22726_ (.B(_06256_),
    .C(_06257_),
    .A(_06255_),
    .Y(_06259_),
    .D(_06258_));
 sg13g2_a22oi_1 _22727_ (.Y(_06260_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[42][28] ),
    .A2(_05264_),
    .A1(\top_ihp.oisc.regs[53][28] ));
 sg13g2_a22oi_1 _22728_ (.Y(_06261_),
    .B1(_05309_),
    .B2(\top_ihp.oisc.regs[58][28] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][28] ));
 sg13g2_a22oi_1 _22729_ (.Y(_06262_),
    .B1(_05031_),
    .B2(\top_ihp.oisc.regs[63][28] ),
    .A2(_05359_),
    .A1(\top_ihp.oisc.regs[49][28] ));
 sg13g2_a22oi_1 _22730_ (.Y(_06263_),
    .B1(net456),
    .B2(\top_ihp.oisc.regs[46][28] ),
    .A2(_05361_),
    .A1(\top_ihp.oisc.regs[50][28] ));
 sg13g2_nand4_1 _22731_ (.B(_06261_),
    .C(_06262_),
    .A(_06260_),
    .Y(_06264_),
    .D(_06263_));
 sg13g2_a22oi_1 _22732_ (.Y(_06265_),
    .B1(_04765_),
    .B2(\top_ihp.oisc.regs[12][28] ),
    .A2(_04763_),
    .A1(\top_ihp.oisc.regs[10][28] ));
 sg13g2_nor2_1 _22733_ (.A(_04896_),
    .B(_06265_),
    .Y(_06266_));
 sg13g2_nor4_1 _22734_ (.A(net678),
    .B(net656),
    .C(net670),
    .D(net691),
    .Y(_06267_));
 sg13g2_a22oi_1 _22735_ (.Y(_06268_),
    .B1(_06267_),
    .B2(\top_ihp.oisc.regs[15][28] ),
    .A2(_04888_),
    .A1(\top_ihp.oisc.regs[13][28] ));
 sg13g2_a22oi_1 _22736_ (.Y(_06269_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[22][28] ),
    .A2(net764),
    .A1(net1028));
 sg13g2_nand2_1 _22737_ (.Y(_06270_),
    .A(_06268_),
    .B(_06269_));
 sg13g2_nor2_1 _22738_ (.A(_06266_),
    .B(_06270_),
    .Y(_06271_));
 sg13g2_a22oi_1 _22739_ (.Y(_06272_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][28] ),
    .A2(_05072_),
    .A1(\top_ihp.oisc.regs[34][28] ));
 sg13g2_a22oi_1 _22740_ (.Y(_06273_),
    .B1(_05080_),
    .B2(\top_ihp.oisc.regs[39][28] ),
    .A2(_05028_),
    .A1(\top_ihp.oisc.regs[43][28] ));
 sg13g2_a22oi_1 _22741_ (.Y(_06274_),
    .B1(_05302_),
    .B2(\top_ihp.oisc.regs[36][28] ),
    .A2(net476),
    .A1(\top_ihp.oisc.regs[47][28] ));
 sg13g2_nand4_1 _22742_ (.B(_06272_),
    .C(_06273_),
    .A(_06271_),
    .Y(_06275_),
    .D(_06274_));
 sg13g2_a22oi_1 _22743_ (.Y(_06276_),
    .B1(net413),
    .B2(\top_ihp.oisc.regs[57][28] ),
    .A2(net268),
    .A1(\top_ihp.oisc.regs[44][28] ));
 sg13g2_a22oi_1 _22744_ (.Y(_06277_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[59][28] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][28] ));
 sg13g2_a22oi_1 _22745_ (.Y(_06278_),
    .B1(_05307_),
    .B2(\top_ihp.oisc.regs[40][28] ),
    .A2(_05047_),
    .A1(\top_ihp.oisc.regs[62][28] ));
 sg13g2_a22oi_1 _22746_ (.Y(_06279_),
    .B1(_05068_),
    .B2(\top_ihp.oisc.regs[52][28] ),
    .A2(net567),
    .A1(\top_ihp.oisc.regs[61][28] ));
 sg13g2_nand4_1 _22747_ (.B(_06277_),
    .C(_06278_),
    .A(_06276_),
    .Y(_06280_),
    .D(_06279_));
 sg13g2_nor4_2 _22748_ (.A(_06259_),
    .B(_06264_),
    .C(_06275_),
    .Y(_06281_),
    .D(_06280_));
 sg13g2_a21oi_1 _22749_ (.A1(_00135_),
    .A2(net75),
    .Y(_06282_),
    .B1(net152));
 sg13g2_a21oi_1 _22750_ (.A1(_07679_),
    .A2(_06228_),
    .Y(_06283_),
    .B1(_06282_));
 sg13g2_a21oi_1 _22751_ (.A1(_06254_),
    .A2(_06281_),
    .Y(_00314_),
    .B1(_06283_));
 sg13g2_nand2_1 _22752_ (.Y(_06284_),
    .A(_07721_),
    .B(net735));
 sg13g2_a21o_1 _22753_ (.A2(_04811_),
    .A1(_00136_),
    .B1(_05105_),
    .X(_06285_));
 sg13g2_nand2_1 _22754_ (.Y(_06286_),
    .A(\top_ihp.oisc.regs[46][29] ),
    .B(net270));
 sg13g2_a22oi_1 _22755_ (.Y(_06287_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][29] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][29] ));
 sg13g2_a22oi_1 _22756_ (.Y(_06288_),
    .B1(net594),
    .B2(\top_ihp.oisc.regs[62][29] ),
    .A2(net580),
    .A1(\top_ihp.oisc.regs[42][29] ));
 sg13g2_a22oi_1 _22757_ (.Y(_06289_),
    .B1(_05590_),
    .B2(\top_ihp.oisc.regs[49][29] ),
    .A2(_05214_),
    .A1(\top_ihp.oisc.regs[54][29] ));
 sg13g2_nand4_1 _22758_ (.B(_06287_),
    .C(_06288_),
    .A(_06286_),
    .Y(_06290_),
    .D(_06289_));
 sg13g2_a22oi_1 _22759_ (.Y(_06291_),
    .B1(_05401_),
    .B2(\top_ihp.oisc.regs[23][29] ),
    .A2(_04847_),
    .A1(\top_ihp.oisc.regs[7][29] ));
 sg13g2_a22oi_1 _22760_ (.Y(_06292_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][29] ),
    .A2(_05462_),
    .A1(\top_ihp.oisc.regs[9][29] ));
 sg13g2_a22oi_1 _22761_ (.Y(_06293_),
    .B1(_04949_),
    .B2(\top_ihp.oisc.regs[28][29] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[17][29] ));
 sg13g2_mux2_1 _22762_ (.A0(\top_ihp.oisc.regs[14][29] ),
    .A1(\top_ihp.oisc.regs[6][29] ),
    .S(net642),
    .X(_06294_));
 sg13g2_nor3_1 _22763_ (.A(net652),
    .B(net656),
    .C(net719),
    .Y(_06295_));
 sg13g2_a22oi_1 _22764_ (.Y(_06296_),
    .B1(_06294_),
    .B2(_06295_),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][29] ));
 sg13g2_nand4_1 _22765_ (.B(_06292_),
    .C(_06293_),
    .A(_06291_),
    .Y(_06297_),
    .D(_06296_));
 sg13g2_mux2_1 _22766_ (.A0(\top_ihp.oisc.regs[24][29] ),
    .A1(\top_ihp.oisc.regs[16][29] ),
    .S(net667),
    .X(_06298_));
 sg13g2_a22oi_1 _22767_ (.Y(_06299_),
    .B1(_06298_),
    .B2(net556),
    .A2(_05472_),
    .A1(\top_ihp.oisc.regs[20][29] ));
 sg13g2_nand2b_1 _22768_ (.Y(_06300_),
    .B(net763),
    .A_N(_06299_));
 sg13g2_mux2_1 _22769_ (.A0(\top_ihp.oisc.regs[3][29] ),
    .A1(\top_ihp.oisc.regs[19][29] ),
    .S(_04953_),
    .X(_06301_));
 sg13g2_a22oi_1 _22770_ (.Y(_06302_),
    .B1(_04959_),
    .B2(_06301_),
    .A2(net472),
    .A1(\top_ihp.oisc.regs[29][29] ));
 sg13g2_a22oi_1 _22771_ (.Y(_06303_),
    .B1(_04937_),
    .B2(\top_ihp.oisc.regs[1][29] ),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[5][29] ));
 sg13g2_nand3_1 _22772_ (.B(_06302_),
    .C(_06303_),
    .A(_06300_),
    .Y(_06304_));
 sg13g2_nor4_1 _22773_ (.A(_05538_),
    .B(_06290_),
    .C(_06297_),
    .D(_06304_),
    .Y(_06305_));
 sg13g2_a22oi_1 _22774_ (.Y(_06306_),
    .B1(_05079_),
    .B2(\top_ihp.oisc.regs[39][29] ),
    .A2(_04988_),
    .A1(\top_ihp.oisc.regs[36][29] ));
 sg13g2_a22oi_1 _22775_ (.Y(_06307_),
    .B1(net600),
    .B2(\top_ihp.oisc.regs[2][29] ),
    .A2(_04965_),
    .A1(\top_ihp.oisc.regs[32][29] ));
 sg13g2_a22oi_1 _22776_ (.Y(_06308_),
    .B1(_05027_),
    .B2(\top_ihp.oisc.regs[43][29] ),
    .A2(_04869_),
    .A1(\top_ihp.oisc.regs[55][29] ));
 sg13g2_a22oi_1 _22777_ (.Y(_06309_),
    .B1(_05061_),
    .B2(\top_ihp.oisc.regs[57][29] ),
    .A2(_05043_),
    .A1(\top_ihp.oisc.regs[44][29] ));
 sg13g2_nand4_1 _22778_ (.B(_06307_),
    .C(_06308_),
    .A(_06306_),
    .Y(_06310_),
    .D(_06309_));
 sg13g2_a22oi_1 _22779_ (.Y(_06311_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[45][29] ),
    .A2(_05039_),
    .A1(\top_ihp.oisc.regs[50][29] ));
 sg13g2_a22oi_1 _22780_ (.Y(_06312_),
    .B1(_05088_),
    .B2(\top_ihp.oisc.regs[37][29] ),
    .A2(_04865_),
    .A1(\top_ihp.oisc.regs[53][29] ));
 sg13g2_a22oi_1 _22781_ (.Y(_06313_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[41][29] ),
    .A2(_05030_),
    .A1(\top_ihp.oisc.regs[63][29] ));
 sg13g2_a22oi_1 _22782_ (.Y(_06314_),
    .B1(_05035_),
    .B2(\top_ihp.oisc.regs[56][29] ),
    .A2(_04994_),
    .A1(\top_ihp.oisc.regs[38][29] ));
 sg13g2_nand4_1 _22783_ (.B(_06312_),
    .C(_06313_),
    .A(_06311_),
    .Y(_06315_),
    .D(_06314_));
 sg13g2_or2_1 _22784_ (.X(_06316_),
    .B(_06315_),
    .A(_06310_));
 sg13g2_a22oi_1 _22785_ (.Y(_06317_),
    .B1(net601),
    .B2(\top_ihp.oisc.regs[48][29] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][29] ));
 sg13g2_a22oi_1 _22786_ (.Y(_06318_),
    .B1(_05097_),
    .B2(\top_ihp.oisc.regs[60][29] ),
    .A2(_05179_),
    .A1(\top_ihp.oisc.regs[33][29] ));
 sg13g2_a22oi_1 _22787_ (.Y(_06319_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][29] ),
    .A2(net559),
    .A1(\top_ihp.oisc.regs[51][29] ));
 sg13g2_nand3_1 _22788_ (.B(net669),
    .C(_04722_),
    .A(\top_ihp.oisc.regs[4][29] ),
    .Y(_06320_));
 sg13g2_nand3_1 _22789_ (.B(net641),
    .C(_04972_),
    .A(\top_ihp.oisc.regs[10][29] ),
    .Y(_06321_));
 sg13g2_a21oi_1 _22790_ (.A1(_06320_),
    .A2(_06321_),
    .Y(_06322_),
    .B1(_05119_));
 sg13g2_a21oi_1 _22791_ (.A1(\top_ihp.oisc.regs[59][29] ),
    .A2(net568),
    .Y(_06323_),
    .B1(_06322_));
 sg13g2_nand4_1 _22792_ (.B(_06318_),
    .C(_06319_),
    .A(_06317_),
    .Y(_06324_),
    .D(_06323_));
 sg13g2_nand2_1 _22793_ (.Y(_06325_),
    .A(\top_ihp.oisc.regs[26][29] ),
    .B(net643));
 sg13g2_nand2_1 _22794_ (.Y(_06326_),
    .A(\top_ihp.oisc.regs[18][29] ),
    .B(net642));
 sg13g2_a21oi_1 _22795_ (.A1(_06325_),
    .A2(_06326_),
    .Y(_06327_),
    .B1(_05573_));
 sg13g2_a21oi_2 _22796_ (.B1(_06327_),
    .Y(_06328_),
    .A2(_04903_),
    .A1(\top_ihp.oisc.regs[21][29] ));
 sg13g2_a22oi_1 _22797_ (.Y(_06329_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][29] ),
    .A2(_05460_),
    .A1(\top_ihp.oisc.regs[11][29] ));
 sg13g2_a22oi_1 _22798_ (.Y(_06330_),
    .B1(net467),
    .B2(\top_ihp.oisc.regs[15][29] ),
    .A2(net473),
    .A1(\top_ihp.oisc.regs[13][29] ));
 sg13g2_a22oi_1 _22799_ (.Y(_06331_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][29] ),
    .A2(_04941_),
    .A1(\top_ihp.oisc.regs[31][29] ));
 sg13g2_nand4_1 _22800_ (.B(_06329_),
    .C(_06330_),
    .A(_06328_),
    .Y(_06332_),
    .D(_06331_));
 sg13g2_a22oi_1 _22801_ (.Y(_06333_),
    .B1(net272),
    .B2(\top_ihp.oisc.regs[34][29] ),
    .A2(net444),
    .A1(\top_ihp.oisc.regs[52][29] ));
 sg13g2_nand2_1 _22802_ (.Y(_06334_),
    .A(\top_ihp.oisc.regs[35][29] ),
    .B(net420));
 sg13g2_a22oi_1 _22803_ (.Y(_06335_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[22][29] ),
    .A2(net576),
    .A1(\top_ihp.oisc.regs[30][29] ));
 sg13g2_nand4_1 _22804_ (.B(_06333_),
    .C(_06334_),
    .A(_06284_),
    .Y(_06336_),
    .D(_06335_));
 sg13g2_nor4_1 _22805_ (.A(_06316_),
    .B(_06324_),
    .C(_06332_),
    .D(_06336_),
    .Y(_06337_));
 sg13g2_a22oi_1 _22806_ (.Y(_00315_),
    .B1(_06305_),
    .B2(_06337_),
    .A2(_06285_),
    .A1(_06284_));
 sg13g2_a22oi_1 _22807_ (.Y(_06338_),
    .B1(_05085_),
    .B2(\top_ihp.oisc.regs[40][2] ),
    .A2(_05058_),
    .A1(\top_ihp.oisc.regs[46][2] ));
 sg13g2_a22oi_1 _22808_ (.Y(_06339_),
    .B1(_05071_),
    .B2(\top_ihp.oisc.regs[34][2] ),
    .A2(_04869_),
    .A1(\top_ihp.oisc.regs[55][2] ));
 sg13g2_a22oi_1 _22809_ (.Y(_06340_),
    .B1(_05051_),
    .B2(\top_ihp.oisc.regs[61][2] ),
    .A2(_04978_),
    .A1(\top_ihp.oisc.regs[49][2] ));
 sg13g2_a22oi_1 _22810_ (.Y(_06341_),
    .B1(_05066_),
    .B2(\top_ihp.oisc.regs[52][2] ),
    .A2(_05027_),
    .A1(\top_ihp.oisc.regs[43][2] ));
 sg13g2_nand4_1 _22811_ (.B(_06339_),
    .C(_06340_),
    .A(_06338_),
    .Y(_06342_),
    .D(_06341_));
 sg13g2_a22oi_1 _22812_ (.Y(_06343_),
    .B1(net561),
    .B2(\top_ihp.oisc.regs[27][2] ),
    .A2(_04898_),
    .A1(\top_ihp.oisc.regs[10][2] ));
 sg13g2_a22oi_1 _22813_ (.Y(_06344_),
    .B1(_05015_),
    .B2(\top_ihp.oisc.regs[4][2] ),
    .A2(_04846_),
    .A1(\top_ihp.oisc.regs[7][2] ));
 sg13g2_a22oi_1 _22814_ (.Y(_06345_),
    .B1(_05254_),
    .B2(\top_ihp.oisc.regs[8][2] ),
    .A2(_05144_),
    .A1(\top_ihp.oisc.regs[17][2] ));
 sg13g2_a22oi_1 _22815_ (.Y(_06346_),
    .B1(_04901_),
    .B2(\top_ihp.oisc.regs[21][2] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][2] ));
 sg13g2_nand4_1 _22816_ (.B(_06344_),
    .C(_06345_),
    .A(_06343_),
    .Y(_06347_),
    .D(_06346_));
 sg13g2_a22oi_1 _22817_ (.Y(_06348_),
    .B1(_04940_),
    .B2(\top_ihp.oisc.regs[31][2] ),
    .A2(net613),
    .A1(\top_ihp.oisc.regs[29][2] ));
 sg13g2_a22oi_1 _22818_ (.Y(_06349_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[22][2] ),
    .A2(net554),
    .A1(\top_ihp.oisc.regs[18][2] ));
 sg13g2_a22oi_1 _22819_ (.Y(_06350_),
    .B1(net576),
    .B2(\top_ihp.oisc.regs[30][2] ),
    .A2(net772),
    .A1(_07482_));
 sg13g2_nand3_1 _22820_ (.B(_06349_),
    .C(_06350_),
    .A(_06348_),
    .Y(_06351_));
 sg13g2_nand2_1 _22821_ (.Y(_06352_),
    .A(\top_ihp.oisc.regs[36][2] ),
    .B(net462));
 sg13g2_nand2_1 _22822_ (.Y(_06353_),
    .A(\top_ihp.oisc.regs[26][2] ),
    .B(_05238_));
 sg13g2_a22oi_1 _22823_ (.Y(_06354_),
    .B1(_05245_),
    .B2(\top_ihp.oisc.regs[3][2] ),
    .A2(_05241_),
    .A1(\top_ihp.oisc.regs[19][2] ));
 sg13g2_nand3_1 _22824_ (.B(_06353_),
    .C(_06354_),
    .A(_06352_),
    .Y(_06355_));
 sg13g2_or4_1 _22825_ (.A(_06342_),
    .B(_06347_),
    .C(_06351_),
    .D(_06355_),
    .X(_06356_));
 sg13g2_a22oi_1 _22826_ (.Y(_06357_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[42][2] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[33][2] ));
 sg13g2_a22oi_1 _22827_ (.Y(_06358_),
    .B1(net434),
    .B2(\top_ihp.oisc.regs[32][2] ),
    .A2(_05191_),
    .A1(\top_ihp.oisc.regs[47][2] ));
 sg13g2_a22oi_1 _22828_ (.Y(_06359_),
    .B1(net581),
    .B2(\top_ihp.oisc.regs[51][2] ),
    .A2(_05180_),
    .A1(\top_ihp.oisc.regs[2][2] ));
 sg13g2_a22oi_1 _22829_ (.Y(_06360_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][2] ),
    .A2(_05215_),
    .A1(\top_ihp.oisc.regs[54][2] ));
 sg13g2_nand4_1 _22830_ (.B(_06358_),
    .C(_06359_),
    .A(_06357_),
    .Y(_06361_),
    .D(_06360_));
 sg13g2_a22oi_1 _22831_ (.Y(_06362_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][2] ),
    .A2(net264),
    .A1(\top_ihp.oisc.regs[45][2] ));
 sg13g2_a22oi_1 _22832_ (.Y(_06363_),
    .B1(_05188_),
    .B2(\top_ihp.oisc.regs[63][2] ),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[48][2] ));
 sg13g2_a22oi_1 _22833_ (.Y(_06364_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][2] ),
    .A2(net255),
    .A1(\top_ihp.oisc.regs[56][2] ));
 sg13g2_a22oi_1 _22834_ (.Y(_06365_),
    .B1(_05090_),
    .B2(\top_ihp.oisc.regs[37][2] ),
    .A2(net595),
    .A1(\top_ihp.oisc.regs[50][2] ));
 sg13g2_nand4_1 _22835_ (.B(_06363_),
    .C(_06364_),
    .A(_06362_),
    .Y(_06366_),
    .D(_06365_));
 sg13g2_nor3_1 _22836_ (.A(_06356_),
    .B(_06361_),
    .C(_06366_),
    .Y(_06367_));
 sg13g2_a22oi_1 _22837_ (.Y(_06368_),
    .B1(net447),
    .B2(\top_ihp.oisc.regs[35][2] ),
    .A2(_05294_),
    .A1(\top_ihp.oisc.regs[44][2] ));
 sg13g2_a22oi_1 _22838_ (.Y(_06369_),
    .B1(net568),
    .B2(\top_ihp.oisc.regs[59][2] ),
    .A2(_04920_),
    .A1(\top_ihp.oisc.regs[6][2] ));
 sg13g2_a22oi_1 _22839_ (.Y(_06370_),
    .B1(net582),
    .B2(\top_ihp.oisc.regs[62][2] ),
    .A2(net616),
    .A1(\top_ihp.oisc.regs[53][2] ));
 sg13g2_a22oi_1 _22840_ (.Y(_06371_),
    .B1(_05268_),
    .B2(\top_ihp.oisc.regs[57][2] ),
    .A2(_04984_),
    .A1(\top_ihp.oisc.regs[58][2] ));
 sg13g2_nand4_1 _22841_ (.B(_06369_),
    .C(_06370_),
    .A(_06368_),
    .Y(_06372_),
    .D(_06371_));
 sg13g2_mux2_1 _22842_ (.A0(\top_ihp.oisc.regs[24][2] ),
    .A1(\top_ihp.oisc.regs[16][2] ),
    .S(net642),
    .X(_06373_));
 sg13g2_a22oi_1 _22843_ (.Y(_06374_),
    .B1(_06373_),
    .B2(net556),
    .A2(net557),
    .A1(\top_ihp.oisc.regs[20][2] ));
 sg13g2_a22oi_1 _22844_ (.Y(_06375_),
    .B1(net267),
    .B2(\top_ihp.oisc.regs[38][2] ),
    .A2(_05485_),
    .A1(\top_ihp.oisc.regs[5][2] ));
 sg13g2_o21ai_1 _22845_ (.B1(_06375_),
    .Y(_06376_),
    .A1(net668),
    .A2(_06374_));
 sg13g2_a22oi_1 _22846_ (.Y(_06377_),
    .B1(_04927_),
    .B2(\top_ihp.oisc.regs[15][2] ),
    .A2(net473),
    .A1(\top_ihp.oisc.regs[13][2] ));
 sg13g2_a22oi_1 _22847_ (.Y(_06378_),
    .B1(net466),
    .B2(\top_ihp.oisc.regs[1][2] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][2] ));
 sg13g2_a22oi_1 _22848_ (.Y(_06379_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][2] ),
    .A2(_04949_),
    .A1(\top_ihp.oisc.regs[28][2] ));
 sg13g2_mux2_1 _22849_ (.A0(\top_ihp.oisc.regs[11][2] ),
    .A1(\top_ihp.oisc.regs[9][2] ),
    .S(net656),
    .X(_06380_));
 sg13g2_nor3_1 _22850_ (.A(net650),
    .B(net644),
    .C(net691),
    .Y(_06381_));
 sg13g2_a22oi_1 _22851_ (.Y(_06382_),
    .B1(_06380_),
    .B2(_06381_),
    .A2(_05142_),
    .A1(\top_ihp.oisc.regs[23][2] ));
 sg13g2_nand4_1 _22852_ (.B(_06378_),
    .C(_06379_),
    .A(_06377_),
    .Y(_06383_),
    .D(_06382_));
 sg13g2_nor4_1 _22853_ (.A(net78),
    .B(_06372_),
    .C(_06376_),
    .D(_06383_),
    .Y(_06384_));
 sg13g2_a21oi_1 _22854_ (.A1(_00109_),
    .A2(_06169_),
    .Y(_06385_),
    .B1(_06065_));
 sg13g2_a21oi_1 _22855_ (.A1(_07482_),
    .A2(_06228_),
    .Y(_06386_),
    .B1(_06385_));
 sg13g2_a21oi_1 _22856_ (.A1(_06367_),
    .A2(_06384_),
    .Y(_00316_),
    .B1(_06386_));
 sg13g2_a22oi_1 _22857_ (.Y(_06387_),
    .B1(net579),
    .B2(\top_ihp.oisc.regs[48][30] ),
    .A2(_05182_),
    .A1(\top_ihp.oisc.regs[42][30] ));
 sg13g2_a22oi_1 _22858_ (.Y(_06388_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][30] ),
    .A2(_05072_),
    .A1(\top_ihp.oisc.regs[34][30] ));
 sg13g2_a22oi_1 _22859_ (.Y(_06389_),
    .B1(net567),
    .B2(\top_ihp.oisc.regs[61][30] ),
    .A2(net474),
    .A1(\top_ihp.oisc.regs[33][30] ));
 sg13g2_a22oi_1 _22860_ (.Y(_06390_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[41][30] ),
    .A2(net582),
    .A1(\top_ihp.oisc.regs[62][30] ));
 sg13g2_nand4_1 _22861_ (.B(_06388_),
    .C(_06389_),
    .A(_06387_),
    .Y(_06391_),
    .D(_06390_));
 sg13g2_a22oi_1 _22862_ (.Y(_06392_),
    .B1(net595),
    .B2(\top_ihp.oisc.regs[50][30] ),
    .A2(net599),
    .A1(\top_ihp.oisc.regs[51][30] ));
 sg13g2_a22oi_1 _22863_ (.Y(_06393_),
    .B1(_05086_),
    .B2(\top_ihp.oisc.regs[40][30] ),
    .A2(net460),
    .A1(\top_ihp.oisc.regs[43][30] ));
 sg13g2_a22oi_1 _22864_ (.Y(_06394_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[45][30] ),
    .A2(_05268_),
    .A1(\top_ihp.oisc.regs[57][30] ));
 sg13g2_a22oi_1 _22865_ (.Y(_06395_),
    .B1(_05037_),
    .B2(\top_ihp.oisc.regs[56][30] ),
    .A2(net476),
    .A1(\top_ihp.oisc.regs[47][30] ));
 sg13g2_nand4_1 _22866_ (.B(_06393_),
    .C(_06394_),
    .A(_06392_),
    .Y(_06396_),
    .D(_06395_));
 sg13g2_a22oi_1 _22867_ (.Y(_06397_),
    .B1(_05127_),
    .B2(\top_ihp.oisc.regs[30][30] ),
    .A2(net797),
    .A1(\top_ihp.oisc.regs[28][30] ));
 sg13g2_nor2_1 _22868_ (.A(_04947_),
    .B(_06397_),
    .Y(_06398_));
 sg13g2_a221oi_1 _22869_ (.B2(\top_ihp.oisc.regs[22][30] ),
    .C1(_06398_),
    .B1(net552),
    .A1(\top_ihp.oisc.regs[3][30] ),
    .Y(_06399_),
    .A2(_05245_));
 sg13g2_a22oi_1 _22870_ (.Y(_06400_),
    .B1(_05241_),
    .B2(\top_ihp.oisc.regs[19][30] ),
    .A2(net574),
    .A1(\top_ihp.oisc.regs[26][30] ));
 sg13g2_a22oi_1 _22871_ (.Y(_06401_),
    .B1(_05520_),
    .B2(\top_ihp.oisc.regs[18][30] ),
    .A2(_03691_),
    .A1(net1026));
 sg13g2_mux2_1 _22872_ (.A0(\top_ihp.oisc.regs[20][30] ),
    .A1(\top_ihp.oisc.regs[16][30] ),
    .S(_04910_),
    .X(_06402_));
 sg13g2_a22oi_1 _22873_ (.Y(_06403_),
    .B1(_06402_),
    .B2(_04853_),
    .A2(_05141_),
    .A1(\top_ihp.oisc.regs[23][30] ));
 sg13g2_a22oi_1 _22874_ (.Y(_06404_),
    .B1(net584),
    .B2(\top_ihp.oisc.regs[27][30] ),
    .A2(net577),
    .A1(\top_ihp.oisc.regs[4][30] ));
 sg13g2_and2_1 _22875_ (.A(_06403_),
    .B(_06404_),
    .X(_06405_));
 sg13g2_nand4_1 _22876_ (.B(_06400_),
    .C(_06401_),
    .A(_06399_),
    .Y(_06406_),
    .D(_06405_));
 sg13g2_a22oi_1 _22877_ (.Y(_06407_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][30] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][30] ));
 sg13g2_a22oi_1 _22878_ (.Y(_06408_),
    .B1(net467),
    .B2(\top_ihp.oisc.regs[15][30] ),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][30] ));
 sg13g2_a22oi_1 _22879_ (.Y(_06409_),
    .B1(net468),
    .B2(\top_ihp.oisc.regs[6][30] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[17][30] ));
 sg13g2_a22oi_1 _22880_ (.Y(_06410_),
    .B1(net465),
    .B2(\top_ihp.oisc.regs[31][30] ),
    .A2(_04890_),
    .A1(\top_ihp.oisc.regs[13][30] ));
 sg13g2_nand4_1 _22881_ (.B(_06408_),
    .C(_06409_),
    .A(_06407_),
    .Y(_06411_),
    .D(_06410_));
 sg13g2_nor4_1 _22882_ (.A(_06391_),
    .B(_06396_),
    .C(_06406_),
    .D(_06411_),
    .Y(_06412_));
 sg13g2_a22oi_1 _22883_ (.Y(_06413_),
    .B1(_05294_),
    .B2(\top_ihp.oisc.regs[44][30] ),
    .A2(_05290_),
    .A1(\top_ihp.oisc.regs[32][30] ));
 sg13g2_a22oi_1 _22884_ (.Y(_06414_),
    .B1(net457),
    .B2(\top_ihp.oisc.regs[35][30] ),
    .A2(_04866_),
    .A1(\top_ihp.oisc.regs[53][30] ));
 sg13g2_a22oi_1 _22885_ (.Y(_06415_),
    .B1(net596),
    .B2(\top_ihp.oisc.regs[63][30] ),
    .A2(net600),
    .A1(\top_ihp.oisc.regs[2][30] ));
 sg13g2_a22oi_1 _22886_ (.Y(_06416_),
    .B1(net589),
    .B2(\top_ihp.oisc.regs[60][30] ),
    .A2(net563),
    .A1(\top_ihp.oisc.regs[49][30] ));
 sg13g2_nand4_1 _22887_ (.B(_06414_),
    .C(_06415_),
    .A(_06413_),
    .Y(_06417_),
    .D(_06416_));
 sg13g2_a22oi_1 _22888_ (.Y(_06418_),
    .B1(_05090_),
    .B2(\top_ihp.oisc.regs[37][30] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[46][30] ));
 sg13g2_a22oi_1 _22889_ (.Y(_06419_),
    .B1(net455),
    .B2(\top_ihp.oisc.regs[52][30] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][30] ));
 sg13g2_a22oi_1 _22890_ (.Y(_06420_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[36][30] ),
    .A2(_05214_),
    .A1(\top_ihp.oisc.regs[54][30] ));
 sg13g2_a22oi_1 _22891_ (.Y(_06421_),
    .B1(net568),
    .B2(\top_ihp.oisc.regs[59][30] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][30] ));
 sg13g2_nand4_1 _22892_ (.B(_06419_),
    .C(_06420_),
    .A(_06418_),
    .Y(_06422_),
    .D(_06421_));
 sg13g2_a22oi_1 _22893_ (.Y(_06423_),
    .B1(_05553_),
    .B2(\top_ihp.oisc.regs[1][30] ),
    .A2(_06111_),
    .A1(\top_ihp.oisc.regs[7][30] ));
 sg13g2_nor3_1 _22894_ (.A(net643),
    .B(net691),
    .C(_06423_),
    .Y(_06424_));
 sg13g2_a21oi_1 _22895_ (.A1(\top_ihp.oisc.regs[58][30] ),
    .A2(net442),
    .Y(_06425_),
    .B1(_06424_));
 sg13g2_mux2_1 _22896_ (.A0(\top_ihp.oisc.regs[12][30] ),
    .A1(\top_ihp.oisc.regs[8][30] ),
    .S(net678),
    .X(_06426_));
 sg13g2_a22oi_1 _22897_ (.Y(_06427_),
    .B1(_04945_),
    .B2(_06426_),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[5][30] ));
 sg13g2_a22oi_1 _22898_ (.Y(_06428_),
    .B1(net569),
    .B2(\top_ihp.oisc.regs[9][30] ),
    .A2(net471),
    .A1(\top_ihp.oisc.regs[10][30] ));
 sg13g2_and2_1 _22899_ (.A(_06427_),
    .B(_06428_),
    .X(_06429_));
 sg13g2_nand2_1 _22900_ (.Y(_06430_),
    .A(\top_ihp.oisc.regs[29][30] ),
    .B(_04894_));
 sg13g2_a22oi_1 _22901_ (.Y(_06431_),
    .B1(net470),
    .B2(\top_ihp.oisc.regs[21][30] ),
    .A2(_05320_),
    .A1(\top_ihp.oisc.regs[14][30] ));
 sg13g2_nand4_1 _22902_ (.B(_06429_),
    .C(_06430_),
    .A(_06425_),
    .Y(_06432_),
    .D(_06431_));
 sg13g2_nor4_1 _22903_ (.A(net78),
    .B(_06417_),
    .C(_06422_),
    .D(_06432_),
    .Y(_06433_));
 sg13g2_a21oi_1 _22904_ (.A1(_00137_),
    .A2(_06169_),
    .Y(_06434_),
    .B1(net152));
 sg13g2_a21oi_1 _22905_ (.A1(_07715_),
    .A2(net685),
    .Y(_06435_),
    .B1(_06434_));
 sg13g2_a21oi_1 _22906_ (.A1(_06412_),
    .A2(_06433_),
    .Y(_00317_),
    .B1(_06435_));
 sg13g2_a22oi_1 _22907_ (.Y(_06436_),
    .B1(net413),
    .B2(\top_ihp.oisc.regs[57][31] ),
    .A2(net571),
    .A1(\top_ihp.oisc.regs[63][31] ));
 sg13g2_a22oi_1 _22908_ (.Y(_06437_),
    .B1(_05297_),
    .B2(\top_ihp.oisc.regs[59][31] ),
    .A2(net572),
    .A1(\top_ihp.oisc.regs[53][31] ));
 sg13g2_a22oi_1 _22909_ (.Y(_06438_),
    .B1(net582),
    .B2(\top_ihp.oisc.regs[62][31] ),
    .A2(net562),
    .A1(\top_ihp.oisc.regs[50][31] ));
 sg13g2_a22oi_1 _22910_ (.Y(_06439_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[46][31] ),
    .A2(_05182_),
    .A1(\top_ihp.oisc.regs[42][31] ));
 sg13g2_nand4_1 _22911_ (.B(_06437_),
    .C(_06438_),
    .A(_06436_),
    .Y(_06440_),
    .D(_06439_));
 sg13g2_a22oi_1 _22912_ (.Y(_06441_),
    .B1(net421),
    .B2(\top_ihp.oisc.regs[12][31] ),
    .A2(net558),
    .A1(\top_ihp.oisc.regs[11][31] ));
 sg13g2_a22oi_1 _22913_ (.Y(_06442_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[9][31] ),
    .A2(net471),
    .A1(\top_ihp.oisc.regs[10][31] ));
 sg13g2_a22oi_1 _22914_ (.Y(_06443_),
    .B1(net468),
    .B2(\top_ihp.oisc.regs[6][31] ),
    .A2(net473),
    .A1(\top_ihp.oisc.regs[13][31] ));
 sg13g2_a22oi_1 _22915_ (.Y(_06444_),
    .B1(net465),
    .B2(\top_ihp.oisc.regs[31][31] ),
    .A2(net612),
    .A1(\top_ihp.oisc.regs[21][31] ));
 sg13g2_nand4_1 _22916_ (.B(_06442_),
    .C(_06443_),
    .A(_06441_),
    .Y(_06445_),
    .D(_06444_));
 sg13g2_mux2_1 _22917_ (.A0(\top_ihp.oisc.regs[28][31] ),
    .A1(\top_ihp.oisc.regs[20][31] ),
    .S(_05281_),
    .X(_06446_));
 sg13g2_a22oi_1 _22918_ (.Y(_06447_),
    .B1(_06446_),
    .B2(_05135_),
    .A2(_05131_),
    .A1(\top_ihp.oisc.regs[24][31] ));
 sg13g2_nand2b_1 _22919_ (.Y(_06448_),
    .B(net763),
    .A_N(_06447_));
 sg13g2_mux2_1 _22920_ (.A0(\top_ihp.oisc.regs[3][31] ),
    .A1(\top_ihp.oisc.regs[19][31] ),
    .S(net676),
    .X(_06449_));
 sg13g2_a22oi_1 _22921_ (.Y(_06450_),
    .B1(net675),
    .B2(_06449_),
    .A2(net419),
    .A1(\top_ihp.oisc.regs[5][31] ));
 sg13g2_a22oi_1 _22922_ (.Y(_06451_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][31] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][31] ));
 sg13g2_nand3_1 _22923_ (.B(_06450_),
    .C(_06451_),
    .A(_06448_),
    .Y(_06452_));
 sg13g2_nor4_1 _22924_ (.A(net76),
    .B(_06440_),
    .C(_06445_),
    .D(_06452_),
    .Y(_06453_));
 sg13g2_a22oi_1 _22925_ (.Y(_06454_),
    .B1(net259),
    .B2(\top_ihp.oisc.regs[40][31] ),
    .A2(_05164_),
    .A1(\top_ihp.oisc.regs[39][31] ));
 sg13g2_a22oi_1 _22926_ (.Y(_06455_),
    .B1(net261),
    .B2(\top_ihp.oisc.regs[44][31] ),
    .A2(net559),
    .A1(\top_ihp.oisc.regs[51][31] ));
 sg13g2_nand2_1 _22927_ (.Y(_06456_),
    .A(\top_ihp.oisc.regs[15][31] ),
    .B(net653));
 sg13g2_a22oi_1 _22928_ (.Y(_06457_),
    .B1(net552),
    .B2(\top_ihp.oisc.regs[22][31] ),
    .A2(net764),
    .A1(_08946_));
 sg13g2_a22oi_1 _22929_ (.Y(_06458_),
    .B1(net645),
    .B2(\top_ihp.oisc.regs[16][31] ),
    .A2(_05237_),
    .A1(\top_ihp.oisc.regs[26][31] ));
 sg13g2_a22oi_1 _22930_ (.Y(_06459_),
    .B1(net554),
    .B2(\top_ihp.oisc.regs[18][31] ),
    .A2(net646),
    .A1(\top_ihp.oisc.regs[30][31] ));
 sg13g2_and4_1 _22931_ (.A(_06456_),
    .B(_06457_),
    .C(_06458_),
    .D(_06459_),
    .X(_06460_));
 sg13g2_a22oi_1 _22932_ (.Y(_06461_),
    .B1(_05139_),
    .B2(\top_ihp.oisc.regs[7][31] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][31] ));
 sg13g2_a22oi_1 _22933_ (.Y(_06462_),
    .B1(_05393_),
    .B2(\top_ihp.oisc.regs[27][31] ),
    .A2(net565),
    .A1(\top_ihp.oisc.regs[1][31] ));
 sg13g2_and2_1 _22934_ (.A(_06461_),
    .B(_06462_),
    .X(_06463_));
 sg13g2_nand4_1 _22935_ (.B(_06455_),
    .C(_06460_),
    .A(_06454_),
    .Y(_06464_),
    .D(_06463_));
 sg13g2_a22oi_1 _22936_ (.Y(_06465_),
    .B1(_05077_),
    .B2(\top_ihp.oisc.regs[45][31] ),
    .A2(net566),
    .A1(\top_ihp.oisc.regs[58][31] ));
 sg13g2_a22oi_1 _22937_ (.Y(_06466_),
    .B1(_04882_),
    .B2(\top_ihp.oisc.regs[4][31] ),
    .A2(_04880_),
    .A1(\top_ihp.oisc.regs[8][31] ));
 sg13g2_nor3_1 _22938_ (.A(net677),
    .B(net719),
    .C(_06466_),
    .Y(_06467_));
 sg13g2_a21oi_1 _22939_ (.A1(\top_ihp.oisc.regs[33][31] ),
    .A2(_05179_),
    .Y(_06468_),
    .B1(_06467_));
 sg13g2_a22oi_1 _22940_ (.Y(_06469_),
    .B1(net604),
    .B2(\top_ihp.oisc.regs[49][31] ),
    .A2(net615),
    .A1(\top_ihp.oisc.regs[55][31] ));
 sg13g2_a22oi_1 _22941_ (.Y(_06470_),
    .B1(_05971_),
    .B2(\top_ihp.oisc.regs[17][31] ),
    .A2(_05609_),
    .A1(\top_ihp.oisc.regs[29][31] ));
 sg13g2_nor3_1 _22942_ (.A(_04944_),
    .B(net696),
    .C(_06470_),
    .Y(_06471_));
 sg13g2_a21oi_1 _22943_ (.A1(\top_ihp.oisc.regs[60][31] ),
    .A2(_05115_),
    .Y(_06472_),
    .B1(_06471_));
 sg13g2_nand4_1 _22944_ (.B(_06468_),
    .C(_06469_),
    .A(_06465_),
    .Y(_06473_),
    .D(_06472_));
 sg13g2_a22oi_1 _22945_ (.Y(_06474_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][31] ),
    .A2(_04970_),
    .A1(\top_ihp.oisc.regs[54][31] ));
 sg13g2_a22oi_1 _22946_ (.Y(_06475_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][31] ),
    .A2(_05055_),
    .A1(\top_ihp.oisc.regs[35][31] ));
 sg13g2_a22oi_1 _22947_ (.Y(_06476_),
    .B1(net440),
    .B2(\top_ihp.oisc.regs[2][31] ),
    .A2(_04989_),
    .A1(\top_ihp.oisc.regs[36][31] ));
 sg13g2_a22oi_1 _22948_ (.Y(_06477_),
    .B1(net455),
    .B2(\top_ihp.oisc.regs[52][31] ),
    .A2(net560),
    .A1(\top_ihp.oisc.regs[48][31] ));
 sg13g2_nand4_1 _22949_ (.B(_06475_),
    .C(_06476_),
    .A(_06474_),
    .Y(_06478_),
    .D(_06477_));
 sg13g2_nand2_1 _22950_ (.Y(_06479_),
    .A(\top_ihp.oisc.regs[56][31] ),
    .B(net255));
 sg13g2_a22oi_1 _22951_ (.Y(_06480_),
    .B1(net434),
    .B2(\top_ihp.oisc.regs[32][31] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][31] ));
 sg13g2_a22oi_1 _22952_ (.Y(_06481_),
    .B1(net269),
    .B2(\top_ihp.oisc.regs[43][31] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[38][31] ));
 sg13g2_a22oi_1 _22953_ (.Y(_06482_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][31] ),
    .A2(net567),
    .A1(\top_ihp.oisc.regs[61][31] ));
 sg13g2_nand4_1 _22954_ (.B(_06480_),
    .C(_06481_),
    .A(_06479_),
    .Y(_06483_),
    .D(_06482_));
 sg13g2_nor4_2 _22955_ (.A(_06464_),
    .B(_06473_),
    .C(_06478_),
    .Y(_06484_),
    .D(_06483_));
 sg13g2_a21oi_1 _22956_ (.A1(_00068_),
    .A2(net75),
    .Y(_06485_),
    .B1(net152));
 sg13g2_a21oi_1 _22957_ (.A1(_08946_),
    .A2(net685),
    .Y(_06486_),
    .B1(_06485_));
 sg13g2_a21oi_1 _22958_ (.A1(_06453_),
    .A2(_06484_),
    .Y(_00318_),
    .B1(_06486_));
 sg13g2_a22oi_1 _22959_ (.Y(_06487_),
    .B1(net673),
    .B2(\top_ihp.oisc.regs[8][3] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[6][3] ));
 sg13g2_nor2_1 _22960_ (.A(net688),
    .B(_06487_),
    .Y(_06488_));
 sg13g2_mux2_1 _22961_ (.A0(\top_ihp.oisc.regs[13][3] ),
    .A1(\top_ihp.oisc.regs[5][3] ),
    .S(net642),
    .X(_06489_));
 sg13g2_nand3_1 _22962_ (.B(net669),
    .C(net690),
    .A(\top_ihp.oisc.regs[30][3] ),
    .Y(_06490_));
 sg13g2_nand3_1 _22963_ (.B(net641),
    .C(net797),
    .A(\top_ihp.oisc.regs[24][3] ),
    .Y(_06491_));
 sg13g2_a21oi_2 _22964_ (.B1(_05655_),
    .Y(_06492_),
    .A2(_06491_),
    .A1(_06490_));
 sg13g2_a221oi_1 _22965_ (.B2(_06489_),
    .C1(_06492_),
    .B1(_04905_),
    .A1(\top_ihp.oisc.regs[29][3] ),
    .Y(_06493_),
    .A2(_05514_));
 sg13g2_a22oi_1 _22966_ (.Y(_06494_),
    .B1(net257),
    .B2(\top_ihp.oisc.regs[10][3] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][3] ));
 sg13g2_nand3_1 _22967_ (.B(_05134_),
    .C(net763),
    .A(\top_ihp.oisc.regs[28][3] ),
    .Y(_06495_));
 sg13g2_nand3_1 _22968_ (.B(_05464_),
    .C(net671),
    .A(\top_ihp.oisc.regs[26][3] ),
    .Y(_06496_));
 sg13g2_nand2_1 _22969_ (.Y(_06497_),
    .A(_06495_),
    .B(_06496_));
 sg13g2_a22oi_1 _22970_ (.Y(_06498_),
    .B1(_06497_),
    .B2(net643),
    .A2(net598),
    .A1(\top_ihp.oisc.regs[4][3] ));
 sg13g2_nand3_1 _22971_ (.B(_06494_),
    .C(_06498_),
    .A(_06493_),
    .Y(_06499_));
 sg13g2_a22oi_1 _22972_ (.Y(_06500_),
    .B1(_05481_),
    .B2(\top_ihp.oisc.regs[35][3] ),
    .A2(net439),
    .A1(\top_ihp.oisc.regs[63][3] ));
 sg13g2_a22oi_1 _22973_ (.Y(_06501_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][3] ),
    .A2(_05177_),
    .A1(\top_ihp.oisc.regs[58][3] ));
 sg13g2_a22oi_1 _22974_ (.Y(_06502_),
    .B1(_05116_),
    .B2(\top_ihp.oisc.regs[60][3] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[54][3] ));
 sg13g2_a22oi_1 _22975_ (.Y(_06503_),
    .B1(_05971_),
    .B2(\top_ihp.oisc.regs[2][3] ),
    .A2(net718),
    .A1(\top_ihp.oisc.regs[14][3] ));
 sg13g2_nor2_1 _22976_ (.A(_04799_),
    .B(_06503_),
    .Y(_06504_));
 sg13g2_a21oi_1 _22977_ (.A1(\top_ihp.oisc.regs[50][3] ),
    .A2(net578),
    .Y(_06505_),
    .B1(_06504_));
 sg13g2_nand4_1 _22978_ (.B(_06501_),
    .C(_06502_),
    .A(_06500_),
    .Y(_06506_),
    .D(_06505_));
 sg13g2_nor4_1 _22979_ (.A(net76),
    .B(_06488_),
    .C(_06499_),
    .D(_06506_),
    .Y(_06507_));
 sg13g2_a22oi_1 _22980_ (.Y(_06508_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[61][3] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[49][3] ));
 sg13g2_a22oi_1 _22981_ (.Y(_06509_),
    .B1(_05219_),
    .B2(\top_ihp.oisc.regs[40][3] ),
    .A2(net431),
    .A1(\top_ihp.oisc.regs[36][3] ));
 sg13g2_a22oi_1 _22982_ (.Y(_06510_),
    .B1(net255),
    .B2(\top_ihp.oisc.regs[56][3] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][3] ));
 sg13g2_a22oi_1 _22983_ (.Y(_06511_),
    .B1(net413),
    .B2(\top_ihp.oisc.regs[57][3] ),
    .A2(net599),
    .A1(\top_ihp.oisc.regs[51][3] ));
 sg13g2_nand4_1 _22984_ (.B(_06509_),
    .C(_06510_),
    .A(_06508_),
    .Y(_06512_),
    .D(_06511_));
 sg13g2_a22oi_1 _22985_ (.Y(_06513_),
    .B1(net270),
    .B2(\top_ihp.oisc.regs[46][3] ),
    .A2(_05109_),
    .A1(\top_ihp.oisc.regs[55][3] ));
 sg13g2_a22oi_1 _22986_ (.Y(_06514_),
    .B1(net553),
    .B2(\top_ihp.oisc.regs[62][3] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[38][3] ));
 sg13g2_a22oi_1 _22987_ (.Y(_06515_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[42][3] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][3] ));
 sg13g2_a22oi_1 _22988_ (.Y(_06516_),
    .B1(net271),
    .B2(\top_ihp.oisc.regs[37][3] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[43][3] ));
 sg13g2_nand4_1 _22989_ (.B(_06514_),
    .C(_06515_),
    .A(_06513_),
    .Y(_06517_),
    .D(_06516_));
 sg13g2_a22oi_1 _22990_ (.Y(_06518_),
    .B1(_05066_),
    .B2(\top_ihp.oisc.regs[52][3] ),
    .A2(_04998_),
    .A1(\top_ihp.oisc.regs[59][3] ));
 sg13g2_a22oi_1 _22991_ (.Y(_06519_),
    .B1(_04965_),
    .B2(\top_ihp.oisc.regs[32][3] ),
    .A2(_04843_),
    .A1(\top_ihp.oisc.regs[47][3] ));
 sg13g2_a22oi_1 _22992_ (.Y(_06520_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[41][3] ),
    .A2(_05043_),
    .A1(\top_ihp.oisc.regs[44][3] ));
 sg13g2_a22oi_1 _22993_ (.Y(_06521_),
    .B1(_05071_),
    .B2(\top_ihp.oisc.regs[34][3] ),
    .A2(_05003_),
    .A1(\top_ihp.oisc.regs[48][3] ));
 sg13g2_nand4_1 _22994_ (.B(_06519_),
    .C(_06520_),
    .A(_06518_),
    .Y(_06522_),
    .D(_06521_));
 sg13g2_nand2_1 _22995_ (.Y(_06523_),
    .A(\top_ihp.oisc.regs[45][3] ),
    .B(net438));
 sg13g2_a22oi_1 _22996_ (.Y(_06524_),
    .B1(net554),
    .B2(\top_ihp.oisc.regs[18][3] ),
    .A2(net645),
    .A1(\top_ihp.oisc.regs[16][3] ));
 sg13g2_a22oi_1 _22997_ (.Y(_06525_),
    .B1(net721),
    .B2(\top_ihp.oisc.regs[22][3] ),
    .A2(net722),
    .A1(\top_ihp.oisc.regs[20][3] ));
 sg13g2_nor2_1 _22998_ (.A(net672),
    .B(_06525_),
    .Y(_06526_));
 sg13g2_a21oi_1 _22999_ (.A1(\top_ihp.oisc.regs[19][3] ),
    .A2(_05241_),
    .Y(_06527_),
    .B1(_06526_));
 sg13g2_nand3_1 _23000_ (.B(_06524_),
    .C(_06527_),
    .A(_06523_),
    .Y(_06528_));
 sg13g2_nand2_1 _23001_ (.Y(_06529_),
    .A(\top_ihp.oisc.regs[27][3] ),
    .B(net584));
 sg13g2_a22oi_1 _23002_ (.Y(_06530_),
    .B1(_05245_),
    .B2(\top_ihp.oisc.regs[3][3] ),
    .A2(net772),
    .A1(_07496_));
 sg13g2_a22oi_1 _23003_ (.Y(_06531_),
    .B1(net607),
    .B2(\top_ihp.oisc.regs[31][3] ),
    .A2(net653),
    .A1(\top_ihp.oisc.regs[15][3] ));
 sg13g2_nand3_1 _23004_ (.B(_06530_),
    .C(_06531_),
    .A(_06529_),
    .Y(_06532_));
 sg13g2_a22oi_1 _23005_ (.Y(_06533_),
    .B1(net569),
    .B2(\top_ihp.oisc.regs[9][3] ),
    .A2(net565),
    .A1(\top_ihp.oisc.regs[1][3] ));
 sg13g2_a22oi_1 _23006_ (.Y(_06534_),
    .B1(net651),
    .B2(\top_ihp.oisc.regs[11][3] ),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][3] ));
 sg13g2_a22oi_1 _23007_ (.Y(_06535_),
    .B1(net585),
    .B2(\top_ihp.oisc.regs[12][3] ),
    .A2(net618),
    .A1(\top_ihp.oisc.regs[17][3] ));
 sg13g2_a22oi_1 _23008_ (.Y(_06536_),
    .B1(net648),
    .B2(\top_ihp.oisc.regs[23][3] ),
    .A2(net649),
    .A1(\top_ihp.oisc.regs[7][3] ));
 sg13g2_nand4_1 _23009_ (.B(_06534_),
    .C(_06535_),
    .A(_06533_),
    .Y(_06537_),
    .D(_06536_));
 sg13g2_or4_1 _23010_ (.A(_06522_),
    .B(_06528_),
    .C(_06532_),
    .D(_06537_),
    .X(_06538_));
 sg13g2_nor3_1 _23011_ (.A(_06512_),
    .B(_06517_),
    .C(_06538_),
    .Y(_06539_));
 sg13g2_a21oi_1 _23012_ (.A1(_00110_),
    .A2(net75),
    .Y(_06540_),
    .B1(net152));
 sg13g2_a21oi_1 _23013_ (.A1(_07496_),
    .A2(net685),
    .Y(_06541_),
    .B1(_06540_));
 sg13g2_a21oi_1 _23014_ (.A1(_06507_),
    .A2(_06539_),
    .Y(_00319_),
    .B1(_06541_));
 sg13g2_a22oi_1 _23015_ (.Y(_06542_),
    .B1(net590),
    .B2(\top_ihp.oisc.regs[60][4] ),
    .A2(net560),
    .A1(\top_ihp.oisc.regs[48][4] ));
 sg13g2_a22oi_1 _23016_ (.Y(_06543_),
    .B1(_05485_),
    .B2(\top_ihp.oisc.regs[5][4] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[33][4] ));
 sg13g2_a22oi_1 _23017_ (.Y(_06544_),
    .B1(net562),
    .B2(\top_ihp.oisc.regs[50][4] ),
    .A2(net459),
    .A1(\top_ihp.oisc.regs[56][4] ));
 sg13g2_a22oi_1 _23018_ (.Y(_06545_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[36][4] ),
    .A2(_04870_),
    .A1(\top_ihp.oisc.regs[55][4] ));
 sg13g2_nand4_1 _23019_ (.B(_06543_),
    .C(_06544_),
    .A(_06542_),
    .Y(_06546_),
    .D(_06545_));
 sg13g2_a22oi_1 _23020_ (.Y(_06547_),
    .B1(net673),
    .B2(\top_ihp.oisc.regs[8][4] ),
    .A2(net674),
    .A1(\top_ihp.oisc.regs[6][4] ));
 sg13g2_a22oi_1 _23021_ (.Y(_06548_),
    .B1(net553),
    .B2(\top_ihp.oisc.regs[62][4] ),
    .A2(net267),
    .A1(\top_ihp.oisc.regs[38][4] ));
 sg13g2_o21ai_1 _23022_ (.B1(_06548_),
    .Y(_06549_),
    .A1(net688),
    .A2(_06547_));
 sg13g2_a22oi_1 _23023_ (.Y(_06550_),
    .B1(net472),
    .B2(\top_ihp.oisc.regs[29][4] ),
    .A2(net418),
    .A1(\top_ihp.oisc.regs[25][4] ));
 sg13g2_a22oi_1 _23024_ (.Y(_06551_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][4] ),
    .A2(net257),
    .A1(\top_ihp.oisc.regs[10][4] ));
 sg13g2_mux2_1 _23025_ (.A0(\top_ihp.oisc.regs[3][4] ),
    .A1(\top_ihp.oisc.regs[19][4] ),
    .S(net676),
    .X(_06552_));
 sg13g2_a22oi_1 _23026_ (.Y(_06553_),
    .B1(net675),
    .B2(_06552_),
    .A2(net470),
    .A1(\top_ihp.oisc.regs[21][4] ));
 sg13g2_mux2_1 _23027_ (.A0(\top_ihp.oisc.regs[30][4] ),
    .A1(\top_ihp.oisc.regs[22][4] ),
    .S(net642),
    .X(_06554_));
 sg13g2_and2_1 _23028_ (.A(_04741_),
    .B(net671),
    .X(_06555_));
 sg13g2_nand3_1 _23029_ (.B(_05409_),
    .C(net671),
    .A(\top_ihp.oisc.regs[26][4] ),
    .Y(_06556_));
 sg13g2_nand3_1 _23030_ (.B(_05412_),
    .C(_05410_),
    .A(\top_ihp.oisc.regs[16][4] ),
    .Y(_06557_));
 sg13g2_nand2_1 _23031_ (.Y(_06558_),
    .A(_06556_),
    .B(_06557_));
 sg13g2_a22oi_1 _23032_ (.Y(_06559_),
    .B1(_06558_),
    .B2(_05474_),
    .A2(_06555_),
    .A1(_06554_));
 sg13g2_nand4_1 _23033_ (.B(_06551_),
    .C(_06553_),
    .A(_06550_),
    .Y(_06560_),
    .D(_06559_));
 sg13g2_nor4_1 _23034_ (.A(net80),
    .B(_06546_),
    .C(_06549_),
    .D(_06560_),
    .Y(_06561_));
 sg13g2_a22oi_1 _23035_ (.Y(_06562_),
    .B1(_05591_),
    .B2(\top_ihp.oisc.regs[37][4] ),
    .A2(_05086_),
    .A1(\top_ihp.oisc.regs[40][4] ));
 sg13g2_a22oi_1 _23036_ (.Y(_06563_),
    .B1(_05031_),
    .B2(\top_ihp.oisc.regs[63][4] ),
    .A2(net602),
    .A1(\top_ihp.oisc.regs[59][4] ));
 sg13g2_a22oi_1 _23037_ (.Y(_06564_),
    .B1(net454),
    .B2(\top_ihp.oisc.regs[34][4] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][4] ));
 sg13g2_a22oi_1 _23038_ (.Y(_06565_),
    .B1(_05059_),
    .B2(\top_ihp.oisc.regs[46][4] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][4] ));
 sg13g2_nand4_1 _23039_ (.B(_06563_),
    .C(_06564_),
    .A(_06562_),
    .Y(_06566_),
    .D(_06565_));
 sg13g2_a22oi_1 _23040_ (.Y(_06567_),
    .B1(net452),
    .B2(\top_ihp.oisc.regs[39][4] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[43][4] ));
 sg13g2_a22oi_1 _23041_ (.Y(_06568_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[41][4] ),
    .A2(_05054_),
    .A1(\top_ihp.oisc.regs[35][4] ));
 sg13g2_a22oi_1 _23042_ (.Y(_06569_),
    .B1(_04979_),
    .B2(\top_ihp.oisc.regs[49][4] ),
    .A2(_04866_),
    .A1(\top_ihp.oisc.regs[53][4] ));
 sg13g2_a22oi_1 _23043_ (.Y(_06570_),
    .B1(net440),
    .B2(\top_ihp.oisc.regs[2][4] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][4] ));
 sg13g2_nand4_1 _23044_ (.B(_06568_),
    .C(_06569_),
    .A(_06567_),
    .Y(_06571_),
    .D(_06570_));
 sg13g2_a22oi_1 _23045_ (.Y(_06572_),
    .B1(net268),
    .B2(\top_ihp.oisc.regs[44][4] ),
    .A2(_05597_),
    .A1(\top_ihp.oisc.regs[47][4] ));
 sg13g2_a22oi_1 _23046_ (.Y(_06573_),
    .B1(net453),
    .B2(\top_ihp.oisc.regs[45][4] ),
    .A2(net570),
    .A1(\top_ihp.oisc.regs[57][4] ));
 sg13g2_a22oi_1 _23047_ (.Y(_06574_),
    .B1(net567),
    .B2(\top_ihp.oisc.regs[61][4] ),
    .A2(net559),
    .A1(\top_ihp.oisc.regs[51][4] ));
 sg13g2_a22oi_1 _23048_ (.Y(_06575_),
    .B1(_05067_),
    .B2(\top_ihp.oisc.regs[52][4] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[58][4] ));
 sg13g2_nand4_1 _23049_ (.B(_06573_),
    .C(_06574_),
    .A(_06572_),
    .Y(_06576_),
    .D(_06575_));
 sg13g2_nand2_1 _23050_ (.Y(_06577_),
    .A(_07487_),
    .B(net764));
 sg13g2_a22oi_1 _23051_ (.Y(_06578_),
    .B1(net554),
    .B2(\top_ihp.oisc.regs[18][4] ),
    .A2(_04855_),
    .A1(\top_ihp.oisc.regs[20][4] ));
 sg13g2_nand2_1 _23052_ (.Y(_06579_),
    .A(_06577_),
    .B(_06578_));
 sg13g2_a221oi_1 _23053_ (.B2(\top_ihp.oisc.regs[11][4] ),
    .C1(_06579_),
    .B1(net651),
    .A1(\top_ihp.oisc.regs[24][4] ),
    .Y(_06580_),
    .A2(net658));
 sg13g2_a22oi_1 _23054_ (.Y(_06581_),
    .B1(net598),
    .B2(\top_ihp.oisc.regs[4][4] ),
    .A2(net466),
    .A1(\top_ihp.oisc.regs[1][4] ));
 sg13g2_a22oi_1 _23055_ (.Y(_06582_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[9][4] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][4] ));
 sg13g2_a22oi_1 _23056_ (.Y(_06583_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[15][4] ),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][4] ));
 sg13g2_a22oi_1 _23057_ (.Y(_06584_),
    .B1(net648),
    .B2(\top_ihp.oisc.regs[23][4] ),
    .A2(net655),
    .A1(\top_ihp.oisc.regs[13][4] ));
 sg13g2_a22oi_1 _23058_ (.Y(_06585_),
    .B1(net585),
    .B2(\top_ihp.oisc.regs[12][4] ),
    .A2(net573),
    .A1(\top_ihp.oisc.regs[31][4] ));
 sg13g2_a22oi_1 _23059_ (.Y(_06586_),
    .B1(_04948_),
    .B2(\top_ihp.oisc.regs[28][4] ),
    .A2(net657),
    .A1(\top_ihp.oisc.regs[7][4] ));
 sg13g2_and4_1 _23060_ (.A(_06583_),
    .B(_06584_),
    .C(_06585_),
    .D(_06586_),
    .X(_06587_));
 sg13g2_nand4_1 _23061_ (.B(_06581_),
    .C(_06582_),
    .A(_06580_),
    .Y(_06588_),
    .D(_06587_));
 sg13g2_nor4_2 _23062_ (.A(_06566_),
    .B(_06571_),
    .C(_06576_),
    .Y(_06589_),
    .D(_06588_));
 sg13g2_a21o_1 _23063_ (.A2(net79),
    .A1(_00111_),
    .B1(net154),
    .X(_06590_));
 sg13g2_a22oi_1 _23064_ (.Y(_00320_),
    .B1(_06590_),
    .B2(_06577_),
    .A2(_06589_),
    .A1(_06561_));
 sg13g2_nand2_1 _23065_ (.Y(_06591_),
    .A(\top_ihp.oisc.regs[48][5] ),
    .B(_05004_));
 sg13g2_a22oi_1 _23066_ (.Y(_06592_),
    .B1(_05077_),
    .B2(\top_ihp.oisc.regs[45][5] ),
    .A2(_05299_),
    .A1(\top_ihp.oisc.regs[61][5] ));
 sg13g2_and2_1 _23067_ (.A(\top_ihp.oisc.regs[6][5] ),
    .B(net610),
    .X(_06593_));
 sg13g2_a221oi_1 _23068_ (.B2(\top_ihp.oisc.regs[5][5] ),
    .C1(_06593_),
    .B1(net611),
    .A1(\top_ihp.oisc.regs[55][5] ),
    .Y(_06594_),
    .A2(net615));
 sg13g2_a22oi_1 _23069_ (.Y(_06595_),
    .B1(net592),
    .B2(\top_ihp.oisc.regs[57][5] ),
    .A2(_05424_),
    .A1(\top_ihp.oisc.regs[51][5] ));
 sg13g2_nand4_1 _23070_ (.B(_06592_),
    .C(_06594_),
    .A(_06591_),
    .Y(_06596_),
    .D(_06595_));
 sg13g2_a22oi_1 _23071_ (.Y(_06597_),
    .B1(net465),
    .B2(\top_ihp.oisc.regs[31][5] ),
    .A2(net617),
    .A1(\top_ihp.oisc.regs[7][5] ));
 sg13g2_a22oi_1 _23072_ (.Y(_06598_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][5] ),
    .A2(net569),
    .A1(\top_ihp.oisc.regs[9][5] ));
 sg13g2_mux2_1 _23073_ (.A0(\top_ihp.oisc.regs[3][5] ),
    .A1(\top_ihp.oisc.regs[19][5] ),
    .S(net676),
    .X(_06599_));
 sg13g2_a22oi_1 _23074_ (.Y(_06600_),
    .B1(net692),
    .B2(_06599_),
    .A2(net473),
    .A1(\top_ihp.oisc.regs[13][5] ));
 sg13g2_a22oi_1 _23075_ (.Y(_06601_),
    .B1(net598),
    .B2(\top_ihp.oisc.regs[4][5] ),
    .A2(net564),
    .A1(\top_ihp.oisc.regs[25][5] ));
 sg13g2_nand4_1 _23076_ (.B(_06598_),
    .C(_06600_),
    .A(_06597_),
    .Y(_06602_),
    .D(_06601_));
 sg13g2_a22oi_1 _23077_ (.Y(_06603_),
    .B1(net467),
    .B2(\top_ihp.oisc.regs[15][5] ),
    .A2(net257),
    .A1(\top_ihp.oisc.regs[10][5] ));
 sg13g2_nand2_1 _23078_ (.Y(_06604_),
    .A(\top_ihp.oisc.regs[17][5] ),
    .B(net429));
 sg13g2_mux2_1 _23079_ (.A0(\top_ihp.oisc.regs[12][5] ),
    .A1(\top_ihp.oisc.regs[8][5] ),
    .S(net654),
    .X(_06605_));
 sg13g2_a22oi_1 _23080_ (.Y(_06606_),
    .B1(_04945_),
    .B2(_06605_),
    .A2(net466),
    .A1(\top_ihp.oisc.regs[1][5] ));
 sg13g2_a22oi_1 _23081_ (.Y(_06607_),
    .B1(net464),
    .B2(\top_ihp.oisc.regs[28][5] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][5] ));
 sg13g2_nand4_1 _23082_ (.B(_06604_),
    .C(_06606_),
    .A(_06603_),
    .Y(_06608_),
    .D(_06607_));
 sg13g2_nor4_1 _23083_ (.A(net76),
    .B(_06596_),
    .C(_06602_),
    .D(_06608_),
    .Y(_06609_));
 sg13g2_a22oi_1 _23084_ (.Y(_06610_),
    .B1(net578),
    .B2(\top_ihp.oisc.regs[50][5] ),
    .A2(_05290_),
    .A1(\top_ihp.oisc.regs[32][5] ));
 sg13g2_a22oi_1 _23085_ (.Y(_06611_),
    .B1(_05094_),
    .B2(\top_ihp.oisc.regs[41][5] ),
    .A2(net458),
    .A1(\top_ihp.oisc.regs[44][5] ));
 sg13g2_a22oi_1 _23086_ (.Y(_06612_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[39][5] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][5] ));
 sg13g2_a22oi_1 _23087_ (.Y(_06613_),
    .B1(_04882_),
    .B2(\top_ihp.oisc.regs[20][5] ),
    .A2(_04880_),
    .A1(\top_ihp.oisc.regs[24][5] ));
 sg13g2_nor2_1 _23088_ (.A(_05130_),
    .B(_06613_),
    .Y(_06614_));
 sg13g2_a21oi_1 _23089_ (.A1(\top_ihp.oisc.regs[33][5] ),
    .A2(_04876_),
    .Y(_06615_),
    .B1(_06614_));
 sg13g2_nand4_1 _23090_ (.B(_06611_),
    .C(_06612_),
    .A(_06610_),
    .Y(_06616_),
    .D(_06615_));
 sg13g2_a22oi_1 _23091_ (.Y(_06617_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[36][5] ),
    .A2(net415),
    .A1(\top_ihp.oisc.regs[47][5] ));
 sg13g2_a22oi_1 _23092_ (.Y(_06618_),
    .B1(net416),
    .B2(\top_ihp.oisc.regs[37][5] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][5] ));
 sg13g2_a22oi_1 _23093_ (.Y(_06619_),
    .B1(net647),
    .B2(\top_ihp.oisc.regs[11][5] ),
    .A2(net613),
    .A1(\top_ihp.oisc.regs[29][5] ));
 sg13g2_a22oi_1 _23094_ (.Y(_06620_),
    .B1(net587),
    .B2(\top_ihp.oisc.regs[23][5] ),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][5] ));
 sg13g2_and2_1 _23095_ (.A(_06619_),
    .B(_06620_),
    .X(_06621_));
 sg13g2_a22oi_1 _23096_ (.Y(_06622_),
    .B1(_05705_),
    .B2(\top_ihp.oisc.regs[22][5] ),
    .A2(_05202_),
    .A1(_07490_));
 sg13g2_inv_1 _23097_ (.Y(_06623_),
    .A(_06622_));
 sg13g2_a221oi_1 _23098_ (.B2(\top_ihp.oisc.regs[30][5] ),
    .C1(_06623_),
    .B1(net576),
    .A1(\top_ihp.oisc.regs[49][5] ),
    .Y(_06624_),
    .A2(net563));
 sg13g2_nand4_1 _23099_ (.B(_06618_),
    .C(_06621_),
    .A(_06617_),
    .Y(_06625_),
    .D(_06624_));
 sg13g2_a22oi_1 _23100_ (.Y(_06626_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][5] ),
    .A2(net571),
    .A1(\top_ihp.oisc.regs[63][5] ));
 sg13g2_a22oi_1 _23101_ (.Y(_06627_),
    .B1(_05047_),
    .B2(\top_ihp.oisc.regs[62][5] ),
    .A2(_05309_),
    .A1(\top_ihp.oisc.regs[58][5] ));
 sg13g2_a22oi_1 _23102_ (.Y(_06628_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][5] ),
    .A2(_05009_),
    .A1(\top_ihp.oisc.regs[2][5] ));
 sg13g2_a22oi_1 _23103_ (.Y(_06629_),
    .B1(net273),
    .B2(\top_ihp.oisc.regs[56][5] ),
    .A2(net461),
    .A1(\top_ihp.oisc.regs[38][5] ));
 sg13g2_nand4_1 _23104_ (.B(_06627_),
    .C(_06628_),
    .A(_06626_),
    .Y(_06630_),
    .D(_06629_));
 sg13g2_nand3_1 _23105_ (.B(_05409_),
    .C(net690),
    .A(\top_ihp.oisc.regs[26][5] ),
    .Y(_06631_));
 sg13g2_nand3_1 _23106_ (.B(_05412_),
    .C(net763),
    .A(\top_ihp.oisc.regs[16][5] ),
    .Y(_06632_));
 sg13g2_nand2_1 _23107_ (.Y(_06633_),
    .A(\top_ihp.oisc.regs[18][5] ),
    .B(_04917_));
 sg13g2_nand3_1 _23108_ (.B(_06632_),
    .C(_06633_),
    .A(_06631_),
    .Y(_06634_));
 sg13g2_a22oi_1 _23109_ (.Y(_06635_),
    .B1(_06634_),
    .B2(_05474_),
    .A2(_05297_),
    .A1(\top_ihp.oisc.regs[59][5] ));
 sg13g2_a22oi_1 _23110_ (.Y(_06636_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][5] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[46][5] ));
 sg13g2_a22oi_1 _23111_ (.Y(_06637_),
    .B1(net455),
    .B2(\top_ihp.oisc.regs[52][5] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][5] ));
 sg13g2_a22oi_1 _23112_ (.Y(_06638_),
    .B1(net420),
    .B2(\top_ihp.oisc.regs[35][5] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[43][5] ));
 sg13g2_nand4_1 _23113_ (.B(_06636_),
    .C(_06637_),
    .A(_06635_),
    .Y(_06639_),
    .D(_06638_));
 sg13g2_nor4_2 _23114_ (.A(_06616_),
    .B(_06625_),
    .C(_06630_),
    .Y(_06640_),
    .D(_06639_));
 sg13g2_a21oi_1 _23115_ (.A1(_00112_),
    .A2(net75),
    .Y(_06641_),
    .B1(net152));
 sg13g2_a21oi_1 _23116_ (.A1(_07490_),
    .A2(net685),
    .Y(_06642_),
    .B1(_06641_));
 sg13g2_a21oi_1 _23117_ (.A1(_06609_),
    .A2(_06640_),
    .Y(_00321_),
    .B1(_06642_));
 sg13g2_a22oi_1 _23118_ (.Y(_06643_),
    .B1(net256),
    .B2(\top_ihp.oisc.regs[34][6] ),
    .A2(net457),
    .A1(\top_ihp.oisc.regs[35][6] ));
 sg13g2_a22oi_1 _23119_ (.Y(_06644_),
    .B1(_05037_),
    .B2(\top_ihp.oisc.regs[56][6] ),
    .A2(_05398_),
    .A1(\top_ihp.oisc.regs[48][6] ));
 sg13g2_a22oi_1 _23120_ (.Y(_06645_),
    .B1(_05089_),
    .B2(\top_ihp.oisc.regs[37][6] ),
    .A2(net593),
    .A1(\top_ihp.oisc.regs[61][6] ));
 sg13g2_a22oi_1 _23121_ (.Y(_06646_),
    .B1(_05062_),
    .B2(\top_ihp.oisc.regs[57][6] ),
    .A2(_04966_),
    .A1(\top_ihp.oisc.regs[32][6] ));
 sg13g2_nand4_1 _23122_ (.B(_06644_),
    .C(_06645_),
    .A(_06643_),
    .Y(_06647_),
    .D(_06646_));
 sg13g2_a22oi_1 _23123_ (.Y(_06648_),
    .B1(net260),
    .B2(\top_ihp.oisc.regs[41][6] ),
    .A2(_05597_),
    .A1(\top_ihp.oisc.regs[47][6] ));
 sg13g2_a22oi_1 _23124_ (.Y(_06649_),
    .B1(net455),
    .B2(\top_ihp.oisc.regs[52][6] ),
    .A2(net606),
    .A1(\top_ihp.oisc.regs[54][6] ));
 sg13g2_a22oi_1 _23125_ (.Y(_06650_),
    .B1(_05012_),
    .B2(\top_ihp.oisc.regs[51][6] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][6] ));
 sg13g2_a22oi_1 _23126_ (.Y(_06651_),
    .B1(_05192_),
    .B2(\top_ihp.oisc.regs[45][6] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[42][6] ));
 sg13g2_nand4_1 _23127_ (.B(_06649_),
    .C(_06650_),
    .A(_06648_),
    .Y(_06652_),
    .D(_06651_));
 sg13g2_mux2_1 _23128_ (.A0(\top_ihp.oisc.regs[3][6] ),
    .A1(\top_ihp.oisc.regs[19][6] ),
    .S(net693),
    .X(_06653_));
 sg13g2_a22oi_1 _23129_ (.Y(_06654_),
    .B1(_06653_),
    .B2(net692),
    .A2(net577),
    .A1(\top_ihp.oisc.regs[4][6] ));
 sg13g2_a22oi_1 _23130_ (.Y(_06655_),
    .B1(net585),
    .B2(\top_ihp.oisc.regs[12][6] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][6] ));
 sg13g2_a22oi_1 _23131_ (.Y(_06656_),
    .B1(net565),
    .B2(\top_ihp.oisc.regs[1][6] ),
    .A2(_04898_),
    .A1(\top_ihp.oisc.regs[10][6] ));
 sg13g2_a22oi_1 _23132_ (.Y(_06657_),
    .B1(net647),
    .B2(\top_ihp.oisc.regs[11][6] ),
    .A2(net573),
    .A1(\top_ihp.oisc.regs[31][6] ));
 sg13g2_and4_1 _23133_ (.A(_06654_),
    .B(_06655_),
    .C(_06656_),
    .D(_06657_),
    .X(_06658_));
 sg13g2_nand2_1 _23134_ (.Y(_06659_),
    .A(\top_ihp.oisc.regs[36][6] ),
    .B(net262));
 sg13g2_a22oi_1 _23135_ (.Y(_06660_),
    .B1(_05620_),
    .B2(\top_ihp.oisc.regs[62][6] ),
    .A2(_05185_),
    .A1(\top_ihp.oisc.regs[50][6] ));
 sg13g2_nand3_1 _23136_ (.B(_06659_),
    .C(_06660_),
    .A(_06658_),
    .Y(_06661_));
 sg13g2_a22oi_1 _23137_ (.Y(_06662_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][6] ),
    .A2(net268),
    .A1(\top_ihp.oisc.regs[44][6] ));
 sg13g2_a22oi_1 _23138_ (.Y(_06663_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[39][6] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[49][6] ));
 sg13g2_a22oi_1 _23139_ (.Y(_06664_),
    .B1(net270),
    .B2(\top_ihp.oisc.regs[46][6] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[43][6] ));
 sg13g2_a22oi_1 _23140_ (.Y(_06665_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[58][6] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[53][6] ));
 sg13g2_nand4_1 _23141_ (.B(_06663_),
    .C(_06664_),
    .A(_06662_),
    .Y(_06666_),
    .D(_06665_));
 sg13g2_nor4_2 _23142_ (.A(_06647_),
    .B(_06652_),
    .C(_06661_),
    .Y(_06667_),
    .D(_06666_));
 sg13g2_and2_1 _23143_ (.A(\top_ihp.oisc.regs[30][6] ),
    .B(net576),
    .X(_06668_));
 sg13g2_a221oi_1 _23144_ (.B2(\top_ihp.oisc.regs[18][6] ),
    .C1(_06668_),
    .B1(_05520_),
    .A1(\top_ihp.oisc.regs[5][6] ),
    .Y(_06669_),
    .A2(net611));
 sg13g2_a22oi_1 _23145_ (.Y(_06670_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[9][6] ),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][6] ));
 sg13g2_a22oi_1 _23146_ (.Y(_06671_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[8][6] ),
    .A2(net612),
    .A1(\top_ihp.oisc.regs[21][6] ));
 sg13g2_a22oi_1 _23147_ (.Y(_06672_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[15][6] ),
    .A2(net618),
    .A1(\top_ihp.oisc.regs[17][6] ));
 sg13g2_nand4_1 _23148_ (.B(_06670_),
    .C(_06671_),
    .A(_06669_),
    .Y(_06673_),
    .D(_06672_));
 sg13g2_nand2_1 _23149_ (.Y(_06674_),
    .A(\top_ihp.oisc.regs[28][6] ),
    .B(net464));
 sg13g2_a22oi_1 _23150_ (.Y(_06675_),
    .B1(net472),
    .B2(\top_ihp.oisc.regs[29][6] ),
    .A2(net617),
    .A1(\top_ihp.oisc.regs[7][6] ));
 sg13g2_a22oi_1 _23151_ (.Y(_06676_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[27][6] ),
    .A2(net587),
    .A1(\top_ihp.oisc.regs[23][6] ));
 sg13g2_nand3_1 _23152_ (.B(_05134_),
    .C(net690),
    .A(\top_ihp.oisc.regs[22][6] ),
    .Y(_06677_));
 sg13g2_nand3_1 _23153_ (.B(_05464_),
    .C(_04851_),
    .A(\top_ihp.oisc.regs[16][6] ),
    .Y(_06678_));
 sg13g2_nand2_1 _23154_ (.Y(_06679_),
    .A(_06677_),
    .B(_06678_));
 sg13g2_a22oi_1 _23155_ (.Y(_06680_),
    .B1(_06679_),
    .B2(net640),
    .A2(net610),
    .A1(\top_ihp.oisc.regs[6][6] ));
 sg13g2_nand4_1 _23156_ (.B(_06675_),
    .C(_06676_),
    .A(_06674_),
    .Y(_06681_),
    .D(_06680_));
 sg13g2_a22oi_1 _23157_ (.Y(_06682_),
    .B1(_05472_),
    .B2(\top_ihp.oisc.regs[20][6] ),
    .A2(_04880_),
    .A1(\top_ihp.oisc.regs[24][6] ));
 sg13g2_and2_1 _23158_ (.A(net1031),
    .B(net803),
    .X(_06683_));
 sg13g2_a221oi_1 _23159_ (.B2(\top_ihp.oisc.regs[26][6] ),
    .C1(_06683_),
    .B1(_05237_),
    .A1(\top_ihp.oisc.regs[14][6] ),
    .Y(_06684_),
    .A2(_04826_));
 sg13g2_o21ai_1 _23160_ (.B1(_06684_),
    .Y(_06685_),
    .A1(net689),
    .A2(_06682_));
 sg13g2_a221oi_1 _23161_ (.B2(\top_ihp.oisc.regs[63][6] ),
    .C1(_06685_),
    .B1(net571),
    .A1(\top_ihp.oisc.regs[2][6] ),
    .Y(_06686_),
    .A2(net440));
 sg13g2_a22oi_1 _23162_ (.Y(_06687_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[59][6] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[33][6] ));
 sg13g2_a22oi_1 _23163_ (.Y(_06688_),
    .B1(net446),
    .B2(\top_ihp.oisc.regs[60][6] ),
    .A2(net267),
    .A1(\top_ihp.oisc.regs[38][6] ));
 sg13g2_nand3_1 _23164_ (.B(_06687_),
    .C(_06688_),
    .A(_06686_),
    .Y(_06689_));
 sg13g2_nor4_1 _23165_ (.A(net78),
    .B(_06673_),
    .C(_06681_),
    .D(_06689_),
    .Y(_06690_));
 sg13g2_a21oi_1 _23166_ (.A1(_00113_),
    .A2(net78),
    .Y(_06691_),
    .B1(net154));
 sg13g2_nor2_1 _23167_ (.A(_06683_),
    .B(_06691_),
    .Y(_06692_));
 sg13g2_a21oi_1 _23168_ (.A1(_06667_),
    .A2(_06690_),
    .Y(_00322_),
    .B1(_06692_));
 sg13g2_a22oi_1 _23169_ (.Y(_06693_),
    .B1(net587),
    .B2(\top_ihp.oisc.regs[23][7] ),
    .A2(net608),
    .A1(\top_ihp.oisc.regs[1][7] ));
 sg13g2_a22oi_1 _23170_ (.Y(_06694_),
    .B1(net612),
    .B2(\top_ihp.oisc.regs[21][7] ),
    .A2(net477),
    .A1(\top_ihp.oisc.regs[14][7] ));
 sg13g2_mux2_1 _23171_ (.A0(\top_ihp.oisc.regs[10][7] ),
    .A1(\top_ihp.oisc.regs[8][7] ),
    .S(net656),
    .X(_06695_));
 sg13g2_nor2_1 _23172_ (.A(net669),
    .B(net679),
    .Y(_06696_));
 sg13g2_a22oi_1 _23173_ (.Y(_06697_),
    .B1(_06695_),
    .B2(_06696_),
    .A2(net647),
    .A1(\top_ihp.oisc.regs[11][7] ));
 sg13g2_a22oi_1 _23174_ (.Y(_06698_),
    .B1(net607),
    .B2(\top_ihp.oisc.regs[31][7] ),
    .A2(net613),
    .A1(\top_ihp.oisc.regs[29][7] ));
 sg13g2_nand4_1 _23175_ (.B(_06694_),
    .C(_06697_),
    .A(_06693_),
    .Y(_06699_),
    .D(_06698_));
 sg13g2_mux2_1 _23176_ (.A0(\top_ihp.oisc.regs[22][7] ),
    .A1(\top_ihp.oisc.regs[18][7] ),
    .S(net678),
    .X(_06700_));
 sg13g2_a22oi_1 _23177_ (.Y(_06701_),
    .B1(_04917_),
    .B2(_06700_),
    .A2(_05344_),
    .A1(\top_ihp.oisc.regs[25][7] ));
 sg13g2_mux2_1 _23178_ (.A0(\top_ihp.oisc.regs[53][7] ),
    .A1(\top_ihp.oisc.regs[52][7] ),
    .S(_04733_),
    .X(_06702_));
 sg13g2_nor4_1 _23179_ (.A(net678),
    .B(_04944_),
    .C(net643),
    .D(_04861_),
    .Y(_06703_));
 sg13g2_a22oi_1 _23180_ (.Y(_06704_),
    .B1(_06702_),
    .B2(_06703_),
    .A2(_04908_),
    .A1(\top_ihp.oisc.regs[5][7] ));
 sg13g2_mux2_1 _23181_ (.A0(\top_ihp.oisc.regs[3][7] ),
    .A1(\top_ihp.oisc.regs[19][7] ),
    .S(_04952_),
    .X(_06705_));
 sg13g2_a22oi_1 _23182_ (.Y(_06706_),
    .B1(net692),
    .B2(_06705_),
    .A2(net614),
    .A1(\top_ihp.oisc.regs[13][7] ));
 sg13g2_mux2_1 _23183_ (.A0(\top_ihp.oisc.regs[6][7] ),
    .A1(\top_ihp.oisc.regs[4][7] ),
    .S(net656),
    .X(_06707_));
 sg13g2_nor2_1 _23184_ (.A(_04772_),
    .B(_05388_),
    .Y(_06708_));
 sg13g2_a22oi_1 _23185_ (.Y(_06709_),
    .B1(_06707_),
    .B2(_06708_),
    .A2(_05393_),
    .A1(\top_ihp.oisc.regs[27][7] ));
 sg13g2_nand4_1 _23186_ (.B(_06704_),
    .C(_06706_),
    .A(_06701_),
    .Y(_06710_),
    .D(_06709_));
 sg13g2_mux2_1 _23187_ (.A0(\top_ihp.oisc.regs[24][7] ),
    .A1(\top_ihp.oisc.regs[16][7] ),
    .S(net667),
    .X(_06711_));
 sg13g2_a22oi_1 _23188_ (.Y(_06712_),
    .B1(_06711_),
    .B2(_04931_),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][7] ));
 sg13g2_nor2_1 _23189_ (.A(net689),
    .B(_06712_),
    .Y(_06713_));
 sg13g2_a22oi_1 _23190_ (.Y(_06714_),
    .B1(_05273_),
    .B2(\top_ihp.oisc.regs[12][7] ),
    .A2(_05007_),
    .A1(\top_ihp.oisc.regs[2][7] ));
 sg13g2_a22oi_1 _23191_ (.Y(_06715_),
    .B1(_05021_),
    .B2(\top_ihp.oisc.regs[9][7] ),
    .A2(net653),
    .A1(\top_ihp.oisc.regs[15][7] ));
 sg13g2_a22oi_1 _23192_ (.Y(_06716_),
    .B1(net657),
    .B2(\top_ihp.oisc.regs[7][7] ),
    .A2(_04820_),
    .A1(\top_ihp.oisc.regs[17][7] ));
 sg13g2_and2_1 _23193_ (.A(_06715_),
    .B(_06716_),
    .X(_06717_));
 sg13g2_o21ai_1 _23194_ (.B1(_06717_),
    .Y(_06718_),
    .A1(net688),
    .A2(_06714_));
 sg13g2_nor4_1 _23195_ (.A(_06699_),
    .B(_06710_),
    .C(_06713_),
    .D(_06718_),
    .Y(_06719_));
 sg13g2_nor2b_1 _23196_ (.A(net79),
    .B_N(_06719_),
    .Y(_06720_));
 sg13g2_a22oi_1 _23197_ (.Y(_06721_),
    .B1(_05307_),
    .B2(\top_ihp.oisc.regs[40][7] ),
    .A2(_05044_),
    .A1(\top_ihp.oisc.regs[44][7] ));
 sg13g2_a22oi_1 _23198_ (.Y(_06722_),
    .B1(_05115_),
    .B2(\top_ihp.oisc.regs[60][7] ),
    .A2(_04876_),
    .A1(\top_ihp.oisc.regs[33][7] ));
 sg13g2_a22oi_1 _23199_ (.Y(_06723_),
    .B1(_05192_),
    .B2(\top_ihp.oisc.regs[45][7] ),
    .A2(net462),
    .A1(\top_ihp.oisc.regs[36][7] ));
 sg13g2_a22oi_1 _23200_ (.Y(_06724_),
    .B1(_05164_),
    .B2(\top_ihp.oisc.regs[39][7] ),
    .A2(_05398_),
    .A1(\top_ihp.oisc.regs[48][7] ));
 sg13g2_nand4_1 _23201_ (.B(_06722_),
    .C(_06723_),
    .A(_06721_),
    .Y(_06725_),
    .D(_06724_));
 sg13g2_a22oi_1 _23202_ (.Y(_06726_),
    .B1(_05310_),
    .B2(\top_ihp.oisc.regs[46][7] ),
    .A2(_04979_),
    .A1(\top_ihp.oisc.regs[49][7] ));
 sg13g2_a22oi_1 _23203_ (.Y(_06727_),
    .B1(_05012_),
    .B2(\top_ihp.oisc.regs[51][7] ),
    .A2(_04984_),
    .A1(\top_ihp.oisc.regs[58][7] ));
 sg13g2_a22oi_1 _23204_ (.Y(_06728_),
    .B1(_05089_),
    .B2(\top_ihp.oisc.regs[37][7] ),
    .A2(_05036_),
    .A1(\top_ihp.oisc.regs[56][7] ));
 sg13g2_nand2_1 _23205_ (.Y(_06729_),
    .A(\top_ihp.oisc.regs[20][7] ),
    .B(_04855_));
 sg13g2_nand3_1 _23206_ (.B(net641),
    .C(net720),
    .A(\top_ihp.oisc.regs[26][7] ),
    .Y(_06730_));
 sg13g2_a22oi_1 _23207_ (.Y(_06731_),
    .B1(net646),
    .B2(\top_ihp.oisc.regs[30][7] ),
    .A2(net803),
    .A1(_07539_));
 sg13g2_nand3_1 _23208_ (.B(_06730_),
    .C(_06731_),
    .A(_06729_),
    .Y(_06732_));
 sg13g2_a21oi_1 _23209_ (.A1(\top_ihp.oisc.regs[43][7] ),
    .A2(net460),
    .Y(_06733_),
    .B1(_06732_));
 sg13g2_nand4_1 _23210_ (.B(_06727_),
    .C(_06728_),
    .A(_06726_),
    .Y(_06734_),
    .D(_06733_));
 sg13g2_a22oi_1 _23211_ (.Y(_06735_),
    .B1(_05383_),
    .B2(\top_ihp.oisc.regs[61][7] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[55][7] ));
 sg13g2_a22oi_1 _23212_ (.Y(_06736_),
    .B1(_05062_),
    .B2(\top_ihp.oisc.regs[57][7] ),
    .A2(net582),
    .A1(\top_ihp.oisc.regs[62][7] ));
 sg13g2_a22oi_1 _23213_ (.Y(_06737_),
    .B1(_05380_),
    .B2(\top_ihp.oisc.regs[42][7] ),
    .A2(net575),
    .A1(\top_ihp.oisc.regs[54][7] ));
 sg13g2_a22oi_1 _23214_ (.Y(_06738_),
    .B1(_05185_),
    .B2(\top_ihp.oisc.regs[50][7] ),
    .A2(_04966_),
    .A1(\top_ihp.oisc.regs[32][7] ));
 sg13g2_nand4_1 _23215_ (.B(_06736_),
    .C(_06737_),
    .A(_06735_),
    .Y(_06739_),
    .D(_06738_));
 sg13g2_a22oi_1 _23216_ (.Y(_06740_),
    .B1(net266),
    .B2(\top_ihp.oisc.regs[41][7] ),
    .A2(_05112_),
    .A1(\top_ihp.oisc.regs[35][7] ));
 sg13g2_a22oi_1 _23217_ (.Y(_06741_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[59][7] ),
    .A2(net265),
    .A1(\top_ihp.oisc.regs[47][7] ));
 sg13g2_nand2_1 _23218_ (.Y(_06742_),
    .A(\top_ihp.oisc.regs[38][7] ),
    .B(net267));
 sg13g2_a22oi_1 _23219_ (.Y(_06743_),
    .B1(_05334_),
    .B2(\top_ihp.oisc.regs[34][7] ),
    .A2(_05266_),
    .A1(\top_ihp.oisc.regs[63][7] ));
 sg13g2_nand4_1 _23220_ (.B(_06741_),
    .C(_06742_),
    .A(_06740_),
    .Y(_06744_),
    .D(_06743_));
 sg13g2_nor4_2 _23221_ (.A(_06725_),
    .B(_06734_),
    .C(_06739_),
    .Y(_06745_),
    .D(_06744_));
 sg13g2_a21oi_1 _23222_ (.A1(_00114_),
    .A2(net75),
    .Y(_06746_),
    .B1(net152));
 sg13g2_a21oi_1 _23223_ (.A1(_07539_),
    .A2(net685),
    .Y(_06747_),
    .B1(_06746_));
 sg13g2_a21oi_1 _23224_ (.A1(_06720_),
    .A2(_06745_),
    .Y(_00323_),
    .B1(_06747_));
 sg13g2_mux2_1 _23225_ (.A0(\top_ihp.oisc.regs[30][8] ),
    .A1(\top_ihp.oisc.regs[26][8] ),
    .S(net704),
    .X(_06748_));
 sg13g2_a22oi_1 _23226_ (.Y(_06749_),
    .B1(_06748_),
    .B2(net720),
    .A2(_04939_),
    .A1(\top_ihp.oisc.regs[31][8] ));
 sg13g2_a22oi_1 _23227_ (.Y(_06750_),
    .B1(_05015_),
    .B2(\top_ihp.oisc.regs[4][8] ),
    .A2(_04901_),
    .A1(\top_ihp.oisc.regs[21][8] ));
 sg13g2_a22oi_1 _23228_ (.Y(_06751_),
    .B1(net657),
    .B2(\top_ihp.oisc.regs[7][8] ),
    .A2(_04833_),
    .A1(\top_ihp.oisc.regs[24][8] ));
 sg13g2_a22oi_1 _23229_ (.Y(_06752_),
    .B1(_05254_),
    .B2(\top_ihp.oisc.regs[8][8] ),
    .A2(_04816_),
    .A1(\top_ihp.oisc.regs[25][8] ));
 sg13g2_nand4_1 _23230_ (.B(_06750_),
    .C(_06751_),
    .A(_06749_),
    .Y(_06753_),
    .D(_06752_));
 sg13g2_a22oi_1 _23231_ (.Y(_06754_),
    .B1(net561),
    .B2(\top_ihp.oisc.regs[27][8] ),
    .A2(net597),
    .A1(\top_ihp.oisc.regs[9][8] ));
 sg13g2_mux2_1 _23232_ (.A0(\top_ihp.oisc.regs[3][8] ),
    .A1(\top_ihp.oisc.regs[19][8] ),
    .S(net725),
    .X(_06755_));
 sg13g2_nand2_1 _23233_ (.Y(_06756_),
    .A(_04957_),
    .B(_06755_));
 sg13g2_nand2_1 _23234_ (.Y(_06757_),
    .A(_06754_),
    .B(_06756_));
 sg13g2_nor2_1 _23235_ (.A(_06753_),
    .B(_06757_),
    .Y(_06758_));
 sg13g2_a22oi_1 _23236_ (.Y(_06759_),
    .B1(net721),
    .B2(\top_ihp.oisc.regs[22][8] ),
    .A2(net722),
    .A1(\top_ihp.oisc.regs[20][8] ));
 sg13g2_nor2_1 _23237_ (.A(net672),
    .B(_06759_),
    .Y(_06760_));
 sg13g2_a21oi_1 _23238_ (.A1(_07580_),
    .A2(net772),
    .Y(_06761_),
    .B1(_06760_));
 sg13g2_a22oi_1 _23239_ (.Y(_06762_),
    .B1(net554),
    .B2(\top_ihp.oisc.regs[18][8] ),
    .A2(net645),
    .A1(\top_ihp.oisc.regs[16][8] ));
 sg13g2_a22oi_1 _23240_ (.Y(_06763_),
    .B1(net610),
    .B2(\top_ihp.oisc.regs[6][8] ),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][8] ));
 sg13g2_a22oi_1 _23241_ (.Y(_06764_),
    .B1(_05093_),
    .B2(\top_ihp.oisc.regs[41][8] ),
    .A2(_05061_),
    .A1(\top_ihp.oisc.regs[57][8] ));
 sg13g2_and4_1 _23242_ (.A(_06761_),
    .B(_06762_),
    .C(_06763_),
    .D(_06764_),
    .X(_06765_));
 sg13g2_a22oi_1 _23243_ (.Y(_06766_),
    .B1(net440),
    .B2(\top_ihp.oisc.regs[2][8] ),
    .A2(net463),
    .A1(\top_ihp.oisc.regs[32][8] ));
 sg13g2_a22oi_1 _23244_ (.Y(_06767_),
    .B1(_04765_),
    .B2(\top_ihp.oisc.regs[12][8] ),
    .A2(_04763_),
    .A1(\top_ihp.oisc.regs[10][8] ));
 sg13g2_nor2_1 _23245_ (.A(net679),
    .B(_06767_),
    .Y(_06768_));
 sg13g2_a21oi_1 _23246_ (.A1(\top_ihp.oisc.regs[37][8] ),
    .A2(net450),
    .Y(_06769_),
    .B1(_06768_));
 sg13g2_nand4_1 _23247_ (.B(_06765_),
    .C(_06766_),
    .A(_06758_),
    .Y(_06770_),
    .D(_06769_));
 sg13g2_a22oi_1 _23248_ (.Y(_06771_),
    .B1(_05112_),
    .B2(\top_ihp.oisc.regs[35][8] ),
    .A2(_04970_),
    .A1(\top_ihp.oisc.regs[54][8] ));
 sg13g2_a22oi_1 _23249_ (.Y(_06772_),
    .B1(_05334_),
    .B2(\top_ihp.oisc.regs[34][8] ),
    .A2(_05424_),
    .A1(\top_ihp.oisc.regs[51][8] ));
 sg13g2_a22oi_1 _23250_ (.Y(_06773_),
    .B1(_05377_),
    .B2(\top_ihp.oisc.regs[38][8] ),
    .A2(net475),
    .A1(\top_ihp.oisc.regs[55][8] ));
 sg13g2_a22oi_1 _23251_ (.Y(_06774_),
    .B1(_05299_),
    .B2(\top_ihp.oisc.regs[61][8] ),
    .A2(_05036_),
    .A1(\top_ihp.oisc.regs[56][8] ));
 sg13g2_nand4_1 _23252_ (.B(_06772_),
    .C(_06773_),
    .A(_06771_),
    .Y(_06775_),
    .D(_06774_));
 sg13g2_a22oi_1 _23253_ (.Y(_06776_),
    .B1(net472),
    .B2(\top_ihp.oisc.regs[29][8] ),
    .A2(net258),
    .A1(\top_ihp.oisc.regs[14][8] ));
 sg13g2_a22oi_1 _23254_ (.Y(_06777_),
    .B1(net558),
    .B2(\top_ihp.oisc.regs[11][8] ),
    .A2(net464),
    .A1(\top_ihp.oisc.regs[28][8] ));
 sg13g2_mux2_1 _23255_ (.A0(\top_ihp.oisc.regs[13][8] ),
    .A1(\top_ihp.oisc.regs[5][8] ),
    .S(net642),
    .X(_06778_));
 sg13g2_a22oi_1 _23256_ (.Y(_06779_),
    .B1(_06778_),
    .B2(_04905_),
    .A2(net467),
    .A1(\top_ihp.oisc.regs[15][8] ));
 sg13g2_a22oi_1 _23257_ (.Y(_06780_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[23][8] ),
    .A2(net608),
    .A1(\top_ihp.oisc.regs[1][8] ));
 sg13g2_nand4_1 _23258_ (.B(_06777_),
    .C(_06779_),
    .A(_06776_),
    .Y(_06781_),
    .D(_06780_));
 sg13g2_a22oi_1 _23259_ (.Y(_06782_),
    .B1(net414),
    .B2(\top_ihp.oisc.regs[59][8] ),
    .A2(_05177_),
    .A1(\top_ihp.oisc.regs[58][8] ));
 sg13g2_a22oi_1 _23260_ (.Y(_06783_),
    .B1(_05193_),
    .B2(\top_ihp.oisc.regs[45][8] ),
    .A2(net269),
    .A1(\top_ihp.oisc.regs[43][8] ));
 sg13g2_nand2_1 _23261_ (.Y(_06784_),
    .A(_06782_),
    .B(_06783_));
 sg13g2_nor4_1 _23262_ (.A(_06770_),
    .B(_06775_),
    .C(_06781_),
    .D(_06784_),
    .Y(_06785_));
 sg13g2_a22oi_1 _23263_ (.Y(_06786_),
    .B1(net268),
    .B2(\top_ihp.oisc.regs[44][8] ),
    .A2(_05191_),
    .A1(\top_ihp.oisc.regs[47][8] ));
 sg13g2_a22oi_1 _23264_ (.Y(_06787_),
    .B1(_05107_),
    .B2(\top_ihp.oisc.regs[46][8] ),
    .A2(_05266_),
    .A1(\top_ihp.oisc.regs[63][8] ));
 sg13g2_a22oi_1 _23265_ (.Y(_06788_),
    .B1(_05221_),
    .B2(\top_ihp.oisc.regs[39][8] ),
    .A2(_05302_),
    .A1(\top_ihp.oisc.regs[36][8] ));
 sg13g2_a22oi_1 _23266_ (.Y(_06789_),
    .B1(_05620_),
    .B2(\top_ihp.oisc.regs[62][8] ),
    .A2(_05380_),
    .A1(\top_ihp.oisc.regs[42][8] ));
 sg13g2_nand4_1 _23267_ (.B(_06787_),
    .C(_06788_),
    .A(_06786_),
    .Y(_06790_),
    .D(_06789_));
 sg13g2_a22oi_1 _23268_ (.Y(_06791_),
    .B1(net595),
    .B2(\top_ihp.oisc.regs[50][8] ),
    .A2(_05217_),
    .A1(\top_ihp.oisc.regs[33][8] ));
 sg13g2_a22oi_1 _23269_ (.Y(_06792_),
    .B1(_05116_),
    .B2(\top_ihp.oisc.regs[60][8] ),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[48][8] ));
 sg13g2_a22oi_1 _23270_ (.Y(_06793_),
    .B1(net417),
    .B2(\top_ihp.oisc.regs[49][8] ),
    .A2(_05173_),
    .A1(\top_ihp.oisc.regs[53][8] ));
 sg13g2_a22oi_1 _23271_ (.Y(_06794_),
    .B1(net263),
    .B2(\top_ihp.oisc.regs[40][8] ),
    .A2(_05068_),
    .A1(\top_ihp.oisc.regs[52][8] ));
 sg13g2_nand4_1 _23272_ (.B(_06792_),
    .C(_06793_),
    .A(_06791_),
    .Y(_06795_),
    .D(_06794_));
 sg13g2_nor3_1 _23273_ (.A(_05101_),
    .B(_06790_),
    .C(_06795_),
    .Y(_06796_));
 sg13g2_a21oi_1 _23274_ (.A1(_00115_),
    .A2(net75),
    .Y(_06797_),
    .B1(_05104_));
 sg13g2_a21oi_1 _23275_ (.A1(_07580_),
    .A2(net685),
    .Y(_06798_),
    .B1(_06797_));
 sg13g2_a21oi_1 _23276_ (.A1(_06785_),
    .A2(_06796_),
    .Y(_00324_),
    .B1(_06798_));
 sg13g2_a22oi_1 _23277_ (.Y(_06799_),
    .B1(net450),
    .B2(\top_ihp.oisc.regs[37][9] ),
    .A2(_04844_),
    .A1(\top_ihp.oisc.regs[47][9] ));
 sg13g2_a22oi_1 _23278_ (.Y(_06800_),
    .B1(net593),
    .B2(\top_ihp.oisc.regs[61][9] ),
    .A2(_04875_),
    .A1(\top_ihp.oisc.regs[33][9] ));
 sg13g2_a22oi_1 _23279_ (.Y(_06801_),
    .B1(_05071_),
    .B2(\top_ihp.oisc.regs[34][9] ),
    .A2(_04969_),
    .A1(\top_ihp.oisc.regs[54][9] ));
 sg13g2_a22oi_1 _23280_ (.Y(_06802_),
    .B1(_05067_),
    .B2(\top_ihp.oisc.regs[52][9] ),
    .A2(_04870_),
    .A1(\top_ihp.oisc.regs[55][9] ));
 sg13g2_nand4_1 _23281_ (.B(_06800_),
    .C(_06801_),
    .A(_06799_),
    .Y(_06803_),
    .D(_06802_));
 sg13g2_a22oi_1 _23282_ (.Y(_06804_),
    .B1(net569),
    .B2(\top_ihp.oisc.regs[9][9] ),
    .A2(net658),
    .A1(\top_ihp.oisc.regs[24][9] ));
 sg13g2_nand2_1 _23283_ (.Y(_06805_),
    .A(\top_ihp.oisc.regs[10][9] ),
    .B(net471));
 sg13g2_a22oi_1 _23284_ (.Y(_06806_),
    .B1(net610),
    .B2(\top_ihp.oisc.regs[6][9] ),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[5][9] ));
 sg13g2_a22oi_1 _23285_ (.Y(_06807_),
    .B1(net584),
    .B2(\top_ihp.oisc.regs[27][9] ),
    .A2(net619),
    .A1(\top_ihp.oisc.regs[25][9] ));
 sg13g2_nand4_1 _23286_ (.B(_06805_),
    .C(_06806_),
    .A(_06804_),
    .Y(_06808_),
    .D(_06807_));
 sg13g2_a22oi_1 _23287_ (.Y(_06809_),
    .B1(_05273_),
    .B2(\top_ihp.oisc.regs[12][9] ),
    .A2(_05007_),
    .A1(\top_ihp.oisc.regs[2][9] ));
 sg13g2_nor2_1 _23288_ (.A(net688),
    .B(_06809_),
    .Y(_06810_));
 sg13g2_mux2_1 _23289_ (.A0(\top_ihp.oisc.regs[20][9] ),
    .A1(\top_ihp.oisc.regs[16][9] ),
    .S(_05122_),
    .X(_06811_));
 sg13g2_a22oi_1 _23290_ (.Y(_06812_),
    .B1(_06811_),
    .B2(net640),
    .A2(net686),
    .A1(\top_ihp.oisc.regs[28][9] ));
 sg13g2_nor2_1 _23291_ (.A(_05280_),
    .B(_06812_),
    .Y(_06813_));
 sg13g2_nor4_1 _23292_ (.A(_06803_),
    .B(_06808_),
    .C(_06810_),
    .D(_06813_),
    .Y(_06814_));
 sg13g2_nor2b_1 _23293_ (.A(net79),
    .B_N(_06814_),
    .Y(_06815_));
 sg13g2_a22oi_1 _23294_ (.Y(_06816_),
    .B1(_05085_),
    .B2(\top_ihp.oisc.regs[40][9] ),
    .A2(_05058_),
    .A1(\top_ihp.oisc.regs[46][9] ));
 sg13g2_a22oi_1 _23295_ (.Y(_06817_),
    .B1(_05093_),
    .B2(\top_ihp.oisc.regs[41][9] ),
    .A2(_04988_),
    .A1(\top_ihp.oisc.regs[36][9] ));
 sg13g2_a22oi_1 _23296_ (.Y(_06818_),
    .B1(_05096_),
    .B2(\top_ihp.oisc.regs[60][9] ),
    .A2(_04974_),
    .A1(\top_ihp.oisc.regs[42][9] ));
 sg13g2_and2_1 _23297_ (.A(\top_ihp.oisc.regs[13][9] ),
    .B(net718),
    .X(_06819_));
 sg13g2_a21o_1 _23298_ (.A2(_05971_),
    .A1(\top_ihp.oisc.regs[1][9] ),
    .B1(_06819_),
    .X(_06820_));
 sg13g2_nor2_1 _23299_ (.A(net694),
    .B(net691),
    .Y(_06821_));
 sg13g2_a22oi_1 _23300_ (.Y(_06822_),
    .B1(_06820_),
    .B2(_06821_),
    .A2(_05043_),
    .A1(\top_ihp.oisc.regs[44][9] ));
 sg13g2_nand4_1 _23301_ (.B(_06817_),
    .C(_06818_),
    .A(_06816_),
    .Y(_06823_),
    .D(_06822_));
 sg13g2_nand2_1 _23302_ (.Y(_06824_),
    .A(\top_ihp.oisc.regs[29][9] ),
    .B(net613));
 sg13g2_a22oi_1 _23303_ (.Y(_06825_),
    .B1(_05245_),
    .B2(\top_ihp.oisc.regs[3][9] ),
    .A2(_03690_),
    .A1(_07547_));
 sg13g2_a22oi_1 _23304_ (.Y(_06826_),
    .B1(_05254_),
    .B2(\top_ihp.oisc.regs[8][9] ),
    .A2(_04826_),
    .A1(\top_ihp.oisc.regs[14][9] ));
 sg13g2_nand3_1 _23305_ (.B(_06825_),
    .C(_06826_),
    .A(_06824_),
    .Y(_06827_));
 sg13g2_nand2_1 _23306_ (.Y(_06828_),
    .A(\top_ihp.oisc.regs[58][9] ),
    .B(_04983_));
 sg13g2_nand2_1 _23307_ (.Y(_06829_),
    .A(\top_ihp.oisc.regs[26][9] ),
    .B(_05238_));
 sg13g2_a22oi_1 _23308_ (.Y(_06830_),
    .B1(_05241_),
    .B2(\top_ihp.oisc.regs[19][9] ),
    .A2(net646),
    .A1(\top_ihp.oisc.regs[30][9] ));
 sg13g2_nand3_1 _23309_ (.B(_06829_),
    .C(_06830_),
    .A(_06828_),
    .Y(_06831_));
 sg13g2_a22oi_1 _23310_ (.Y(_06832_),
    .B1(net651),
    .B2(\top_ihp.oisc.regs[11][9] ),
    .A2(net583),
    .A1(\top_ihp.oisc.regs[21][9] ));
 sg13g2_a22oi_1 _23311_ (.Y(_06833_),
    .B1(net577),
    .B2(\top_ihp.oisc.regs[4][9] ),
    .A2(net586),
    .A1(\top_ihp.oisc.regs[17][9] ));
 sg13g2_mux2_1 _23312_ (.A0(\top_ihp.oisc.regs[22][9] ),
    .A1(\top_ihp.oisc.regs[18][9] ),
    .S(_05326_),
    .X(_06834_));
 sg13g2_a22oi_1 _23313_ (.Y(_06835_),
    .B1(_06834_),
    .B2(net695),
    .A2(_05141_),
    .A1(\top_ihp.oisc.regs[23][9] ));
 sg13g2_mux2_1 _23314_ (.A0(\top_ihp.oisc.regs[15][9] ),
    .A1(\top_ihp.oisc.regs[7][9] ),
    .S(net670),
    .X(_06836_));
 sg13g2_a22oi_1 _23315_ (.Y(_06837_),
    .B1(_06184_),
    .B2(_06836_),
    .A2(net573),
    .A1(\top_ihp.oisc.regs[31][9] ));
 sg13g2_nand4_1 _23316_ (.B(_06833_),
    .C(_06835_),
    .A(_06832_),
    .Y(_06838_),
    .D(_06837_));
 sg13g2_or4_1 _23317_ (.A(_06823_),
    .B(_06827_),
    .C(_06831_),
    .D(_06838_),
    .X(_06839_));
 sg13g2_a22oi_1 _23318_ (.Y(_06840_),
    .B1(_05481_),
    .B2(\top_ihp.oisc.regs[35][9] ),
    .A2(_05174_),
    .A1(\top_ihp.oisc.regs[51][9] ));
 sg13g2_a22oi_1 _23319_ (.Y(_06841_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[63][9] ),
    .A2(net417),
    .A1(\top_ihp.oisc.regs[49][9] ));
 sg13g2_a22oi_1 _23320_ (.Y(_06842_),
    .B1(_05040_),
    .B2(\top_ihp.oisc.regs[50][9] ),
    .A2(_05226_),
    .A1(\top_ihp.oisc.regs[32][9] ));
 sg13g2_a22oi_1 _23321_ (.Y(_06843_),
    .B1(net553),
    .B2(\top_ihp.oisc.regs[62][9] ),
    .A2(_05377_),
    .A1(\top_ihp.oisc.regs[38][9] ));
 sg13g2_nand4_1 _23322_ (.B(_06841_),
    .C(_06842_),
    .A(_06840_),
    .Y(_06844_),
    .D(_06843_));
 sg13g2_a22oi_1 _23323_ (.Y(_06845_),
    .B1(net269),
    .B2(\top_ihp.oisc.regs[43][9] ),
    .A2(net414),
    .A1(\top_ihp.oisc.regs[59][9] ));
 sg13g2_a22oi_1 _23324_ (.Y(_06846_),
    .B1(_05193_),
    .B2(\top_ihp.oisc.regs[45][9] ),
    .A2(net413),
    .A1(\top_ihp.oisc.regs[57][9] ));
 sg13g2_a22oi_1 _23325_ (.Y(_06847_),
    .B1(_05221_),
    .B2(\top_ihp.oisc.regs[39][9] ),
    .A2(_05173_),
    .A1(\top_ihp.oisc.regs[53][9] ));
 sg13g2_a22oi_1 _23326_ (.Y(_06848_),
    .B1(_05758_),
    .B2(\top_ihp.oisc.regs[56][9] ),
    .A2(_05183_),
    .A1(\top_ihp.oisc.regs[48][9] ));
 sg13g2_nand4_1 _23327_ (.B(_06846_),
    .C(_06847_),
    .A(_06845_),
    .Y(_06849_),
    .D(_06848_));
 sg13g2_nor3_1 _23328_ (.A(_06839_),
    .B(_06844_),
    .C(_06849_),
    .Y(_06850_));
 sg13g2_a21oi_1 _23329_ (.A1(_00116_),
    .A2(_04810_),
    .Y(_06851_),
    .B1(_05104_));
 sg13g2_a21oi_1 _23330_ (.A1(_07547_),
    .A2(net685),
    .Y(_06852_),
    .B1(_06851_));
 sg13g2_a21oi_1 _23331_ (.A1(_06815_),
    .A2(_06850_),
    .Y(_00325_),
    .B1(_06852_));
 sg13g2_buf_1 _23332_ (.A(net735),
    .X(_06853_));
 sg13g2_nor2_1 _23333_ (.A(net879),
    .B(net939),
    .Y(_06854_));
 sg13g2_buf_1 _23334_ (.A(_06854_),
    .X(_06855_));
 sg13g2_buf_1 _23335_ (.A(net828),
    .X(_06856_));
 sg13g2_buf_1 _23336_ (.A(net812),
    .X(_06857_));
 sg13g2_or2_1 _23337_ (.X(_06858_),
    .B(_08233_),
    .A(_08227_));
 sg13g2_buf_1 _23338_ (.A(_06858_),
    .X(_06859_));
 sg13g2_nor3_1 _23339_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_06859_),
    .Y(_06860_));
 sg13g2_buf_1 _23340_ (.A(_06860_),
    .X(_06861_));
 sg13g2_or2_1 _23341_ (.X(_06862_),
    .B(_08231_),
    .A(_08232_));
 sg13g2_buf_1 _23342_ (.A(_06862_),
    .X(_06863_));
 sg13g2_nor3_1 _23343_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_06863_),
    .Y(_06864_));
 sg13g2_buf_1 _23344_ (.A(_06864_),
    .X(_06865_));
 sg13g2_buf_1 _23345_ (.A(_06865_),
    .X(_06866_));
 sg13g2_a22oi_1 _23346_ (.Y(_06867_),
    .B1(_06866_),
    .B2(\top_ihp.oisc.regs[2][0] ),
    .A2(_06861_),
    .A1(\top_ihp.oisc.regs[1][0] ));
 sg13g2_nand2_2 _23347_ (.Y(_06868_),
    .A(_08227_),
    .B(\top_ihp.oisc.reg_rb[0] ));
 sg13g2_nor3_1 _23348_ (.A(\top_ihp.oisc.reg_rb[3] ),
    .B(\top_ihp.oisc.reg_rb[2] ),
    .C(_06868_),
    .Y(_06869_));
 sg13g2_buf_1 _23349_ (.A(_06869_),
    .X(_06870_));
 sg13g2_nand2_1 _23350_ (.Y(_06871_),
    .A(\top_ihp.oisc.regs[3][0] ),
    .B(_06870_));
 sg13g2_nand2_1 _23351_ (.Y(_06872_),
    .A(_08238_),
    .B(\top_ihp.oisc.reg_rb[3] ));
 sg13g2_nor2_1 _23352_ (.A(_06859_),
    .B(_06872_),
    .Y(_06873_));
 sg13g2_buf_2 _23353_ (.A(_06873_),
    .X(_06874_));
 sg13g2_buf_1 _23354_ (.A(_06874_),
    .X(_06875_));
 sg13g2_nor3_1 _23355_ (.A(_08238_),
    .B(_08235_),
    .C(_06863_),
    .Y(_06876_));
 sg13g2_buf_1 _23356_ (.A(_06876_),
    .X(_06877_));
 sg13g2_buf_1 _23357_ (.A(_06877_),
    .X(_06878_));
 sg13g2_a22oi_1 _23358_ (.Y(_06879_),
    .B1(net794),
    .B2(\top_ihp.oisc.regs[10][0] ),
    .A2(_06875_),
    .A1(\top_ihp.oisc.regs[13][0] ));
 sg13g2_nand2_1 _23359_ (.Y(_06880_),
    .A(_08231_),
    .B(_08233_));
 sg13g2_nor2_1 _23360_ (.A(_06872_),
    .B(_06880_),
    .Y(_06881_));
 sg13g2_buf_1 _23361_ (.A(_06881_),
    .X(_06882_));
 sg13g2_buf_2 _23362_ (.A(_06882_),
    .X(_06883_));
 sg13g2_nor2_1 _23363_ (.A(_06863_),
    .B(_06872_),
    .Y(_06884_));
 sg13g2_buf_1 _23364_ (.A(_06884_),
    .X(_06885_));
 sg13g2_buf_2 _23365_ (.A(_06885_),
    .X(_06886_));
 sg13g2_a22oi_1 _23366_ (.Y(_06887_),
    .B1(_06886_),
    .B2(\top_ihp.oisc.regs[14][0] ),
    .A2(net761),
    .A1(\top_ihp.oisc.regs[12][0] ));
 sg13g2_nand4_1 _23367_ (.B(_06871_),
    .C(_06879_),
    .A(_06867_),
    .Y(_06888_),
    .D(_06887_));
 sg13g2_nor2_1 _23368_ (.A(_06868_),
    .B(_06872_),
    .Y(_06889_));
 sg13g2_buf_2 _23369_ (.A(_06889_),
    .X(_06890_));
 sg13g2_buf_1 _23370_ (.A(_06890_),
    .X(_06891_));
 sg13g2_nor3_1 _23371_ (.A(_08238_),
    .B(_08235_),
    .C(_06868_),
    .Y(_06892_));
 sg13g2_buf_1 _23372_ (.A(_06892_),
    .X(_06893_));
 sg13g2_buf_1 _23373_ (.A(_06893_),
    .X(_06894_));
 sg13g2_a22oi_1 _23374_ (.Y(_06895_),
    .B1(net793),
    .B2(\top_ihp.oisc.regs[11][0] ),
    .A2(net759),
    .A1(\top_ihp.oisc.regs[15][0] ));
 sg13g2_nor3_1 _23375_ (.A(_08238_),
    .B(_08235_),
    .C(_06880_),
    .Y(_06896_));
 sg13g2_buf_1 _23376_ (.A(_06896_),
    .X(_06897_));
 sg13g2_buf_1 _23377_ (.A(_06897_),
    .X(_06898_));
 sg13g2_a22oi_1 _23378_ (.Y(_06899_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[8][0] ),
    .A2(_06856_),
    .A1(\top_ihp.oisc.regs[32][0] ));
 sg13g2_nor3_1 _23379_ (.A(_08238_),
    .B(_08235_),
    .C(_06859_),
    .Y(_06900_));
 sg13g2_buf_2 _23380_ (.A(_06900_),
    .X(_06901_));
 sg13g2_buf_1 _23381_ (.A(_06901_),
    .X(_06902_));
 sg13g2_nor4_1 _23382_ (.A(_08238_),
    .B(\top_ihp.oisc.micro_op[11] ),
    .C(_08232_),
    .D(_08227_),
    .Y(_06903_));
 sg13g2_and2_1 _23383_ (.A(net939),
    .B(_06903_),
    .X(_06904_));
 sg13g2_buf_1 _23384_ (.A(_06904_),
    .X(_06905_));
 sg13g2_buf_1 _23385_ (.A(net865),
    .X(_06906_));
 sg13g2_a21oi_1 _23386_ (.A1(\top_ihp.oisc.regs[9][0] ),
    .A2(_06902_),
    .Y(_06907_),
    .B1(net848));
 sg13g2_nand3_1 _23387_ (.B(_06899_),
    .C(_06907_),
    .A(_06895_),
    .Y(_06908_));
 sg13g2_nand2_1 _23388_ (.Y(_06909_),
    .A(_08235_),
    .B(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_nor2_1 _23389_ (.A(_06880_),
    .B(_06909_),
    .Y(_06910_));
 sg13g2_buf_1 _23390_ (.A(_06910_),
    .X(_06911_));
 sg13g2_nor2_1 _23391_ (.A(_06868_),
    .B(_06909_),
    .Y(_06912_));
 sg13g2_buf_1 _23392_ (.A(_06912_),
    .X(_06913_));
 sg13g2_a22oi_1 _23393_ (.Y(_06914_),
    .B1(_06913_),
    .B2(\top_ihp.oisc.regs[7][0] ),
    .A2(_06911_),
    .A1(\top_ihp.oisc.regs[4][0] ));
 sg13g2_nor2_1 _23394_ (.A(_06863_),
    .B(_06909_),
    .Y(_06915_));
 sg13g2_buf_1 _23395_ (.A(_06915_),
    .X(_06916_));
 sg13g2_nor2_1 _23396_ (.A(_06859_),
    .B(_06909_),
    .Y(_06917_));
 sg13g2_buf_1 _23397_ (.A(_06917_),
    .X(_06918_));
 sg13g2_a22oi_1 _23398_ (.Y(_06919_),
    .B1(_06918_),
    .B2(\top_ihp.oisc.regs[5][0] ),
    .A2(_06916_),
    .A1(\top_ihp.oisc.regs[6][0] ));
 sg13g2_nand2_1 _23399_ (.Y(_06920_),
    .A(_06914_),
    .B(_06919_));
 sg13g2_nor3_1 _23400_ (.A(_06888_),
    .B(_06908_),
    .C(_06920_),
    .Y(_06921_));
 sg13g2_nand2_1 _23401_ (.Y(_06922_),
    .A(net939),
    .B(_06903_));
 sg13g2_buf_1 _23402_ (.A(_06922_),
    .X(_06923_));
 sg13g2_buf_1 _23403_ (.A(_06923_),
    .X(_06924_));
 sg13g2_nor2_1 _23404_ (.A(\top_ihp.oisc.regs[0][0] ),
    .B(_06924_),
    .Y(_06925_));
 sg13g2_nor4_1 _23405_ (.A(net735),
    .B(net796),
    .C(_06921_),
    .D(_06925_),
    .Y(_06926_));
 sg13g2_a21o_1 _23406_ (.A2(net684),
    .A1(_07474_),
    .B1(_06926_),
    .X(_00326_));
 sg13g2_buf_1 _23407_ (.A(net773),
    .X(_06927_));
 sg13g2_buf_1 _23408_ (.A(_06916_),
    .X(_06928_));
 sg13g2_buf_1 _23409_ (.A(_06918_),
    .X(_06929_));
 sg13g2_a22oi_1 _23410_ (.Y(_06930_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][10] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][10] ));
 sg13g2_buf_1 _23411_ (.A(_06861_),
    .X(_06931_));
 sg13g2_buf_1 _23412_ (.A(_06911_),
    .X(_06932_));
 sg13g2_a22oi_1 _23413_ (.Y(_06933_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][10] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][10] ));
 sg13g2_nand2_1 _23414_ (.Y(_06934_),
    .A(_06930_),
    .B(_06933_));
 sg13g2_buf_1 _23415_ (.A(_06897_),
    .X(_06935_));
 sg13g2_buf_1 _23416_ (.A(net810),
    .X(_06936_));
 sg13g2_nand2_1 _23417_ (.Y(_06937_),
    .A(\top_ihp.oisc.regs[8][10] ),
    .B(net790));
 sg13g2_buf_1 _23418_ (.A(_06891_),
    .X(_06938_));
 sg13g2_buf_1 _23419_ (.A(net792),
    .X(_06939_));
 sg13g2_a22oi_1 _23420_ (.Y(_06940_),
    .B1(net755),
    .B2(\top_ihp.oisc.regs[9][10] ),
    .A2(net716),
    .A1(\top_ihp.oisc.regs[15][10] ));
 sg13g2_buf_1 _23421_ (.A(_06870_),
    .X(_06941_));
 sg13g2_buf_1 _23422_ (.A(_06913_),
    .X(_06942_));
 sg13g2_a22oi_1 _23423_ (.Y(_06943_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[7][10] ),
    .A2(net789),
    .A1(\top_ihp.oisc.regs[3][10] ));
 sg13g2_buf_1 _23424_ (.A(net795),
    .X(_06944_));
 sg13g2_buf_2 _23425_ (.A(_06885_),
    .X(_06945_));
 sg13g2_a22oi_1 _23426_ (.Y(_06946_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[32][10] ),
    .A2(net752),
    .A1(\top_ihp.oisc.regs[14][10] ));
 sg13g2_buf_1 _23427_ (.A(_06877_),
    .X(_06947_));
 sg13g2_buf_1 _23428_ (.A(_06893_),
    .X(_06948_));
 sg13g2_a22oi_1 _23429_ (.Y(_06949_),
    .B1(net787),
    .B2(\top_ihp.oisc.regs[11][10] ),
    .A2(net788),
    .A1(\top_ihp.oisc.regs[10][10] ));
 sg13g2_buf_1 _23430_ (.A(_06874_),
    .X(_06950_));
 sg13g2_buf_2 _23431_ (.A(_06882_),
    .X(_06951_));
 sg13g2_a22oi_1 _23432_ (.Y(_06952_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][10] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][10] ));
 sg13g2_nand4_1 _23433_ (.B(_06946_),
    .C(_06949_),
    .A(net847),
    .Y(_06953_),
    .D(_06952_));
 sg13g2_a21oi_1 _23434_ (.A1(\top_ihp.oisc.regs[2][10] ),
    .A2(net753),
    .Y(_06954_),
    .B1(_06953_));
 sg13g2_nand4_1 _23435_ (.B(_06940_),
    .C(_06943_),
    .A(_06937_),
    .Y(_06955_),
    .D(_06954_));
 sg13g2_buf_1 _23436_ (.A(net848),
    .X(_06956_));
 sg13g2_buf_1 _23437_ (.A(net812),
    .X(_06957_));
 sg13g2_a21oi_1 _23438_ (.A1(_00117_),
    .A2(net827),
    .Y(_06958_),
    .B1(net786));
 sg13g2_o21ai_1 _23439_ (.B1(_06958_),
    .Y(_06959_),
    .A1(_06934_),
    .A2(_06955_));
 sg13g2_buf_1 _23440_ (.A(net773),
    .X(_06960_));
 sg13g2_nor2_1 _23441_ (.A(_07535_),
    .B(net715),
    .Y(_06961_));
 sg13g2_a21oi_1 _23442_ (.A1(net717),
    .A2(_06959_),
    .Y(_00327_),
    .B1(_06961_));
 sg13g2_buf_1 _23443_ (.A(_06870_),
    .X(_06962_));
 sg13g2_a22oi_1 _23444_ (.Y(_06963_),
    .B1(net785),
    .B2(\top_ihp.oisc.regs[3][11] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][11] ));
 sg13g2_nand2_1 _23445_ (.Y(_06964_),
    .A(\top_ihp.oisc.regs[12][11] ),
    .B(net761));
 sg13g2_a22oi_1 _23446_ (.Y(_06965_),
    .B1(net793),
    .B2(\top_ihp.oisc.regs[11][11] ),
    .A2(net759),
    .A1(\top_ihp.oisc.regs[15][11] ));
 sg13g2_buf_1 _23447_ (.A(net795),
    .X(_06966_));
 sg13g2_buf_1 _23448_ (.A(_06885_),
    .X(_06967_));
 sg13g2_buf_1 _23449_ (.A(net828),
    .X(_06968_));
 sg13g2_a22oi_1 _23450_ (.Y(_06969_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][11] ),
    .A2(net748),
    .A1(\top_ihp.oisc.regs[14][11] ));
 sg13g2_a22oi_1 _23451_ (.Y(_06970_),
    .B1(_06901_),
    .B2(\top_ihp.oisc.regs[9][11] ),
    .A2(_06897_),
    .A1(\top_ihp.oisc.regs[8][11] ));
 sg13g2_a22oi_1 _23452_ (.Y(_06971_),
    .B1(net788),
    .B2(\top_ihp.oisc.regs[10][11] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][11] ));
 sg13g2_nand4_1 _23453_ (.B(_06969_),
    .C(_06970_),
    .A(net864),
    .Y(_06972_),
    .D(_06971_));
 sg13g2_a21oi_1 _23454_ (.A1(\top_ihp.oisc.regs[2][11] ),
    .A2(net749),
    .Y(_06973_),
    .B1(_06972_));
 sg13g2_nand4_1 _23455_ (.B(_06964_),
    .C(_06965_),
    .A(_06963_),
    .Y(_06974_),
    .D(_06973_));
 sg13g2_buf_1 _23456_ (.A(_06911_),
    .X(_06975_));
 sg13g2_buf_1 _23457_ (.A(_06918_),
    .X(_06976_));
 sg13g2_a22oi_1 _23458_ (.Y(_06977_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][11] ),
    .A2(net747),
    .A1(\top_ihp.oisc.regs[4][11] ));
 sg13g2_buf_1 _23459_ (.A(_06916_),
    .X(_06978_));
 sg13g2_a22oi_1 _23460_ (.Y(_06979_),
    .B1(net745),
    .B2(\top_ihp.oisc.regs[6][11] ),
    .A2(net754),
    .A1(\top_ihp.oisc.regs[7][11] ));
 sg13g2_nand2_1 _23461_ (.Y(_06980_),
    .A(_06977_),
    .B(_06979_));
 sg13g2_a21oi_1 _23462_ (.A1(_00118_),
    .A2(net827),
    .Y(_06981_),
    .B1(net786));
 sg13g2_o21ai_1 _23463_ (.B1(_06981_),
    .Y(_06982_),
    .A1(_06974_),
    .A2(_06980_));
 sg13g2_nor2_1 _23464_ (.A(_07532_),
    .B(net715),
    .Y(_06983_));
 sg13g2_a21oi_1 _23465_ (.A1(net717),
    .A2(_06982_),
    .Y(_00328_),
    .B1(_06983_));
 sg13g2_buf_1 _23466_ (.A(_06911_),
    .X(_06984_));
 sg13g2_buf_1 _23467_ (.A(_06913_),
    .X(_06985_));
 sg13g2_a22oi_1 _23468_ (.Y(_06986_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][12] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][12] ));
 sg13g2_buf_1 _23469_ (.A(_06916_),
    .X(_06987_));
 sg13g2_buf_1 _23470_ (.A(_06918_),
    .X(_06988_));
 sg13g2_a22oi_1 _23471_ (.Y(_06989_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][12] ),
    .A2(net742),
    .A1(\top_ihp.oisc.regs[6][12] ));
 sg13g2_nand2_1 _23472_ (.Y(_06990_),
    .A(_06986_),
    .B(_06989_));
 sg13g2_nand2_1 _23473_ (.Y(_06991_),
    .A(\top_ihp.oisc.regs[8][12] ),
    .B(net790));
 sg13g2_a22oi_1 _23474_ (.Y(_06992_),
    .B1(net761),
    .B2(\top_ihp.oisc.regs[12][12] ),
    .A2(net794),
    .A1(\top_ihp.oisc.regs[10][12] ));
 sg13g2_buf_1 _23475_ (.A(_06861_),
    .X(_06993_));
 sg13g2_a22oi_1 _23476_ (.Y(_06994_),
    .B1(net785),
    .B2(\top_ihp.oisc.regs[3][12] ),
    .A2(net784),
    .A1(\top_ihp.oisc.regs[1][12] ));
 sg13g2_buf_1 _23477_ (.A(_06893_),
    .X(_06995_));
 sg13g2_a22oi_1 _23478_ (.Y(_06996_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[32][12] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][12] ));
 sg13g2_a22oi_1 _23479_ (.Y(_06997_),
    .B1(net759),
    .B2(\top_ihp.oisc.regs[15][12] ),
    .A2(net748),
    .A1(\top_ihp.oisc.regs[14][12] ));
 sg13g2_buf_1 _23480_ (.A(_06901_),
    .X(_06998_));
 sg13g2_a22oi_1 _23481_ (.Y(_06999_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][12] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][12] ));
 sg13g2_nand4_1 _23482_ (.B(_06996_),
    .C(_06997_),
    .A(net847),
    .Y(_07000_),
    .D(_06999_));
 sg13g2_a21oi_1 _23483_ (.A1(\top_ihp.oisc.regs[2][12] ),
    .A2(net753),
    .Y(_07001_),
    .B1(_07000_));
 sg13g2_nand4_1 _23484_ (.B(_06992_),
    .C(_06994_),
    .A(_06991_),
    .Y(_07002_),
    .D(_07001_));
 sg13g2_a21oi_1 _23485_ (.A1(_00119_),
    .A2(net827),
    .Y(_07003_),
    .B1(net786));
 sg13g2_o21ai_1 _23486_ (.B1(_07003_),
    .Y(_07004_),
    .A1(_06990_),
    .A2(_07002_));
 sg13g2_buf_1 _23487_ (.A(net773),
    .X(_07005_));
 sg13g2_nor2_1 _23488_ (.A(_07529_),
    .B(net714),
    .Y(_07006_));
 sg13g2_a21oi_1 _23489_ (.A1(net717),
    .A2(_07004_),
    .Y(_00329_),
    .B1(_07006_));
 sg13g2_a22oi_1 _23490_ (.Y(_07007_),
    .B1(_06929_),
    .B2(\top_ihp.oisc.regs[5][13] ),
    .A2(_06928_),
    .A1(\top_ihp.oisc.regs[6][13] ));
 sg13g2_a22oi_1 _23491_ (.Y(_07008_),
    .B1(net747),
    .B2(\top_ihp.oisc.regs[4][13] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][13] ));
 sg13g2_nand2_1 _23492_ (.Y(_07009_),
    .A(_07007_),
    .B(_07008_));
 sg13g2_nand2_1 _23493_ (.Y(_07010_),
    .A(\top_ihp.oisc.regs[14][13] ),
    .B(_06886_));
 sg13g2_buf_2 _23494_ (.A(net759),
    .X(_07011_));
 sg13g2_a22oi_1 _23495_ (.Y(_07012_),
    .B1(net713),
    .B2(\top_ihp.oisc.regs[15][13] ),
    .A2(net794),
    .A1(\top_ihp.oisc.regs[10][13] ));
 sg13g2_a22oi_1 _23496_ (.Y(_07013_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[7][13] ),
    .A2(net789),
    .A1(\top_ihp.oisc.regs[3][13] ));
 sg13g2_a22oi_1 _23497_ (.Y(_07014_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][13] ),
    .A2(net809),
    .A1(\top_ihp.oisc.regs[32][13] ));
 sg13g2_a22oi_1 _23498_ (.Y(_07015_),
    .B1(_06898_),
    .B2(\top_ihp.oisc.regs[8][13] ),
    .A2(_06950_),
    .A1(\top_ihp.oisc.regs[13][13] ));
 sg13g2_buf_1 _23499_ (.A(_06882_),
    .X(_07016_));
 sg13g2_a22oi_1 _23500_ (.Y(_07017_),
    .B1(net787),
    .B2(\top_ihp.oisc.regs[11][13] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][13] ));
 sg13g2_nand4_1 _23501_ (.B(_07014_),
    .C(_07015_),
    .A(net847),
    .Y(_07018_),
    .D(_07017_));
 sg13g2_a21oi_1 _23502_ (.A1(\top_ihp.oisc.regs[2][13] ),
    .A2(net753),
    .Y(_07019_),
    .B1(_07018_));
 sg13g2_nand4_1 _23503_ (.B(_07012_),
    .C(_07013_),
    .A(_07010_),
    .Y(_07020_),
    .D(_07019_));
 sg13g2_a21oi_1 _23504_ (.A1(_00120_),
    .A2(net827),
    .Y(_07021_),
    .B1(_06957_));
 sg13g2_o21ai_1 _23505_ (.B1(_07021_),
    .Y(_07022_),
    .A1(_07009_),
    .A2(_07020_));
 sg13g2_nor2_1 _23506_ (.A(_07526_),
    .B(net714),
    .Y(_07023_));
 sg13g2_a21oi_1 _23507_ (.A1(net717),
    .A2(_07022_),
    .Y(_00330_),
    .B1(_07023_));
 sg13g2_buf_1 _23508_ (.A(net735),
    .X(_07024_));
 sg13g2_a22oi_1 _23509_ (.Y(_07025_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][14] ),
    .A2(net747),
    .A1(\top_ihp.oisc.regs[4][14] ));
 sg13g2_a22oi_1 _23510_ (.Y(_07026_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][14] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][14] ));
 sg13g2_buf_1 _23511_ (.A(net762),
    .X(_07027_));
 sg13g2_and2_1 _23512_ (.A(\top_ihp.oisc.regs[9][14] ),
    .B(net792),
    .X(_07028_));
 sg13g2_a221oi_1 _23513_ (.B2(\top_ihp.oisc.regs[10][14] ),
    .C1(_07028_),
    .B1(net794),
    .A1(\top_ihp.oisc.regs[13][14] ),
    .Y(_07029_),
    .A2(net712));
 sg13g2_nand2_1 _23514_ (.Y(_07030_),
    .A(\top_ihp.oisc.regs[2][14] ),
    .B(net795));
 sg13g2_buf_1 _23515_ (.A(_06855_),
    .X(_07031_));
 sg13g2_a221oi_1 _23516_ (.B2(\top_ihp.oisc.regs[32][14] ),
    .C1(net848),
    .B1(net808),
    .A1(\top_ihp.oisc.regs[11][14] ),
    .Y(_07032_),
    .A2(net783));
 sg13g2_a22oi_1 _23517_ (.Y(_07033_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[8][14] ),
    .A2(net759),
    .A1(\top_ihp.oisc.regs[15][14] ));
 sg13g2_a22oi_1 _23518_ (.Y(_07034_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[14][14] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][14] ));
 sg13g2_nand4_1 _23519_ (.B(_07032_),
    .C(_07033_),
    .A(_07030_),
    .Y(_07035_),
    .D(_07034_));
 sg13g2_a221oi_1 _23520_ (.B2(\top_ihp.oisc.regs[3][14] ),
    .C1(_07035_),
    .B1(net789),
    .A1(\top_ihp.oisc.regs[1][14] ),
    .Y(_07036_),
    .A2(_06861_));
 sg13g2_nand4_1 _23521_ (.B(_07026_),
    .C(_07029_),
    .A(_07025_),
    .Y(_07037_),
    .D(_07036_));
 sg13g2_buf_1 _23522_ (.A(net848),
    .X(_07038_));
 sg13g2_a21oi_1 _23523_ (.A1(_00121_),
    .A2(net826),
    .Y(_07039_),
    .B1(net796));
 sg13g2_a21oi_1 _23524_ (.A1(_07037_),
    .A2(_07039_),
    .Y(_07040_),
    .B1(net684));
 sg13g2_a21oi_1 _23525_ (.A1(_07898_),
    .A2(net683),
    .Y(_00331_),
    .B1(_07040_));
 sg13g2_a22oi_1 _23526_ (.Y(_07041_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][15] ),
    .A2(net745),
    .A1(\top_ihp.oisc.regs[6][15] ));
 sg13g2_buf_1 _23527_ (.A(_06861_),
    .X(_07042_));
 sg13g2_a22oi_1 _23528_ (.Y(_07043_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][15] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][15] ));
 sg13g2_and2_1 _23529_ (.A(\top_ihp.oisc.regs[8][15] ),
    .B(net790),
    .X(_07044_));
 sg13g2_a221oi_1 _23530_ (.B2(\top_ihp.oisc.regs[12][15] ),
    .C1(_07044_),
    .B1(net761),
    .A1(\top_ihp.oisc.regs[13][15] ),
    .Y(_07045_),
    .A2(net712));
 sg13g2_buf_1 _23531_ (.A(_06870_),
    .X(_07046_));
 sg13g2_buf_1 _23532_ (.A(_06913_),
    .X(_07047_));
 sg13g2_nand2_1 _23533_ (.Y(_07048_),
    .A(\top_ihp.oisc.regs[2][15] ),
    .B(net795));
 sg13g2_a221oi_1 _23534_ (.B2(\top_ihp.oisc.regs[32][15] ),
    .C1(net865),
    .B1(net808),
    .A1(\top_ihp.oisc.regs[14][15] ),
    .Y(_07049_),
    .A2(net748));
 sg13g2_buf_1 _23535_ (.A(_06877_),
    .X(_07050_));
 sg13g2_a22oi_1 _23536_ (.Y(_07051_),
    .B1(net759),
    .B2(\top_ihp.oisc.regs[15][15] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][15] ));
 sg13g2_a22oi_1 _23537_ (.Y(_07052_),
    .B1(net792),
    .B2(\top_ihp.oisc.regs[9][15] ),
    .A2(net787),
    .A1(\top_ihp.oisc.regs[11][15] ));
 sg13g2_nand4_1 _23538_ (.B(_07049_),
    .C(_07051_),
    .A(_07048_),
    .Y(_07053_),
    .D(_07052_));
 sg13g2_a221oi_1 _23539_ (.B2(\top_ihp.oisc.regs[7][15] ),
    .C1(_07053_),
    .B1(net739),
    .A1(\top_ihp.oisc.regs[3][15] ),
    .Y(_07054_),
    .A2(net780));
 sg13g2_nand4_1 _23540_ (.B(_07043_),
    .C(_07045_),
    .A(_07041_),
    .Y(_07055_),
    .D(_07054_));
 sg13g2_a21oi_1 _23541_ (.A1(_00122_),
    .A2(net826),
    .Y(_07056_),
    .B1(net796));
 sg13g2_a21oi_1 _23542_ (.A1(_07055_),
    .A2(_07056_),
    .Y(_07057_),
    .B1(net684));
 sg13g2_a21oi_1 _23543_ (.A1(_07559_),
    .A2(net683),
    .Y(_00332_),
    .B1(_07057_));
 sg13g2_a22oi_1 _23544_ (.Y(_07058_),
    .B1(net742),
    .B2(\top_ihp.oisc.regs[6][16] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][16] ));
 sg13g2_nand2_1 _23545_ (.Y(_07059_),
    .A(\top_ihp.oisc.regs[9][16] ),
    .B(net755));
 sg13g2_a22oi_1 _23546_ (.Y(_07060_),
    .B1(net713),
    .B2(\top_ihp.oisc.regs[15][16] ),
    .A2(net712),
    .A1(\top_ihp.oisc.regs[13][16] ));
 sg13g2_a22oi_1 _23547_ (.Y(_07061_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][16] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][16] ));
 sg13g2_a22oi_1 _23548_ (.Y(_07062_),
    .B1(_06935_),
    .B2(\top_ihp.oisc.regs[8][16] ),
    .A2(_06995_),
    .A1(\top_ihp.oisc.regs[11][16] ));
 sg13g2_a22oi_1 _23549_ (.Y(_07063_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[14][16] ),
    .A2(_06877_),
    .A1(\top_ihp.oisc.regs[10][16] ));
 sg13g2_nand4_1 _23550_ (.B(_07061_),
    .C(_07062_),
    .A(net864),
    .Y(_07064_),
    .D(_07063_));
 sg13g2_a21oi_1 _23551_ (.A1(\top_ihp.oisc.regs[2][16] ),
    .A2(_06966_),
    .Y(_07065_),
    .B1(_07064_));
 sg13g2_nand4_1 _23552_ (.B(_07059_),
    .C(_07060_),
    .A(_07058_),
    .Y(_07066_),
    .D(_07065_));
 sg13g2_a22oi_1 _23553_ (.Y(_07067_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][16] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][16] ));
 sg13g2_a22oi_1 _23554_ (.Y(_07068_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][16] ),
    .A2(net785),
    .A1(\top_ihp.oisc.regs[3][16] ));
 sg13g2_nand2_1 _23555_ (.Y(_07069_),
    .A(_07067_),
    .B(_07068_));
 sg13g2_a21oi_1 _23556_ (.A1(_00123_),
    .A2(_06956_),
    .Y(_07070_),
    .B1(net786));
 sg13g2_o21ai_1 _23557_ (.B1(_07070_),
    .Y(_07071_),
    .A1(_07066_),
    .A2(_07069_));
 sg13g2_nor2_1 _23558_ (.A(_07508_),
    .B(net714),
    .Y(_07072_));
 sg13g2_a21oi_1 _23559_ (.A1(net717),
    .A2(_07071_),
    .Y(_00333_),
    .B1(_07072_));
 sg13g2_and2_1 _23560_ (.A(\top_ihp.oisc.regs[9][17] ),
    .B(net792),
    .X(_07073_));
 sg13g2_a221oi_1 _23561_ (.B2(\top_ihp.oisc.regs[15][17] ),
    .C1(_07073_),
    .B1(net713),
    .A1(\top_ihp.oisc.regs[13][17] ),
    .Y(_07074_),
    .A2(net712));
 sg13g2_nand2_1 _23562_ (.Y(_07075_),
    .A(\top_ihp.oisc.regs[3][17] ),
    .B(_06870_));
 sg13g2_a221oi_1 _23563_ (.B2(\top_ihp.oisc.regs[32][17] ),
    .C1(net848),
    .B1(net808),
    .A1(\top_ihp.oisc.regs[12][17] ),
    .Y(_07076_),
    .A2(_06882_));
 sg13g2_a22oi_1 _23564_ (.Y(_07077_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[8][17] ),
    .A2(net787),
    .A1(\top_ihp.oisc.regs[11][17] ));
 sg13g2_a22oi_1 _23565_ (.Y(_07078_),
    .B1(net760),
    .B2(\top_ihp.oisc.regs[14][17] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][17] ));
 sg13g2_nand4_1 _23566_ (.B(_07076_),
    .C(_07077_),
    .A(_07075_),
    .Y(_07079_),
    .D(_07078_));
 sg13g2_a221oi_1 _23567_ (.B2(\top_ihp.oisc.regs[6][17] ),
    .C1(_07079_),
    .B1(net742),
    .A1(\top_ihp.oisc.regs[7][17] ),
    .Y(_07080_),
    .A2(net739));
 sg13g2_a22oi_1 _23568_ (.Y(_07081_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][17] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][17] ));
 sg13g2_a22oi_1 _23569_ (.Y(_07082_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][17] ),
    .A2(net753),
    .A1(\top_ihp.oisc.regs[2][17] ));
 sg13g2_nand4_1 _23570_ (.B(_07080_),
    .C(_07081_),
    .A(_07074_),
    .Y(_07083_),
    .D(_07082_));
 sg13g2_a21oi_1 _23571_ (.A1(_00124_),
    .A2(net826),
    .Y(_07084_),
    .B1(net796));
 sg13g2_a21oi_1 _23572_ (.A1(_07083_),
    .A2(_07084_),
    .Y(_07085_),
    .B1(net684));
 sg13g2_a21oi_1 _23573_ (.A1(_07558_),
    .A2(net683),
    .Y(_00334_),
    .B1(_07085_));
 sg13g2_a22oi_1 _23574_ (.Y(_07086_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][18] ),
    .A2(net745),
    .A1(\top_ihp.oisc.regs[6][18] ));
 sg13g2_a22oi_1 _23575_ (.Y(_07087_),
    .B1(_06932_),
    .B2(\top_ihp.oisc.regs[4][18] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][18] ));
 sg13g2_and2_1 _23576_ (.A(\top_ihp.oisc.regs[8][18] ),
    .B(net790),
    .X(_07088_));
 sg13g2_a221oi_1 _23577_ (.B2(\top_ihp.oisc.regs[15][18] ),
    .C1(_07088_),
    .B1(net713),
    .A1(\top_ihp.oisc.regs[13][18] ),
    .Y(_07089_),
    .A2(net762));
 sg13g2_nand2_1 _23578_ (.Y(_07090_),
    .A(\top_ihp.oisc.regs[2][18] ),
    .B(net795));
 sg13g2_a221oi_1 _23579_ (.B2(\top_ihp.oisc.regs[32][18] ),
    .C1(net865),
    .B1(net828),
    .A1(\top_ihp.oisc.regs[11][18] ),
    .Y(_07091_),
    .A2(_06893_));
 sg13g2_a22oi_1 _23580_ (.Y(_07092_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][18] ),
    .A2(_07050_),
    .A1(\top_ihp.oisc.regs[10][18] ));
 sg13g2_a22oi_1 _23581_ (.Y(_07093_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][18] ),
    .A2(net752),
    .A1(\top_ihp.oisc.regs[14][18] ));
 sg13g2_nand4_1 _23582_ (.B(_07091_),
    .C(_07092_),
    .A(_07090_),
    .Y(_07094_),
    .D(_07093_));
 sg13g2_a221oi_1 _23583_ (.B2(\top_ihp.oisc.regs[7][18] ),
    .C1(_07094_),
    .B1(net739),
    .A1(\top_ihp.oisc.regs[3][18] ),
    .Y(_07095_),
    .A2(net780));
 sg13g2_nand4_1 _23584_ (.B(_07087_),
    .C(_07089_),
    .A(_07086_),
    .Y(_07096_),
    .D(_07095_));
 sg13g2_a21oi_1 _23585_ (.A1(_00125_),
    .A2(net826),
    .Y(_07097_),
    .B1(net796));
 sg13g2_a21oi_1 _23586_ (.A1(_07096_),
    .A2(_07097_),
    .Y(_07098_),
    .B1(net684));
 sg13g2_a21oi_1 _23587_ (.A1(_07890_),
    .A2(net683),
    .Y(_00335_),
    .B1(_07098_));
 sg13g2_a22oi_1 _23588_ (.Y(_07099_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][19] ),
    .A2(net745),
    .A1(\top_ihp.oisc.regs[6][19] ));
 sg13g2_a22oi_1 _23589_ (.Y(_07100_),
    .B1(_06932_),
    .B2(\top_ihp.oisc.regs[4][19] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][19] ));
 sg13g2_and2_1 _23590_ (.A(\top_ihp.oisc.regs[12][19] ),
    .B(net761),
    .X(_07101_));
 sg13g2_a221oi_1 _23591_ (.B2(\top_ihp.oisc.regs[11][19] ),
    .C1(_07101_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[15][19] ),
    .Y(_07102_),
    .A2(net759));
 sg13g2_nand2_1 _23592_ (.Y(_07103_),
    .A(\top_ihp.oisc.regs[7][19] ),
    .B(_06913_));
 sg13g2_a221oi_1 _23593_ (.B2(\top_ihp.oisc.regs[32][19] ),
    .C1(net865),
    .B1(net828),
    .A1(\top_ihp.oisc.regs[14][19] ),
    .Y(_07104_),
    .A2(net748));
 sg13g2_a22oi_1 _23594_ (.Y(_07105_),
    .B1(net792),
    .B2(\top_ihp.oisc.regs[9][19] ),
    .A2(net810),
    .A1(\top_ihp.oisc.regs[8][19] ));
 sg13g2_a22oi_1 _23595_ (.Y(_07106_),
    .B1(net794),
    .B2(\top_ihp.oisc.regs[10][19] ),
    .A2(net762),
    .A1(\top_ihp.oisc.regs[13][19] ));
 sg13g2_nand4_1 _23596_ (.B(_07104_),
    .C(_07105_),
    .A(_07103_),
    .Y(_07107_),
    .D(_07106_));
 sg13g2_a221oi_1 _23597_ (.B2(\top_ihp.oisc.regs[3][19] ),
    .C1(_07107_),
    .B1(net789),
    .A1(\top_ihp.oisc.regs[2][19] ),
    .Y(_07108_),
    .A2(net749));
 sg13g2_nand4_1 _23598_ (.B(_07100_),
    .C(_07102_),
    .A(_07099_),
    .Y(_07109_),
    .D(_07108_));
 sg13g2_a21oi_1 _23599_ (.A1(_00126_),
    .A2(net826),
    .Y(_07110_),
    .B1(net796));
 sg13g2_a21oi_1 _23600_ (.A1(_07109_),
    .A2(_07110_),
    .Y(_07111_),
    .B1(_06853_));
 sg13g2_a21oi_1 _23601_ (.A1(_07454_),
    .A2(net683),
    .Y(_00336_),
    .B1(_07111_));
 sg13g2_and2_1 _23602_ (.A(\top_ihp.oisc.regs[8][1] ),
    .B(net790),
    .X(_07112_));
 sg13g2_a221oi_1 _23603_ (.B2(\top_ihp.oisc.regs[9][1] ),
    .C1(_07112_),
    .B1(_06939_),
    .A1(\top_ihp.oisc.regs[15][1] ),
    .Y(_07113_),
    .A2(net716));
 sg13g2_nand2_1 _23604_ (.Y(_07114_),
    .A(\top_ihp.oisc.regs[2][1] ),
    .B(net795));
 sg13g2_a221oi_1 _23605_ (.B2(\top_ihp.oisc.regs[32][1] ),
    .C1(net848),
    .B1(_07031_),
    .A1(\top_ihp.oisc.regs[14][1] ),
    .Y(_07115_),
    .A2(net748));
 sg13g2_a22oi_1 _23606_ (.Y(_07116_),
    .B1(net793),
    .B2(\top_ihp.oisc.regs[11][1] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][1] ));
 sg13g2_a22oi_1 _23607_ (.Y(_07117_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][1] ),
    .A2(net762),
    .A1(\top_ihp.oisc.regs[13][1] ));
 sg13g2_nand4_1 _23608_ (.B(_07115_),
    .C(_07116_),
    .A(_07114_),
    .Y(_07118_),
    .D(_07117_));
 sg13g2_a221oi_1 _23609_ (.B2(\top_ihp.oisc.regs[6][1] ),
    .C1(_07118_),
    .B1(net742),
    .A1(\top_ihp.oisc.regs[1][1] ),
    .Y(_07119_),
    .A2(net784));
 sg13g2_a22oi_1 _23610_ (.Y(_07120_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][1] ),
    .A2(net754),
    .A1(\top_ihp.oisc.regs[7][1] ));
 sg13g2_a22oi_1 _23611_ (.Y(_07121_),
    .B1(_06975_),
    .B2(\top_ihp.oisc.regs[4][1] ),
    .A2(net785),
    .A1(\top_ihp.oisc.regs[3][1] ));
 sg13g2_nand4_1 _23612_ (.B(_07119_),
    .C(_07120_),
    .A(_07113_),
    .Y(_07122_),
    .D(_07121_));
 sg13g2_a21oi_1 _23613_ (.A1(_00108_),
    .A2(_07038_),
    .Y(_07123_),
    .B1(net796));
 sg13g2_a21oi_1 _23614_ (.A1(_07122_),
    .A2(_07123_),
    .Y(_07124_),
    .B1(_06853_));
 sg13g2_a21oi_1 _23615_ (.A1(_07850_),
    .A2(_07024_),
    .Y(_00337_),
    .B1(_07124_));
 sg13g2_a22oi_1 _23616_ (.Y(_07125_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][20] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][20] ));
 sg13g2_a22oi_1 _23617_ (.Y(_07126_),
    .B1(net747),
    .B2(\top_ihp.oisc.regs[4][20] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][20] ));
 sg13g2_nand2_1 _23618_ (.Y(_07127_),
    .A(_07125_),
    .B(_07126_));
 sg13g2_nand2_1 _23619_ (.Y(_07128_),
    .A(\top_ihp.oisc.regs[8][20] ),
    .B(net790));
 sg13g2_a22oi_1 _23620_ (.Y(_07129_),
    .B1(net793),
    .B2(\top_ihp.oisc.regs[11][20] ),
    .A2(net716),
    .A1(\top_ihp.oisc.regs[15][20] ));
 sg13g2_a22oi_1 _23621_ (.Y(_07130_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[7][20] ),
    .A2(_06941_),
    .A1(\top_ihp.oisc.regs[3][20] ));
 sg13g2_a22oi_1 _23622_ (.Y(_07131_),
    .B1(_06856_),
    .B2(\top_ihp.oisc.regs[32][20] ),
    .A2(net752),
    .A1(\top_ihp.oisc.regs[14][20] ));
 sg13g2_a22oi_1 _23623_ (.Y(_07132_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][20] ),
    .A2(net788),
    .A1(\top_ihp.oisc.regs[10][20] ));
 sg13g2_a22oi_1 _23624_ (.Y(_07133_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][20] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][20] ));
 sg13g2_nand4_1 _23625_ (.B(_07131_),
    .C(_07132_),
    .A(net847),
    .Y(_07134_),
    .D(_07133_));
 sg13g2_a21oi_1 _23626_ (.A1(\top_ihp.oisc.regs[2][20] ),
    .A2(_06944_),
    .Y(_07135_),
    .B1(_07134_));
 sg13g2_nand4_1 _23627_ (.B(_07129_),
    .C(_07130_),
    .A(_07128_),
    .Y(_07136_),
    .D(_07135_));
 sg13g2_a21oi_1 _23628_ (.A1(_00127_),
    .A2(_06956_),
    .Y(_07137_),
    .B1(_06957_));
 sg13g2_o21ai_1 _23629_ (.B1(_07137_),
    .Y(_07138_),
    .A1(_07127_),
    .A2(_07136_));
 sg13g2_nor2_1 _23630_ (.A(_07452_),
    .B(net714),
    .Y(_07139_));
 sg13g2_a21oi_1 _23631_ (.A1(net717),
    .A2(_07138_),
    .Y(_00338_),
    .B1(_07139_));
 sg13g2_a22oi_1 _23632_ (.Y(_07140_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][21] ),
    .A2(_06928_),
    .A1(\top_ihp.oisc.regs[6][21] ));
 sg13g2_a22oi_1 _23633_ (.Y(_07141_),
    .B1(net747),
    .B2(\top_ihp.oisc.regs[4][21] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][21] ));
 sg13g2_nand2_1 _23634_ (.Y(_07142_),
    .A(_07140_),
    .B(_07141_));
 sg13g2_nand2_1 _23635_ (.Y(_07143_),
    .A(\top_ihp.oisc.regs[14][21] ),
    .B(net760));
 sg13g2_a22oi_1 _23636_ (.Y(_07144_),
    .B1(_06894_),
    .B2(\top_ihp.oisc.regs[11][21] ),
    .A2(net716),
    .A1(\top_ihp.oisc.regs[15][21] ));
 sg13g2_a22oi_1 _23637_ (.Y(_07145_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[7][21] ),
    .A2(net789),
    .A1(\top_ihp.oisc.regs[3][21] ));
 sg13g2_a22oi_1 _23638_ (.Y(_07146_),
    .B1(_06898_),
    .B2(\top_ihp.oisc.regs[8][21] ),
    .A2(net808),
    .A1(\top_ihp.oisc.regs[32][21] ));
 sg13g2_a22oi_1 _23639_ (.Y(_07147_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][21] ),
    .A2(net788),
    .A1(\top_ihp.oisc.regs[10][21] ));
 sg13g2_a22oi_1 _23640_ (.Y(_07148_),
    .B1(net740),
    .B2(\top_ihp.oisc.regs[12][21] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][21] ));
 sg13g2_nand4_1 _23641_ (.B(_07146_),
    .C(_07147_),
    .A(net847),
    .Y(_07149_),
    .D(_07148_));
 sg13g2_a21oi_1 _23642_ (.A1(\top_ihp.oisc.regs[2][21] ),
    .A2(net753),
    .Y(_07150_),
    .B1(_07149_));
 sg13g2_nand4_1 _23643_ (.B(_07144_),
    .C(_07145_),
    .A(_07143_),
    .Y(_07151_),
    .D(_07150_));
 sg13g2_buf_1 _23644_ (.A(net812),
    .X(_07152_));
 sg13g2_a21oi_1 _23645_ (.A1(_00128_),
    .A2(net827),
    .Y(_07153_),
    .B1(net778));
 sg13g2_o21ai_1 _23646_ (.B1(_07153_),
    .Y(_07154_),
    .A1(_07142_),
    .A2(_07151_));
 sg13g2_nor2_1 _23647_ (.A(_07462_),
    .B(net714),
    .Y(_07155_));
 sg13g2_a21oi_1 _23648_ (.A1(net717),
    .A2(_07154_),
    .Y(_00339_),
    .B1(_07155_));
 sg13g2_a22oi_1 _23649_ (.Y(_07156_),
    .B1(net785),
    .B2(\top_ihp.oisc.regs[3][22] ),
    .A2(net784),
    .A1(\top_ihp.oisc.regs[1][22] ));
 sg13g2_nand2_1 _23650_ (.Y(_07157_),
    .A(\top_ihp.oisc.regs[9][22] ),
    .B(net755));
 sg13g2_a22oi_1 _23651_ (.Y(_07158_),
    .B1(net713),
    .B2(\top_ihp.oisc.regs[15][22] ),
    .A2(net712),
    .A1(\top_ihp.oisc.regs[13][22] ));
 sg13g2_a22oi_1 _23652_ (.Y(_07159_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][22] ),
    .A2(_07016_),
    .A1(\top_ihp.oisc.regs[12][22] ));
 sg13g2_a22oi_1 _23653_ (.Y(_07160_),
    .B1(net810),
    .B2(\top_ihp.oisc.regs[8][22] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][22] ));
 sg13g2_a22oi_1 _23654_ (.Y(_07161_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[14][22] ),
    .A2(_06877_),
    .A1(\top_ihp.oisc.regs[10][22] ));
 sg13g2_nand4_1 _23655_ (.B(_07159_),
    .C(_07160_),
    .A(net864),
    .Y(_07162_),
    .D(_07161_));
 sg13g2_a21oi_1 _23656_ (.A1(\top_ihp.oisc.regs[2][22] ),
    .A2(net749),
    .Y(_07163_),
    .B1(_07162_));
 sg13g2_nand4_1 _23657_ (.B(_07157_),
    .C(_07158_),
    .A(_07156_),
    .Y(_07164_),
    .D(_07163_));
 sg13g2_a22oi_1 _23658_ (.Y(_07165_),
    .B1(_06976_),
    .B2(\top_ihp.oisc.regs[5][22] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][22] ));
 sg13g2_a22oi_1 _23659_ (.Y(_07166_),
    .B1(net745),
    .B2(\top_ihp.oisc.regs[6][22] ),
    .A2(_06942_),
    .A1(\top_ihp.oisc.regs[7][22] ));
 sg13g2_nand2_1 _23660_ (.Y(_07167_),
    .A(_07165_),
    .B(_07166_));
 sg13g2_buf_1 _23661_ (.A(_06906_),
    .X(_07168_));
 sg13g2_a21oi_1 _23662_ (.A1(_00129_),
    .A2(net825),
    .Y(_07169_),
    .B1(net778));
 sg13g2_o21ai_1 _23663_ (.B1(_07169_),
    .Y(_07170_),
    .A1(_07164_),
    .A2(_07167_));
 sg13g2_nor2_1 _23664_ (.A(_07445_),
    .B(net714),
    .Y(_07171_));
 sg13g2_a21oi_1 _23665_ (.A1(net717),
    .A2(_07170_),
    .Y(_00340_),
    .B1(_07171_));
 sg13g2_a22oi_1 _23666_ (.Y(_07172_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][23] ),
    .A2(_06987_),
    .A1(\top_ihp.oisc.regs[6][23] ));
 sg13g2_a22oi_1 _23667_ (.Y(_07173_),
    .B1(net747),
    .B2(\top_ihp.oisc.regs[4][23] ),
    .A2(_06931_),
    .A1(\top_ihp.oisc.regs[1][23] ));
 sg13g2_nand2_1 _23668_ (.Y(_07174_),
    .A(_07172_),
    .B(_07173_));
 sg13g2_nand2_1 _23669_ (.Y(_07175_),
    .A(\top_ihp.oisc.regs[12][23] ),
    .B(net761));
 sg13g2_a22oi_1 _23670_ (.Y(_07176_),
    .B1(net713),
    .B2(\top_ihp.oisc.regs[15][23] ),
    .A2(net712),
    .A1(\top_ihp.oisc.regs[13][23] ));
 sg13g2_a22oi_1 _23671_ (.Y(_07177_),
    .B1(_06942_),
    .B2(\top_ihp.oisc.regs[7][23] ),
    .A2(_06941_),
    .A1(\top_ihp.oisc.regs[3][23] ));
 sg13g2_a22oi_1 _23672_ (.Y(_07178_),
    .B1(net812),
    .B2(\top_ihp.oisc.regs[32][23] ),
    .A2(_06945_),
    .A1(\top_ihp.oisc.regs[14][23] ));
 sg13g2_a22oi_1 _23673_ (.Y(_07179_),
    .B1(_06948_),
    .B2(\top_ihp.oisc.regs[11][23] ),
    .A2(_06947_),
    .A1(\top_ihp.oisc.regs[10][23] ));
 sg13g2_a22oi_1 _23674_ (.Y(_07180_),
    .B1(_06998_),
    .B2(\top_ihp.oisc.regs[9][23] ),
    .A2(_06897_),
    .A1(\top_ihp.oisc.regs[8][23] ));
 sg13g2_nand4_1 _23675_ (.B(_07178_),
    .C(_07179_),
    .A(net847),
    .Y(_07181_),
    .D(_07180_));
 sg13g2_a21oi_1 _23676_ (.A1(\top_ihp.oisc.regs[2][23] ),
    .A2(net749),
    .Y(_07182_),
    .B1(_07181_));
 sg13g2_nand4_1 _23677_ (.B(_07176_),
    .C(_07177_),
    .A(_07175_),
    .Y(_07183_),
    .D(_07182_));
 sg13g2_a21oi_1 _23678_ (.A1(_00130_),
    .A2(net825),
    .Y(_07184_),
    .B1(net778));
 sg13g2_o21ai_1 _23679_ (.B1(_07184_),
    .Y(_07185_),
    .A1(_07174_),
    .A2(_07183_));
 sg13g2_nor2_1 _23680_ (.A(_07443_),
    .B(net714),
    .Y(_07186_));
 sg13g2_a21oi_1 _23681_ (.A1(_06927_),
    .A2(_07185_),
    .Y(_00341_),
    .B1(_07186_));
 sg13g2_and2_1 _23682_ (.A(\top_ihp.oisc.regs[12][24] ),
    .B(net761),
    .X(_07187_));
 sg13g2_a221oi_1 _23683_ (.B2(\top_ihp.oisc.regs[11][24] ),
    .C1(_07187_),
    .B1(_06894_),
    .A1(\top_ihp.oisc.regs[15][24] ),
    .Y(_07188_),
    .A2(net716));
 sg13g2_nand2_1 _23684_ (.Y(_07189_),
    .A(\top_ihp.oisc.regs[2][24] ),
    .B(_06866_));
 sg13g2_a221oi_1 _23685_ (.B2(\top_ihp.oisc.regs[32][24] ),
    .C1(_06906_),
    .B1(_07031_),
    .A1(\top_ihp.oisc.regs[14][24] ),
    .Y(_07190_),
    .A2(net748));
 sg13g2_a22oi_1 _23686_ (.Y(_07191_),
    .B1(net792),
    .B2(\top_ihp.oisc.regs[9][24] ),
    .A2(net811),
    .A1(\top_ihp.oisc.regs[8][24] ));
 sg13g2_a22oi_1 _23687_ (.Y(_07192_),
    .B1(net794),
    .B2(\top_ihp.oisc.regs[10][24] ),
    .A2(net762),
    .A1(\top_ihp.oisc.regs[13][24] ));
 sg13g2_nand4_1 _23688_ (.B(_07190_),
    .C(_07191_),
    .A(_07189_),
    .Y(_07193_),
    .D(_07192_));
 sg13g2_a221oi_1 _23689_ (.B2(\top_ihp.oisc.regs[3][24] ),
    .C1(_07193_),
    .B1(net785),
    .A1(\top_ihp.oisc.regs[1][24] ),
    .Y(_07194_),
    .A2(net784));
 sg13g2_a22oi_1 _23690_ (.Y(_07195_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][24] ),
    .A2(net754),
    .A1(\top_ihp.oisc.regs[7][24] ));
 sg13g2_a22oi_1 _23691_ (.Y(_07196_),
    .B1(net745),
    .B2(\top_ihp.oisc.regs[6][24] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][24] ));
 sg13g2_nand4_1 _23692_ (.B(_07194_),
    .C(_07195_),
    .A(_07188_),
    .Y(_07197_),
    .D(_07196_));
 sg13g2_a21oi_1 _23693_ (.A1(_00131_),
    .A2(_07038_),
    .Y(_07198_),
    .B1(_06857_));
 sg13g2_a21oi_1 _23694_ (.A1(_07197_),
    .A2(_07198_),
    .Y(_07199_),
    .B1(_03692_));
 sg13g2_a21oi_1 _23695_ (.A1(_07613_),
    .A2(net683),
    .Y(_00342_),
    .B1(_07199_));
 sg13g2_a22oi_1 _23696_ (.Y(_07200_),
    .B1(_06929_),
    .B2(\top_ihp.oisc.regs[5][25] ),
    .A2(net742),
    .A1(\top_ihp.oisc.regs[6][25] ));
 sg13g2_a22oi_1 _23697_ (.Y(_07201_),
    .B1(_06975_),
    .B2(\top_ihp.oisc.regs[4][25] ),
    .A2(_06931_),
    .A1(\top_ihp.oisc.regs[1][25] ));
 sg13g2_nand2_1 _23698_ (.Y(_07202_),
    .A(_07200_),
    .B(_07201_));
 sg13g2_nand2_1 _23699_ (.Y(_07203_),
    .A(\top_ihp.oisc.regs[8][25] ),
    .B(net790));
 sg13g2_a22oi_1 _23700_ (.Y(_07204_),
    .B1(_07011_),
    .B2(\top_ihp.oisc.regs[15][25] ),
    .A2(_07027_),
    .A1(\top_ihp.oisc.regs[13][25] ));
 sg13g2_a22oi_1 _23701_ (.Y(_07205_),
    .B1(_07047_),
    .B2(\top_ihp.oisc.regs[7][25] ),
    .A2(net789),
    .A1(\top_ihp.oisc.regs[3][25] ));
 sg13g2_a22oi_1 _23702_ (.Y(_07206_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][25] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][25] ));
 sg13g2_a22oi_1 _23703_ (.Y(_07207_),
    .B1(_06951_),
    .B2(\top_ihp.oisc.regs[12][25] ),
    .A2(_06947_),
    .A1(\top_ihp.oisc.regs[10][25] ));
 sg13g2_a22oi_1 _23704_ (.Y(_07208_),
    .B1(_06998_),
    .B2(\top_ihp.oisc.regs[9][25] ),
    .A2(_06967_),
    .A1(\top_ihp.oisc.regs[14][25] ));
 sg13g2_nand4_1 _23705_ (.B(_07206_),
    .C(_07207_),
    .A(net847),
    .Y(_07209_),
    .D(_07208_));
 sg13g2_a21oi_1 _23706_ (.A1(\top_ihp.oisc.regs[2][25] ),
    .A2(net749),
    .Y(_07210_),
    .B1(_07209_));
 sg13g2_nand4_1 _23707_ (.B(_07204_),
    .C(_07205_),
    .A(_07203_),
    .Y(_07211_),
    .D(_07210_));
 sg13g2_a21oi_1 _23708_ (.A1(_00132_),
    .A2(net825),
    .Y(_07212_),
    .B1(net778));
 sg13g2_o21ai_1 _23709_ (.B1(_07212_),
    .Y(_07213_),
    .A1(_07202_),
    .A2(_07211_));
 sg13g2_nor2_1 _23710_ (.A(_07622_),
    .B(net714),
    .Y(_07214_));
 sg13g2_a21oi_1 _23711_ (.A1(_06927_),
    .A2(_07213_),
    .Y(_00343_),
    .B1(_07214_));
 sg13g2_a22oi_1 _23712_ (.Y(_07215_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][26] ),
    .A2(net753),
    .A1(\top_ihp.oisc.regs[2][26] ));
 sg13g2_nand2_1 _23713_ (.Y(_07216_),
    .A(\top_ihp.oisc.regs[14][26] ),
    .B(net760));
 sg13g2_a22oi_1 _23714_ (.Y(_07217_),
    .B1(_07011_),
    .B2(\top_ihp.oisc.regs[15][26] ),
    .A2(net794),
    .A1(\top_ihp.oisc.regs[10][26] ));
 sg13g2_a22oi_1 _23715_ (.Y(_07218_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][26] ),
    .A2(net808),
    .A1(\top_ihp.oisc.regs[32][26] ));
 sg13g2_a22oi_1 _23716_ (.Y(_07219_),
    .B1(net787),
    .B2(\top_ihp.oisc.regs[11][26] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][26] ));
 sg13g2_a22oi_1 _23717_ (.Y(_07220_),
    .B1(_06897_),
    .B2(\top_ihp.oisc.regs[8][26] ),
    .A2(_06874_),
    .A1(\top_ihp.oisc.regs[13][26] ));
 sg13g2_nand4_1 _23718_ (.B(_07218_),
    .C(_07219_),
    .A(net864),
    .Y(_07221_),
    .D(_07220_));
 sg13g2_a21oi_1 _23719_ (.A1(\top_ihp.oisc.regs[3][26] ),
    .A2(_07046_),
    .Y(_07222_),
    .B1(_07221_));
 sg13g2_nand4_1 _23720_ (.B(_07216_),
    .C(_07217_),
    .A(_07215_),
    .Y(_07223_),
    .D(_07222_));
 sg13g2_a22oi_1 _23721_ (.Y(_07224_),
    .B1(net745),
    .B2(\top_ihp.oisc.regs[6][26] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][26] ));
 sg13g2_a22oi_1 _23722_ (.Y(_07225_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][26] ),
    .A2(_07042_),
    .A1(\top_ihp.oisc.regs[1][26] ));
 sg13g2_nand2_1 _23723_ (.Y(_07226_),
    .A(_07224_),
    .B(_07225_));
 sg13g2_a21oi_1 _23724_ (.A1(_00133_),
    .A2(_07168_),
    .Y(_07227_),
    .B1(_07152_));
 sg13g2_o21ai_1 _23725_ (.B1(_07227_),
    .Y(_07228_),
    .A1(_07223_),
    .A2(_07226_));
 sg13g2_nor2_1 _23726_ (.A(_07615_),
    .B(_07005_),
    .Y(_07229_));
 sg13g2_a21oi_1 _23727_ (.A1(net715),
    .A2(_07228_),
    .Y(_00344_),
    .B1(_07229_));
 sg13g2_a22oi_1 _23728_ (.Y(_07230_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][27] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][27] ));
 sg13g2_a22oi_1 _23729_ (.Y(_07231_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][27] ),
    .A2(net742),
    .A1(\top_ihp.oisc.regs[6][27] ));
 sg13g2_nand2_1 _23730_ (.Y(_07232_),
    .A(_07230_),
    .B(_07231_));
 sg13g2_nand2_1 _23731_ (.Y(_07233_),
    .A(\top_ihp.oisc.regs[9][27] ),
    .B(_06939_));
 sg13g2_a22oi_1 _23732_ (.Y(_07234_),
    .B1(_06878_),
    .B2(\top_ihp.oisc.regs[10][27] ),
    .A2(_07027_),
    .A1(\top_ihp.oisc.regs[13][27] ));
 sg13g2_a22oi_1 _23733_ (.Y(_07235_),
    .B1(net785),
    .B2(\top_ihp.oisc.regs[3][27] ),
    .A2(net784),
    .A1(\top_ihp.oisc.regs[1][27] ));
 sg13g2_a22oi_1 _23734_ (.Y(_07236_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][27] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][27] ));
 sg13g2_a22oi_1 _23735_ (.Y(_07237_),
    .B1(_06935_),
    .B2(\top_ihp.oisc.regs[8][27] ),
    .A2(_06890_),
    .A1(\top_ihp.oisc.regs[15][27] ));
 sg13g2_a22oi_1 _23736_ (.Y(_07238_),
    .B1(_06945_),
    .B2(\top_ihp.oisc.regs[14][27] ),
    .A2(_07016_),
    .A1(\top_ihp.oisc.regs[12][27] ));
 sg13g2_nand4_1 _23737_ (.B(_07236_),
    .C(_07237_),
    .A(_06924_),
    .Y(_07239_),
    .D(_07238_));
 sg13g2_a21oi_1 _23738_ (.A1(\top_ihp.oisc.regs[2][27] ),
    .A2(net749),
    .Y(_07240_),
    .B1(_07239_));
 sg13g2_nand4_1 _23739_ (.B(_07234_),
    .C(_07235_),
    .A(_07233_),
    .Y(_07241_),
    .D(_07240_));
 sg13g2_a21oi_1 _23740_ (.A1(_00134_),
    .A2(_07168_),
    .Y(_07242_),
    .B1(_07152_));
 sg13g2_o21ai_1 _23741_ (.B1(_07242_),
    .Y(_07243_),
    .A1(_07232_),
    .A2(_07241_));
 sg13g2_nor2_1 _23742_ (.A(_07682_),
    .B(_07005_),
    .Y(_07244_));
 sg13g2_a21oi_1 _23743_ (.A1(net715),
    .A2(_07243_),
    .Y(_00345_),
    .B1(_07244_));
 sg13g2_a22oi_1 _23744_ (.Y(_07245_),
    .B1(_06985_),
    .B2(\top_ihp.oisc.regs[7][28] ),
    .A2(_06984_),
    .A1(\top_ihp.oisc.regs[4][28] ));
 sg13g2_a22oi_1 _23745_ (.Y(_07246_),
    .B1(_06978_),
    .B2(\top_ihp.oisc.regs[6][28] ),
    .A2(_06962_),
    .A1(\top_ihp.oisc.regs[3][28] ));
 sg13g2_nand2_1 _23746_ (.Y(_07247_),
    .A(_07245_),
    .B(_07246_));
 sg13g2_nand2_1 _23747_ (.Y(_07248_),
    .A(\top_ihp.oisc.regs[14][28] ),
    .B(net760));
 sg13g2_a22oi_1 _23748_ (.Y(_07249_),
    .B1(net755),
    .B2(\top_ihp.oisc.regs[9][28] ),
    .A2(net716),
    .A1(\top_ihp.oisc.regs[15][28] ));
 sg13g2_a22oi_1 _23749_ (.Y(_07250_),
    .B1(_06944_),
    .B2(\top_ihp.oisc.regs[2][28] ),
    .A2(_06993_),
    .A1(\top_ihp.oisc.regs[1][28] ));
 sg13g2_a22oi_1 _23750_ (.Y(_07251_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][28] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][28] ));
 sg13g2_a22oi_1 _23751_ (.Y(_07252_),
    .B1(_06951_),
    .B2(\top_ihp.oisc.regs[12][28] ),
    .A2(net788),
    .A1(\top_ihp.oisc.regs[10][28] ));
 sg13g2_a22oi_1 _23752_ (.Y(_07253_),
    .B1(net810),
    .B2(\top_ihp.oisc.regs[8][28] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][28] ));
 sg13g2_nand4_1 _23753_ (.B(_07251_),
    .C(_07252_),
    .A(net847),
    .Y(_07254_),
    .D(_07253_));
 sg13g2_a21oi_1 _23754_ (.A1(\top_ihp.oisc.regs[5][28] ),
    .A2(_06988_),
    .Y(_07255_),
    .B1(_07254_));
 sg13g2_nand4_1 _23755_ (.B(_07249_),
    .C(_07250_),
    .A(_07248_),
    .Y(_07256_),
    .D(_07255_));
 sg13g2_a21oi_1 _23756_ (.A1(_00135_),
    .A2(net825),
    .Y(_07257_),
    .B1(net778));
 sg13g2_o21ai_1 _23757_ (.B1(_07257_),
    .Y(_07258_),
    .A1(_07247_),
    .A2(_07256_));
 sg13g2_nor2_1 _23758_ (.A(_07680_),
    .B(net773),
    .Y(_07259_));
 sg13g2_a21oi_1 _23759_ (.A1(net715),
    .A2(_07258_),
    .Y(_00346_),
    .B1(_07259_));
 sg13g2_a22oi_1 _23760_ (.Y(_07260_),
    .B1(_06985_),
    .B2(\top_ihp.oisc.regs[7][29] ),
    .A2(_06984_),
    .A1(\top_ihp.oisc.regs[4][29] ));
 sg13g2_a22oi_1 _23761_ (.Y(_07261_),
    .B1(_06988_),
    .B2(\top_ihp.oisc.regs[5][29] ),
    .A2(_06987_),
    .A1(\top_ihp.oisc.regs[6][29] ));
 sg13g2_nand2_1 _23762_ (.Y(_07262_),
    .A(_07260_),
    .B(_07261_));
 sg13g2_nand2_1 _23763_ (.Y(_07263_),
    .A(\top_ihp.oisc.regs[8][29] ),
    .B(_06936_));
 sg13g2_a22oi_1 _23764_ (.Y(_07264_),
    .B1(_06883_),
    .B2(\top_ihp.oisc.regs[12][29] ),
    .A2(_06878_),
    .A1(\top_ihp.oisc.regs[10][29] ));
 sg13g2_a22oi_1 _23765_ (.Y(_07265_),
    .B1(_06962_),
    .B2(\top_ihp.oisc.regs[3][29] ),
    .A2(_06993_),
    .A1(\top_ihp.oisc.regs[1][29] ));
 sg13g2_a22oi_1 _23766_ (.Y(_07266_),
    .B1(_06968_),
    .B2(\top_ihp.oisc.regs[32][29] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][29] ));
 sg13g2_a22oi_1 _23767_ (.Y(_07267_),
    .B1(_06891_),
    .B2(\top_ihp.oisc.regs[15][29] ),
    .A2(_06967_),
    .A1(\top_ihp.oisc.regs[14][29] ));
 sg13g2_a22oi_1 _23768_ (.Y(_07268_),
    .B1(_06901_),
    .B2(\top_ihp.oisc.regs[9][29] ),
    .A2(_06950_),
    .A1(\top_ihp.oisc.regs[13][29] ));
 sg13g2_nand4_1 _23769_ (.B(_07266_),
    .C(_07267_),
    .A(_06923_),
    .Y(_07269_),
    .D(_07268_));
 sg13g2_a21oi_1 _23770_ (.A1(\top_ihp.oisc.regs[2][29] ),
    .A2(_06966_),
    .Y(_07270_),
    .B1(_07269_));
 sg13g2_nand4_1 _23771_ (.B(_07264_),
    .C(_07265_),
    .A(_07263_),
    .Y(_07271_),
    .D(_07270_));
 sg13g2_a21oi_1 _23772_ (.A1(_00136_),
    .A2(net825),
    .Y(_07272_),
    .B1(net778));
 sg13g2_o21ai_1 _23773_ (.B1(_07272_),
    .Y(_07273_),
    .A1(_07262_),
    .A2(_07271_));
 sg13g2_nor2_1 _23774_ (.A(_07722_),
    .B(_03680_),
    .Y(_07274_));
 sg13g2_a21oi_1 _23775_ (.A1(_06960_),
    .A2(_07273_),
    .Y(_00347_),
    .B1(_07274_));
 sg13g2_a22oi_1 _23776_ (.Y(_07275_),
    .B1(_06976_),
    .B2(\top_ihp.oisc.regs[5][2] ),
    .A2(_06978_),
    .A1(\top_ihp.oisc.regs[6][2] ));
 sg13g2_a22oi_1 _23777_ (.Y(_07276_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][2] ),
    .A2(_07042_),
    .A1(\top_ihp.oisc.regs[1][2] ));
 sg13g2_and2_1 _23778_ (.A(\top_ihp.oisc.regs[8][2] ),
    .B(_06936_),
    .X(_07277_));
 sg13g2_a221oi_1 _23779_ (.B2(\top_ihp.oisc.regs[15][2] ),
    .C1(_07277_),
    .B1(_06938_),
    .A1(\top_ihp.oisc.regs[12][2] ),
    .Y(_07278_),
    .A2(_06883_));
 sg13g2_nand2_1 _23780_ (.Y(_07279_),
    .A(\top_ihp.oisc.regs[2][2] ),
    .B(_06865_));
 sg13g2_a221oi_1 _23781_ (.B2(\top_ihp.oisc.regs[32][2] ),
    .C1(_06905_),
    .B1(_06855_),
    .A1(\top_ihp.oisc.regs[14][2] ),
    .Y(_07280_),
    .A2(net748));
 sg13g2_a22oi_1 _23782_ (.Y(_07281_),
    .B1(_06902_),
    .B2(\top_ihp.oisc.regs[9][2] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][2] ));
 sg13g2_a22oi_1 _23783_ (.Y(_07282_),
    .B1(_06948_),
    .B2(\top_ihp.oisc.regs[11][2] ),
    .A2(_06875_),
    .A1(\top_ihp.oisc.regs[13][2] ));
 sg13g2_nand4_1 _23784_ (.B(_07280_),
    .C(_07281_),
    .A(_07279_),
    .Y(_07283_),
    .D(_07282_));
 sg13g2_a221oi_1 _23785_ (.B2(\top_ihp.oisc.regs[7][2] ),
    .C1(_07283_),
    .B1(_07047_),
    .A1(\top_ihp.oisc.regs[3][2] ),
    .Y(_07284_),
    .A2(net780));
 sg13g2_nand4_1 _23786_ (.B(_07276_),
    .C(_07278_),
    .A(_07275_),
    .Y(_07285_),
    .D(_07284_));
 sg13g2_a21oi_1 _23787_ (.A1(_00109_),
    .A2(net826),
    .Y(_07286_),
    .B1(_06857_));
 sg13g2_a21oi_1 _23788_ (.A1(_07285_),
    .A2(_07286_),
    .Y(_07287_),
    .B1(net709));
 sg13g2_a21oi_1 _23789_ (.A1(_07847_),
    .A2(_07024_),
    .Y(_00348_),
    .B1(_07287_));
 sg13g2_a22oi_1 _23790_ (.Y(_07288_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][30] ),
    .A2(net742),
    .A1(\top_ihp.oisc.regs[6][30] ));
 sg13g2_a22oi_1 _23791_ (.Y(_07289_),
    .B1(net747),
    .B2(\top_ihp.oisc.regs[4][30] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][30] ));
 sg13g2_nand2_1 _23792_ (.Y(_07290_),
    .A(_07288_),
    .B(_07289_));
 sg13g2_nand2_1 _23793_ (.Y(_07291_),
    .A(\top_ihp.oisc.regs[14][30] ),
    .B(net760));
 sg13g2_a22oi_1 _23794_ (.Y(_07292_),
    .B1(net755),
    .B2(\top_ihp.oisc.regs[9][30] ),
    .A2(_06938_),
    .A1(\top_ihp.oisc.regs[15][30] ));
 sg13g2_a22oi_1 _23795_ (.Y(_07293_),
    .B1(net739),
    .B2(\top_ihp.oisc.regs[7][30] ),
    .A2(net789),
    .A1(\top_ihp.oisc.regs[3][30] ));
 sg13g2_a22oi_1 _23796_ (.Y(_07294_),
    .B1(_06968_),
    .B2(\top_ihp.oisc.regs[32][30] ),
    .A2(_06995_),
    .A1(\top_ihp.oisc.regs[11][30] ));
 sg13g2_a22oi_1 _23797_ (.Y(_07295_),
    .B1(net810),
    .B2(\top_ihp.oisc.regs[8][30] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][30] ));
 sg13g2_a22oi_1 _23798_ (.Y(_07296_),
    .B1(_07050_),
    .B2(\top_ihp.oisc.regs[10][30] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][30] ));
 sg13g2_nand4_1 _23799_ (.B(_07294_),
    .C(_07295_),
    .A(net864),
    .Y(_07297_),
    .D(_07296_));
 sg13g2_a21oi_1 _23800_ (.A1(\top_ihp.oisc.regs[2][30] ),
    .A2(net749),
    .Y(_07298_),
    .B1(_07297_));
 sg13g2_nand4_1 _23801_ (.B(_07292_),
    .C(_07293_),
    .A(_07291_),
    .Y(_07299_),
    .D(_07298_));
 sg13g2_a21oi_1 _23802_ (.A1(_00137_),
    .A2(net825),
    .Y(_07300_),
    .B1(net778));
 sg13g2_o21ai_1 _23803_ (.B1(_07300_),
    .Y(_07301_),
    .A1(_07290_),
    .A2(_07299_));
 sg13g2_nor2_1 _23804_ (.A(_07719_),
    .B(net773),
    .Y(_07302_));
 sg13g2_a21oi_1 _23805_ (.A1(_06960_),
    .A2(_07301_),
    .Y(_00349_),
    .B1(_07302_));
 sg13g2_a22oi_1 _23806_ (.Y(_07303_),
    .B1(net753),
    .B2(\top_ihp.oisc.regs[2][31] ),
    .A2(net784),
    .A1(\top_ihp.oisc.regs[1][31] ));
 sg13g2_nand2_1 _23807_ (.Y(_07304_),
    .A(\top_ihp.oisc.regs[14][31] ),
    .B(net760));
 sg13g2_a22oi_1 _23808_ (.Y(_07305_),
    .B1(net755),
    .B2(\top_ihp.oisc.regs[9][31] ),
    .A2(net793),
    .A1(\top_ihp.oisc.regs[11][31] ));
 sg13g2_a22oi_1 _23809_ (.Y(_07306_),
    .B1(net810),
    .B2(\top_ihp.oisc.regs[8][31] ),
    .A2(net808),
    .A1(\top_ihp.oisc.regs[32][31] ));
 sg13g2_a22oi_1 _23810_ (.Y(_07307_),
    .B1(_06890_),
    .B2(\top_ihp.oisc.regs[15][31] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][31] ));
 sg13g2_a22oi_1 _23811_ (.Y(_07308_),
    .B1(net788),
    .B2(\top_ihp.oisc.regs[10][31] ),
    .A2(_06874_),
    .A1(\top_ihp.oisc.regs[13][31] ));
 sg13g2_nand4_1 _23812_ (.B(_07306_),
    .C(_07307_),
    .A(net864),
    .Y(_07309_),
    .D(_07308_));
 sg13g2_a21oi_1 _23813_ (.A1(\top_ihp.oisc.regs[3][31] ),
    .A2(_07046_),
    .Y(_07310_),
    .B1(_07309_));
 sg13g2_nand4_1 _23814_ (.B(_07304_),
    .C(_07305_),
    .A(_07303_),
    .Y(_07311_),
    .D(_07310_));
 sg13g2_a22oi_1 _23815_ (.Y(_07312_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][31] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][31] ));
 sg13g2_a22oi_1 _23816_ (.Y(_07313_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][31] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][31] ));
 sg13g2_nand2_1 _23817_ (.Y(_07314_),
    .A(_07312_),
    .B(_07313_));
 sg13g2_a21oi_1 _23818_ (.A1(_00068_),
    .A2(net825),
    .Y(_07315_),
    .B1(net778));
 sg13g2_o21ai_1 _23819_ (.B1(_07315_),
    .Y(_07316_),
    .A1(_07311_),
    .A2(_07314_));
 sg13g2_nor2_1 _23820_ (.A(\top_ihp.oisc.op_b[31] ),
    .B(net773),
    .Y(_07317_));
 sg13g2_a21oi_1 _23821_ (.A1(net715),
    .A2(_07316_),
    .Y(_00350_),
    .B1(_07317_));
 sg13g2_a22oi_1 _23822_ (.Y(_07318_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][3] ),
    .A2(net742),
    .A1(\top_ihp.oisc.regs[6][3] ));
 sg13g2_a22oi_1 _23823_ (.Y(_07319_),
    .B1(net747),
    .B2(\top_ihp.oisc.regs[4][3] ),
    .A2(net791),
    .A1(\top_ihp.oisc.regs[1][3] ));
 sg13g2_nand2_1 _23824_ (.Y(_07320_),
    .A(_07318_),
    .B(_07319_));
 sg13g2_nand2_1 _23825_ (.Y(_07321_),
    .A(\top_ihp.oisc.regs[8][3] ),
    .B(net790));
 sg13g2_a22oi_1 _23826_ (.Y(_07322_),
    .B1(net713),
    .B2(\top_ihp.oisc.regs[15][3] ),
    .A2(net712),
    .A1(\top_ihp.oisc.regs[13][3] ));
 sg13g2_a22oi_1 _23827_ (.Y(_07323_),
    .B1(net739),
    .B2(\top_ihp.oisc.regs[7][3] ),
    .A2(net780),
    .A1(\top_ihp.oisc.regs[3][3] ));
 sg13g2_a22oi_1 _23828_ (.Y(_07324_),
    .B1(net809),
    .B2(\top_ihp.oisc.regs[32][3] ),
    .A2(net783),
    .A1(\top_ihp.oisc.regs[11][3] ));
 sg13g2_a22oi_1 _23829_ (.Y(_07325_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][3] ),
    .A2(net788),
    .A1(\top_ihp.oisc.regs[10][3] ));
 sg13g2_a22oi_1 _23830_ (.Y(_07326_),
    .B1(_06901_),
    .B2(\top_ihp.oisc.regs[9][3] ),
    .A2(net748),
    .A1(\top_ihp.oisc.regs[14][3] ));
 sg13g2_nand4_1 _23831_ (.B(_07324_),
    .C(_07325_),
    .A(net864),
    .Y(_07327_),
    .D(_07326_));
 sg13g2_a21oi_1 _23832_ (.A1(\top_ihp.oisc.regs[2][3] ),
    .A2(net749),
    .Y(_07328_),
    .B1(_07327_));
 sg13g2_nand4_1 _23833_ (.B(_07322_),
    .C(_07323_),
    .A(_07321_),
    .Y(_07329_),
    .D(_07328_));
 sg13g2_a21oi_1 _23834_ (.A1(_00110_),
    .A2(net825),
    .Y(_07330_),
    .B1(net812));
 sg13g2_o21ai_1 _23835_ (.B1(_07330_),
    .Y(_07331_),
    .A1(_07320_),
    .A2(_07329_));
 sg13g2_nor2_1 _23836_ (.A(_07485_),
    .B(net773),
    .Y(_07332_));
 sg13g2_a21oi_1 _23837_ (.A1(net715),
    .A2(_07331_),
    .Y(_00351_),
    .B1(_07332_));
 sg13g2_a22oi_1 _23838_ (.Y(_07333_),
    .B1(net753),
    .B2(\top_ihp.oisc.regs[2][4] ),
    .A2(net784),
    .A1(\top_ihp.oisc.regs[1][4] ));
 sg13g2_nand2_1 _23839_ (.Y(_07334_),
    .A(\top_ihp.oisc.regs[14][4] ),
    .B(net760));
 sg13g2_a22oi_1 _23840_ (.Y(_07335_),
    .B1(net755),
    .B2(\top_ihp.oisc.regs[9][4] ),
    .A2(net793),
    .A1(\top_ihp.oisc.regs[11][4] ));
 sg13g2_a22oi_1 _23841_ (.Y(_07336_),
    .B1(net810),
    .B2(\top_ihp.oisc.regs[8][4] ),
    .A2(net808),
    .A1(\top_ihp.oisc.regs[32][4] ));
 sg13g2_a22oi_1 _23842_ (.Y(_07337_),
    .B1(_06890_),
    .B2(\top_ihp.oisc.regs[15][4] ),
    .A2(net740),
    .A1(\top_ihp.oisc.regs[12][4] ));
 sg13g2_a22oi_1 _23843_ (.Y(_07338_),
    .B1(net788),
    .B2(\top_ihp.oisc.regs[10][4] ),
    .A2(_06874_),
    .A1(\top_ihp.oisc.regs[13][4] ));
 sg13g2_nand4_1 _23844_ (.B(_07336_),
    .C(_07337_),
    .A(net864),
    .Y(_07339_),
    .D(_07338_));
 sg13g2_a21oi_1 _23845_ (.A1(\top_ihp.oisc.regs[3][4] ),
    .A2(net780),
    .Y(_07340_),
    .B1(_07339_));
 sg13g2_nand4_1 _23846_ (.B(_07334_),
    .C(_07335_),
    .A(_07333_),
    .Y(_07341_),
    .D(_07340_));
 sg13g2_a22oi_1 _23847_ (.Y(_07342_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][4] ),
    .A2(net744),
    .A1(\top_ihp.oisc.regs[4][4] ));
 sg13g2_a22oi_1 _23848_ (.Y(_07343_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[5][4] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][4] ));
 sg13g2_nand2_1 _23849_ (.Y(_07344_),
    .A(_07342_),
    .B(_07343_));
 sg13g2_a21oi_1 _23850_ (.A1(_00111_),
    .A2(net848),
    .Y(_07345_),
    .B1(net812));
 sg13g2_o21ai_1 _23851_ (.B1(_07345_),
    .Y(_07346_),
    .A1(_07341_),
    .A2(_07344_));
 sg13g2_nor2_1 _23852_ (.A(_07486_),
    .B(net773),
    .Y(_07347_));
 sg13g2_a21oi_1 _23853_ (.A1(net715),
    .A2(_07346_),
    .Y(_00352_),
    .B1(_07347_));
 sg13g2_a22oi_1 _23854_ (.Y(_07348_),
    .B1(net743),
    .B2(\top_ihp.oisc.regs[7][5] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][5] ));
 sg13g2_a22oi_1 _23855_ (.Y(_07349_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][5] ),
    .A2(net785),
    .A1(\top_ihp.oisc.regs[3][5] ));
 sg13g2_and2_1 _23856_ (.A(\top_ihp.oisc.regs[8][5] ),
    .B(net811),
    .X(_07350_));
 sg13g2_a221oi_1 _23857_ (.B2(\top_ihp.oisc.regs[9][5] ),
    .C1(_07350_),
    .B1(net755),
    .A1(\top_ihp.oisc.regs[10][5] ),
    .Y(_07351_),
    .A2(net794));
 sg13g2_nand2_1 _23858_ (.Y(_07352_),
    .A(\top_ihp.oisc.regs[5][5] ),
    .B(_06918_));
 sg13g2_a221oi_1 _23859_ (.B2(\top_ihp.oisc.regs[32][5] ),
    .C1(net865),
    .B1(net828),
    .A1(\top_ihp.oisc.regs[15][5] ),
    .Y(_07353_),
    .A2(_06890_));
 sg13g2_a22oi_1 _23860_ (.Y(_07354_),
    .B1(net787),
    .B2(\top_ihp.oisc.regs[11][5] ),
    .A2(net752),
    .A1(\top_ihp.oisc.regs[14][5] ));
 sg13g2_a22oi_1 _23861_ (.Y(_07355_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][5] ),
    .A2(net762),
    .A1(\top_ihp.oisc.regs[13][5] ));
 sg13g2_nand4_1 _23862_ (.B(_07353_),
    .C(_07354_),
    .A(_07352_),
    .Y(_07356_),
    .D(_07355_));
 sg13g2_a221oi_1 _23863_ (.B2(\top_ihp.oisc.regs[6][5] ),
    .C1(_07356_),
    .B1(_06916_),
    .A1(\top_ihp.oisc.regs[2][5] ),
    .Y(_07357_),
    .A2(net795));
 sg13g2_nand4_1 _23864_ (.B(_07349_),
    .C(_07351_),
    .A(_07348_),
    .Y(_07358_),
    .D(_07357_));
 sg13g2_a21oi_1 _23865_ (.A1(_00112_),
    .A2(net826),
    .Y(_07359_),
    .B1(net796));
 sg13g2_a21oi_1 _23866_ (.A1(_07358_),
    .A2(_07359_),
    .Y(_07360_),
    .B1(net709));
 sg13g2_a21oi_1 _23867_ (.A1(_07502_),
    .A2(net683),
    .Y(_00353_),
    .B1(_07360_));
 sg13g2_a22oi_1 _23868_ (.Y(_07361_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][6] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][6] ));
 sg13g2_a22oi_1 _23869_ (.Y(_07362_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][6] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][6] ));
 sg13g2_and2_1 _23870_ (.A(\top_ihp.oisc.regs[8][6] ),
    .B(net811),
    .X(_07363_));
 sg13g2_a221oi_1 _23871_ (.B2(\top_ihp.oisc.regs[11][6] ),
    .C1(_07363_),
    .B1(net793),
    .A1(\top_ihp.oisc.regs[15][6] ),
    .Y(_07364_),
    .A2(net759));
 sg13g2_nand2_1 _23872_ (.Y(_07365_),
    .A(\top_ihp.oisc.regs[2][6] ),
    .B(_06865_));
 sg13g2_a221oi_1 _23873_ (.B2(\top_ihp.oisc.regs[32][6] ),
    .C1(net865),
    .B1(net828),
    .A1(\top_ihp.oisc.regs[14][6] ),
    .Y(_07366_),
    .A2(_06885_));
 sg13g2_a22oi_1 _23874_ (.Y(_07367_),
    .B1(net792),
    .B2(\top_ihp.oisc.regs[9][6] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][6] ));
 sg13g2_a22oi_1 _23875_ (.Y(_07368_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][6] ),
    .A2(net751),
    .A1(\top_ihp.oisc.regs[13][6] ));
 sg13g2_nand4_1 _23876_ (.B(_07366_),
    .C(_07367_),
    .A(_07365_),
    .Y(_07369_),
    .D(_07368_));
 sg13g2_a221oi_1 _23877_ (.B2(\top_ihp.oisc.regs[7][6] ),
    .C1(_07369_),
    .B1(net739),
    .A1(\top_ihp.oisc.regs[3][6] ),
    .Y(_07370_),
    .A2(net780));
 sg13g2_nand4_1 _23878_ (.B(_07362_),
    .C(_07364_),
    .A(_07361_),
    .Y(_07371_),
    .D(_07370_));
 sg13g2_a21oi_1 _23879_ (.A1(_00113_),
    .A2(net826),
    .Y(_07372_),
    .B1(net786));
 sg13g2_a21oi_1 _23880_ (.A1(_07371_),
    .A2(_07372_),
    .Y(_07373_),
    .B1(net709));
 sg13g2_a21oi_1 _23881_ (.A1(_07552_),
    .A2(net683),
    .Y(_00354_),
    .B1(_07373_));
 sg13g2_a22oi_1 _23882_ (.Y(_07374_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][7] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][7] ));
 sg13g2_a22oi_1 _23883_ (.Y(_07375_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][7] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][7] ));
 sg13g2_and2_1 _23884_ (.A(\top_ihp.oisc.regs[8][7] ),
    .B(net811),
    .X(_07376_));
 sg13g2_a221oi_1 _23885_ (.B2(\top_ihp.oisc.regs[15][7] ),
    .C1(_07376_),
    .B1(net716),
    .A1(\top_ihp.oisc.regs[13][7] ),
    .Y(_07377_),
    .A2(net762));
 sg13g2_nand2_1 _23886_ (.Y(_07378_),
    .A(\top_ihp.oisc.regs[2][7] ),
    .B(_06865_));
 sg13g2_a221oi_1 _23887_ (.B2(\top_ihp.oisc.regs[32][7] ),
    .C1(net865),
    .B1(net828),
    .A1(\top_ihp.oisc.regs[11][7] ),
    .Y(_07379_),
    .A2(_06893_));
 sg13g2_a22oi_1 _23888_ (.Y(_07380_),
    .B1(net750),
    .B2(\top_ihp.oisc.regs[12][7] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][7] ));
 sg13g2_a22oi_1 _23889_ (.Y(_07381_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][7] ),
    .A2(net752),
    .A1(\top_ihp.oisc.regs[14][7] ));
 sg13g2_nand4_1 _23890_ (.B(_07379_),
    .C(_07380_),
    .A(_07378_),
    .Y(_07382_),
    .D(_07381_));
 sg13g2_a221oi_1 _23891_ (.B2(\top_ihp.oisc.regs[7][7] ),
    .C1(_07382_),
    .B1(net739),
    .A1(\top_ihp.oisc.regs[3][7] ),
    .Y(_07383_),
    .A2(net780));
 sg13g2_nand4_1 _23892_ (.B(_07375_),
    .C(_07377_),
    .A(_07374_),
    .Y(_07384_),
    .D(_07383_));
 sg13g2_a21oi_1 _23893_ (.A1(_00114_),
    .A2(net827),
    .Y(_07385_),
    .B1(net786));
 sg13g2_a21oi_1 _23894_ (.A1(_07384_),
    .A2(_07385_),
    .Y(_07386_),
    .B1(net709));
 sg13g2_a21oi_1 _23895_ (.A1(_07583_),
    .A2(net684),
    .Y(_00355_),
    .B1(_07386_));
 sg13g2_and2_1 _23896_ (.A(\top_ihp.oisc.regs[9][8] ),
    .B(net792),
    .X(_07387_));
 sg13g2_a221oi_1 _23897_ (.B2(\top_ihp.oisc.regs[15][8] ),
    .C1(_07387_),
    .B1(net713),
    .A1(\top_ihp.oisc.regs[13][8] ),
    .Y(_07388_),
    .A2(net712));
 sg13g2_nand2_1 _23898_ (.Y(_07389_),
    .A(\top_ihp.oisc.regs[2][8] ),
    .B(net795));
 sg13g2_a221oi_1 _23899_ (.B2(\top_ihp.oisc.regs[32][8] ),
    .C1(net848),
    .B1(net808),
    .A1(\top_ihp.oisc.regs[12][8] ),
    .Y(_07390_),
    .A2(_06882_));
 sg13g2_a22oi_1 _23900_ (.Y(_07391_),
    .B1(net811),
    .B2(\top_ihp.oisc.regs[8][8] ),
    .A2(net787),
    .A1(\top_ihp.oisc.regs[11][8] ));
 sg13g2_a22oi_1 _23901_ (.Y(_07392_),
    .B1(net760),
    .B2(\top_ihp.oisc.regs[14][8] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][8] ));
 sg13g2_nand4_1 _23902_ (.B(_07390_),
    .C(_07391_),
    .A(_07389_),
    .Y(_07393_),
    .D(_07392_));
 sg13g2_a221oi_1 _23903_ (.B2(\top_ihp.oisc.regs[3][8] ),
    .C1(_07393_),
    .B1(net789),
    .A1(\top_ihp.oisc.regs[1][8] ),
    .Y(_07394_),
    .A2(net784));
 sg13g2_a22oi_1 _23904_ (.Y(_07395_),
    .B1(net741),
    .B2(\top_ihp.oisc.regs[5][8] ),
    .A2(net754),
    .A1(\top_ihp.oisc.regs[7][8] ));
 sg13g2_a22oi_1 _23905_ (.Y(_07396_),
    .B1(net745),
    .B2(\top_ihp.oisc.regs[6][8] ),
    .A2(_06911_),
    .A1(\top_ihp.oisc.regs[4][8] ));
 sg13g2_nand4_1 _23906_ (.B(_07394_),
    .C(_07395_),
    .A(_07388_),
    .Y(_07397_),
    .D(_07396_));
 sg13g2_a21oi_1 _23907_ (.A1(_00115_),
    .A2(net827),
    .Y(_07398_),
    .B1(net786));
 sg13g2_a21oi_1 _23908_ (.A1(_07397_),
    .A2(_07398_),
    .Y(_07399_),
    .B1(net709));
 sg13g2_a21oi_1 _23909_ (.A1(_07581_),
    .A2(net684),
    .Y(_00356_),
    .B1(_07399_));
 sg13g2_a22oi_1 _23910_ (.Y(_07400_),
    .B1(net746),
    .B2(\top_ihp.oisc.regs[5][9] ),
    .A2(net758),
    .A1(\top_ihp.oisc.regs[6][9] ));
 sg13g2_a22oi_1 _23911_ (.Y(_07401_),
    .B1(net756),
    .B2(\top_ihp.oisc.regs[4][9] ),
    .A2(net781),
    .A1(\top_ihp.oisc.regs[1][9] ));
 sg13g2_and2_1 _23912_ (.A(\top_ihp.oisc.regs[12][9] ),
    .B(net761),
    .X(_07402_));
 sg13g2_a221oi_1 _23913_ (.B2(\top_ihp.oisc.regs[15][9] ),
    .C1(_07402_),
    .B1(net716),
    .A1(\top_ihp.oisc.regs[13][9] ),
    .Y(_07403_),
    .A2(net762));
 sg13g2_nand2_1 _23914_ (.Y(_07404_),
    .A(\top_ihp.oisc.regs[2][9] ),
    .B(_06865_));
 sg13g2_a221oi_1 _23915_ (.B2(\top_ihp.oisc.regs[32][9] ),
    .C1(net865),
    .B1(net828),
    .A1(\top_ihp.oisc.regs[14][9] ),
    .Y(_07405_),
    .A2(_06885_));
 sg13g2_a22oi_1 _23916_ (.Y(_07406_),
    .B1(net787),
    .B2(\top_ihp.oisc.regs[11][9] ),
    .A2(net779),
    .A1(\top_ihp.oisc.regs[10][9] ));
 sg13g2_a22oi_1 _23917_ (.Y(_07407_),
    .B1(net782),
    .B2(\top_ihp.oisc.regs[9][9] ),
    .A2(net810),
    .A1(\top_ihp.oisc.regs[8][9] ));
 sg13g2_nand4_1 _23918_ (.B(_07405_),
    .C(_07406_),
    .A(_07404_),
    .Y(_07408_),
    .D(_07407_));
 sg13g2_a221oi_1 _23919_ (.B2(\top_ihp.oisc.regs[7][9] ),
    .C1(_07408_),
    .B1(net739),
    .A1(\top_ihp.oisc.regs[3][9] ),
    .Y(_07409_),
    .A2(net780));
 sg13g2_nand4_1 _23920_ (.B(_07401_),
    .C(_07403_),
    .A(_07400_),
    .Y(_07410_),
    .D(_07409_));
 sg13g2_a21oi_1 _23921_ (.A1(_00116_),
    .A2(net827),
    .Y(_07411_),
    .B1(net786));
 sg13g2_a21oi_1 _23922_ (.A1(_07410_),
    .A2(_07411_),
    .Y(_07412_),
    .B1(net709));
 sg13g2_a21oi_1 _23923_ (.A1(_07592_),
    .A2(net684),
    .Y(_00357_),
    .B1(_07412_));
 sg13g2_a21oi_1 _23924_ (.A1(_07713_),
    .A2(_07741_),
    .Y(_00229_),
    .B1(_08213_));
 sg13g2_mux4_1 _23925_ (.S0(_08043_),
    .A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ),
    .A2(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ),
    .A3(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ),
    .S1(_08044_),
    .X(_07413_));
 sg13g2_mux4_1 _23926_ (.S0(_08043_),
    .A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ),
    .A2(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ),
    .A3(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ),
    .S1(_08044_),
    .X(_07414_));
 sg13g2_mux2_1 _23927_ (.A0(_07413_),
    .A1(_07414_),
    .S(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .X(_07415_));
 sg13g2_nand2b_1 _23928_ (.Y(_07416_),
    .B(_08040_),
    .A_N(net1024));
 sg13g2_o21ai_1 _23929_ (.B1(_07416_),
    .Y(_00230_),
    .A1(_04518_),
    .A2(_07415_));
 sg13g2_nor2_1 _23930_ (.A(net907),
    .B(net2097),
    .Y(\top_ihp.ram_clk_o ));
 sg13g2_and2_1 _23931_ (.A(_03933_),
    .B(\top_ihp.wb_emem.cmd[63] ),
    .X(\top_ihp.ram_data_o ));
 sg13g2_nor2_1 _23932_ (.A(net2096),
    .B(\top_ihp.rom_cs_o ),
    .Y(\top_ihp.rom_clk_o ));
 sg13g2_and2_1 _23933_ (.A(_07750_),
    .B(\top_ihp.wb_dati_rom[7] ),
    .X(\top_ihp.rom_data_o ));
 sg13g2_and2_1 _23934_ (.A(net983),
    .B(\top_ihp.wb_dati_spi[31] ),
    .X(\top_ihp.spi_data_o ));
 sg13g2_inv_1 _14128__1 (.Y(net1980),
    .A(clknet_leaf_57_clk));
 sg13g2_buf_1 _23936_ (.A(net1395),
    .X(uio_oe[0]));
 sg13g2_buf_1 _23937_ (.A(net1396),
    .X(uio_oe[1]));
 sg13g2_buf_1 _23938_ (.A(net1397),
    .X(uio_oe[2]));
 sg13g2_buf_1 _23939_ (.A(net1398),
    .X(uio_oe[3]));
 sg13g2_buf_1 _23940_ (.A(net1399),
    .X(uio_oe[4]));
 sg13g2_buf_1 _23941_ (.A(net1400),
    .X(uio_oe[5]));
 sg13g2_buf_1 _23942_ (.A(net1401),
    .X(uio_oe[6]));
 sg13g2_buf_1 _23943_ (.A(net1402),
    .X(uio_oe[7]));
 sg13g2_buf_1 _23944_ (.A(\top_ihp.spi_data_o ),
    .X(net9));
 sg13g2_buf_1 _23945_ (.A(\top_ihp.spi_cs_o_1 ),
    .X(net10));
 sg13g2_buf_1 _23946_ (.A(\top_ihp.spi_cs_o_2 ),
    .X(net11));
 sg13g2_buf_1 _23947_ (.A(\top_ihp.spi_cs_o_3 ),
    .X(net12));
 sg13g2_buf_1 _23948_ (.A(\top_ihp.gpio_o_1 ),
    .X(net13));
 sg13g2_buf_1 _23949_ (.A(\top_ihp.gpio_o_2 ),
    .X(net14));
 sg13g2_buf_1 _23950_ (.A(\top_ihp.gpio_o_3 ),
    .X(net15));
 sg13g2_buf_1 _23951_ (.A(\top_ihp.gpio_o_4 ),
    .X(net16));
 sg13g2_buf_1 _23952_ (.A(\top_ihp.tx ),
    .X(net17));
 sg13g2_buf_1 _23953_ (.A(\top_ihp.rom_clk_o ),
    .X(net18));
 sg13g2_buf_1 _23954_ (.A(\top_ihp.rom_data_o ),
    .X(net19));
 sg13g2_buf_1 _23955_ (.A(\top_ihp.rom_cs_o ),
    .X(net20));
 sg13g2_buf_1 _23956_ (.A(\top_ihp.ram_clk_o ),
    .X(net21));
 sg13g2_buf_1 _23957_ (.A(\top_ihp.ram_data_o ),
    .X(net22));
 sg13g2_buf_1 _23958_ (.A(\top_ihp.ram_cs_o ),
    .X(net23));
 sg13g2_buf_1 _23959_ (.A(\top_ihp.spi_clk_o ),
    .X(net24));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_00231_),
    .Q_N(_13128_),
    .Q(\top_ihp.oisc.decoder.decoded[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_00232_),
    .Q_N(_13127_),
    .Q(\top_ihp.oisc.decoder.decoded[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1100),
    .D(_00233_),
    .Q_N(_13126_),
    .Q(\top_ihp.oisc.decoder.decoded[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1100),
    .D(_00234_),
    .Q_N(_13125_),
    .Q(\top_ihp.oisc.decoder.decoded[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1100),
    .D(_00235_),
    .Q_N(_13124_),
    .Q(\top_ihp.oisc.decoder.decoded[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1100),
    .D(_00236_),
    .Q_N(_13123_),
    .Q(\top_ihp.oisc.decoder.decoded[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1100),
    .D(_00237_),
    .Q_N(_00073_),
    .Q(\top_ihp.oisc.decoder.decoded[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1098),
    .D(_00238_),
    .Q_N(_13122_),
    .Q(\top_ihp.oisc.decoder.decoded[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_00239_),
    .Q_N(_13121_),
    .Q(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1092),
    .D(_00240_),
    .Q_N(_13120_),
    .Q(\top_ihp.oisc.decoder.decoded[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1102),
    .D(_00241_),
    .Q_N(_13119_),
    .Q(\top_ihp.oisc.decoder.decoded[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1092),
    .D(_00242_),
    .Q_N(_13118_),
    .Q(\top_ihp.oisc.decoder.decoded[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1098),
    .D(_00243_),
    .Q_N(_13117_),
    .Q(\top_ihp.oisc.decoder.decoded[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1098),
    .D(_00244_),
    .Q_N(_13116_),
    .Q(\top_ihp.oisc.decoder.decoded[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1100),
    .D(_00245_),
    .Q_N(_13115_),
    .Q(\top_ihp.oisc.decoder.instruction[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1104),
    .D(_00246_),
    .Q_N(_13114_),
    .Q(\top_ihp.oisc.decoder.instruction[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1095),
    .D(_00247_),
    .Q_N(_13113_),
    .Q(\top_ihp.oisc.decoder.instruction[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1096),
    .D(_00248_),
    .Q_N(_13112_),
    .Q(\top_ihp.oisc.decoder.instruction[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1095),
    .D(_00249_),
    .Q_N(_00070_),
    .Q(\top_ihp.oisc.decoder.instruction[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1095),
    .D(_00107_),
    .Q_N(_13111_),
    .Q(\top_ihp.oisc.decoder.instruction[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1097),
    .D(_00250_),
    .Q_N(_00103_),
    .Q(\top_ihp.oisc.decoder.instruction[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1097),
    .D(_00251_),
    .Q_N(_00104_),
    .Q(\top_ihp.oisc.decoder.instruction[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1097),
    .D(_00252_),
    .Q_N(_00105_),
    .Q(\top_ihp.oisc.decoder.instruction[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1095),
    .D(_00253_),
    .Q_N(_00106_),
    .Q(\top_ihp.oisc.decoder.instruction[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1105),
    .D(_00254_),
    .Q_N(_13110_),
    .Q(\top_ihp.oisc.decoder.instruction[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1104),
    .D(_00255_),
    .Q_N(_00099_),
    .Q(\top_ihp.oisc.decoder.instruction[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1105),
    .D(_00256_),
    .Q_N(_00100_),
    .Q(\top_ihp.oisc.decoder.instruction[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1105),
    .D(_00257_),
    .Q_N(_00101_),
    .Q(\top_ihp.oisc.decoder.instruction[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1104),
    .D(_00258_),
    .Q_N(_00102_),
    .Q(\top_ihp.oisc.decoder.instruction[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1078),
    .D(_00259_),
    .Q_N(_13109_),
    .Q(\top_ihp.oisc.decoder.instruction[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1078),
    .D(_00260_),
    .Q_N(_13108_),
    .Q(\top_ihp.oisc.decoder.instruction[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_00261_),
    .Q_N(_13107_),
    .Q(\top_ihp.oisc.decoder.instruction[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1078),
    .D(_00262_),
    .Q_N(_13106_),
    .Q(\top_ihp.oisc.decoder.instruction[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1078),
    .D(_00263_),
    .Q_N(_13105_),
    .Q(\top_ihp.oisc.decoder.instruction[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1097),
    .D(_00264_),
    .Q_N(_13104_),
    .Q(\top_ihp.oisc.decoder.instruction[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_00265_),
    .Q_N(_13103_),
    .Q(\top_ihp.oisc.decoder.instruction[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1100),
    .D(_00266_),
    .Q_N(_13102_),
    .Q(\top_ihp.oisc.decoder.instruction[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1104),
    .D(_00267_),
    .Q_N(_13101_),
    .Q(\top_ihp.oisc.decoder.instruction[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1100),
    .D(_00268_),
    .Q_N(_13129_),
    .Q(\top_ihp.oisc.decoder.instruction[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.mem_addr_lowbits[0]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1403),
    .D(\top_ihp.oisc.wb_adr_o[0] ),
    .Q_N(_13130_),
    .Q(\top_ihp.oisc.mem_addr_lowbits[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.mem_addr_lowbits[1]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1404),
    .D(\top_ihp.oisc.wb_adr_o[1] ),
    .Q_N(_13100_),
    .Q(\top_ihp.oisc.mem_addr_lowbits[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1092),
    .D(_00269_),
    .Q_N(_13099_),
    .Q(\top_ihp.oisc.micro_op[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1098),
    .D(_00270_),
    .Q_N(_13098_),
    .Q(\top_ihp.oisc.micro_op[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1092),
    .D(_00271_),
    .Q_N(_13097_),
    .Q(\top_ihp.oisc.micro_op[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1098),
    .D(_00272_),
    .Q_N(_13096_),
    .Q(\top_ihp.oisc.micro_op[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1098),
    .D(_00273_),
    .Q_N(_13095_),
    .Q(\top_ihp.oisc.micro_op[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1098),
    .D(_00274_),
    .Q_N(_13094_),
    .Q(\top_ihp.oisc.micro_op[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1092),
    .D(_00275_),
    .Q_N(_13093_),
    .Q(\top_ihp.oisc.micro_op[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1092),
    .D(_00276_),
    .Q_N(_13092_),
    .Q(\top_ihp.oisc.micro_op[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1092),
    .D(_00277_),
    .Q_N(_13091_),
    .Q(\top_ihp.oisc.micro_op[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1092),
    .D(_00278_),
    .Q_N(_13090_),
    .Q(\top_ihp.oisc.micro_op[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1099),
    .D(_00279_),
    .Q_N(_13089_),
    .Q(\top_ihp.oisc.micro_op[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1093),
    .D(_00280_),
    .Q_N(_13088_),
    .Q(\top_ihp.oisc.micro_op[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1098),
    .D(_00281_),
    .Q_N(_13087_),
    .Q(\top_ihp.oisc.micro_op[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1099),
    .D(_00282_),
    .Q_N(_13086_),
    .Q(\top_ihp.oisc.micro_op[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1405),
    .D(_00283_),
    .Q_N(_00087_),
    .Q(\top_ihp.oisc.micro_pc[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1406),
    .D(_00284_),
    .Q_N(_00088_),
    .Q(\top_ihp.oisc.micro_pc[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1407),
    .D(_00285_),
    .Q_N(_00086_),
    .Q(\top_ihp.oisc.micro_pc[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1408),
    .D(_00286_),
    .Q_N(_00085_),
    .Q(\top_ihp.oisc.micro_pc[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1409),
    .D(_00287_),
    .Q_N(_00084_),
    .Q(\top_ihp.oisc.micro_pc[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1410),
    .D(_00288_),
    .Q_N(_00083_),
    .Q(\top_ihp.oisc.micro_pc[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1411),
    .D(_00289_),
    .Q_N(_00082_),
    .Q(\top_ihp.oisc.micro_pc[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1412),
    .D(_00290_),
    .Q_N(_00081_),
    .Q(\top_ihp.oisc.micro_pc[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[0]$_DFF_PN0_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1145),
    .D(\top_ihp.oisc.reg_rb[0] ),
    .Q_N(_13131_),
    .Q(\top_ihp.oisc.micro_res_addr[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[1]$_DFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1145),
    .D(\top_ihp.oisc.reg_rb[1] ),
    .Q_N(_13132_),
    .Q(\top_ihp.oisc.micro_res_addr[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[2]$_DFF_PN0_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1145),
    .D(\top_ihp.oisc.reg_rb[2] ),
    .Q_N(_13133_),
    .Q(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[3]$_DFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1145),
    .D(\top_ihp.oisc.reg_rb[3] ),
    .Q_N(_13085_),
    .Q(\top_ihp.oisc.micro_res_addr[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1103),
    .D(_00291_),
    .Q_N(\top_ihp.oisc.micro_state[0] ),
    .Q(_13204_));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1103),
    .D(_00292_),
    .Q_N(_13084_),
    .Q(\top_ihp.oisc.micro_state[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1103),
    .D(_00293_),
    .Q_N(_13083_),
    .Q(\top_ihp.oisc.micro_state[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1144),
    .D(_00294_),
    .Q_N(_13082_),
    .Q(\top_ihp.oisc.op_a[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1174),
    .D(_00295_),
    .Q_N(_13081_),
    .Q(\top_ihp.oisc.op_a[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1107),
    .D(_00296_),
    .Q_N(_13080_),
    .Q(\top_ihp.oisc.op_a[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1176),
    .D(_00297_),
    .Q_N(_13079_),
    .Q(\top_ihp.oisc.op_a[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1228),
    .D(_00298_),
    .Q_N(_13078_),
    .Q(\top_ihp.oisc.op_a[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1113),
    .D(_00299_),
    .Q_N(_13077_),
    .Q(\top_ihp.oisc.op_a[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1107),
    .D(_00300_),
    .Q_N(_13076_),
    .Q(\top_ihp.oisc.op_a[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1228),
    .D(_00301_),
    .Q_N(_13075_),
    .Q(\top_ihp.oisc.op_a[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1181),
    .D(_00302_),
    .Q_N(_13074_),
    .Q(\top_ihp.oisc.op_a[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1187),
    .D(_00303_),
    .Q_N(_13073_),
    .Q(\top_ihp.oisc.op_a[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1186),
    .D(_00304_),
    .Q_N(_13072_),
    .Q(\top_ihp.oisc.op_a[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1139),
    .D(_00305_),
    .Q_N(_13071_),
    .Q(\top_ihp.oisc.op_a[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1257),
    .D(_00306_),
    .Q_N(_13070_),
    .Q(\top_ihp.oisc.op_a[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1140),
    .D(_00307_),
    .Q_N(_13069_),
    .Q(\top_ihp.oisc.op_a[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1241),
    .D(_00308_),
    .Q_N(_13068_),
    .Q(\top_ihp.oisc.op_a[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1238),
    .D(_00309_),
    .Q_N(_13067_),
    .Q(\top_ihp.oisc.op_a[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1233),
    .D(_00310_),
    .Q_N(_13066_),
    .Q(\top_ihp.oisc.op_a[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1144),
    .D(_00311_),
    .Q_N(_13065_),
    .Q(\top_ihp.oisc.op_a[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1248),
    .D(_00312_),
    .Q_N(_13064_),
    .Q(\top_ihp.oisc.op_a[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1238),
    .D(_00313_),
    .Q_N(_13063_),
    .Q(\top_ihp.oisc.op_a[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1238),
    .D(_00314_),
    .Q_N(_13062_),
    .Q(\top_ihp.oisc.op_a[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1231),
    .D(_00315_),
    .Q_N(_13061_),
    .Q(\top_ihp.oisc.op_a[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1139),
    .D(_00316_),
    .Q_N(_13060_),
    .Q(\top_ihp.oisc.op_a[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1228),
    .D(_00317_),
    .Q_N(_13059_),
    .Q(\top_ihp.oisc.op_a[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1187),
    .D(_00318_),
    .Q_N(_13058_),
    .Q(\top_ihp.oisc.op_a[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1112),
    .D(_00319_),
    .Q_N(_13057_),
    .Q(\top_ihp.oisc.op_a[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1114),
    .D(_00320_),
    .Q_N(_13056_),
    .Q(\top_ihp.oisc.op_a[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1186),
    .D(_00321_),
    .Q_N(_13055_),
    .Q(\top_ihp.oisc.op_a[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1107),
    .D(_00322_),
    .Q_N(_13054_),
    .Q(\top_ihp.oisc.op_a[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1107),
    .D(_00323_),
    .Q_N(_13053_),
    .Q(\top_ihp.oisc.op_a[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1107),
    .D(_00324_),
    .Q_N(_13052_),
    .Q(\top_ihp.oisc.op_a[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1178),
    .D(_00325_),
    .Q_N(_13051_),
    .Q(\top_ihp.oisc.op_a[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1139),
    .D(_00326_),
    .Q_N(_13050_),
    .Q(\top_ihp.oisc.op_b[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1113),
    .D(_00327_),
    .Q_N(_13049_),
    .Q(\top_ihp.oisc.op_b[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1113),
    .D(_00328_),
    .Q_N(_13048_),
    .Q(\top_ihp.oisc.op_b[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1113),
    .D(_00329_),
    .Q_N(_13047_),
    .Q(\top_ihp.oisc.op_b[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1113),
    .D(_00330_),
    .Q_N(_13046_),
    .Q(\top_ihp.oisc.op_b[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1081),
    .D(_00331_),
    .Q_N(_13045_),
    .Q(\top_ihp.oisc.op_b[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1073),
    .D(_00332_),
    .Q_N(_13044_),
    .Q(\top_ihp.oisc.op_b[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1112),
    .D(_00333_),
    .Q_N(_13043_),
    .Q(\top_ihp.oisc.op_b[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1113),
    .D(_00334_),
    .Q_N(_13042_),
    .Q(\top_ihp.oisc.op_b[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1112),
    .D(_00335_),
    .Q_N(_13041_),
    .Q(\top_ihp.oisc.op_b[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1112),
    .D(_00336_),
    .Q_N(_13040_),
    .Q(\top_ihp.oisc.op_b[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1139),
    .D(_00337_),
    .Q_N(_13039_),
    .Q(\top_ihp.oisc.op_b[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1139),
    .D(_00338_),
    .Q_N(_13038_),
    .Q(\top_ihp.oisc.op_b[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1139),
    .D(_00339_),
    .Q_N(_13037_),
    .Q(\top_ihp.oisc.op_b[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1144),
    .D(_00340_),
    .Q_N(_13036_),
    .Q(\top_ihp.oisc.op_b[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1145),
    .D(_00341_),
    .Q_N(_13035_),
    .Q(\top_ihp.oisc.op_b[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1139),
    .D(_00342_),
    .Q_N(_13034_),
    .Q(\top_ihp.oisc.op_b[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1144),
    .D(_00343_),
    .Q_N(_13033_),
    .Q(\top_ihp.oisc.op_b[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1143),
    .D(_00344_),
    .Q_N(_13032_),
    .Q(\top_ihp.oisc.op_b[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1144),
    .D(_00345_),
    .Q_N(_13031_),
    .Q(\top_ihp.oisc.op_b[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1144),
    .D(_00346_),
    .Q_N(_13030_),
    .Q(\top_ihp.oisc.op_b[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1144),
    .D(_00347_),
    .Q_N(_13029_),
    .Q(\top_ihp.oisc.op_b[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1139),
    .D(_00348_),
    .Q_N(_13028_),
    .Q(\top_ihp.oisc.op_b[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1144),
    .D(_00349_),
    .Q_N(_13027_),
    .Q(\top_ihp.oisc.op_b[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1112),
    .D(_00350_),
    .Q_N(_13026_),
    .Q(\top_ihp.oisc.op_b[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1112),
    .D(_00351_),
    .Q_N(_13025_),
    .Q(\top_ihp.oisc.op_b[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1112),
    .D(_00352_),
    .Q_N(_13024_),
    .Q(\top_ihp.oisc.op_b[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1113),
    .D(_00353_),
    .Q_N(_13023_),
    .Q(\top_ihp.oisc.op_b[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1107),
    .D(_00354_),
    .Q_N(_13022_),
    .Q(\top_ihp.oisc.op_b[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1107),
    .D(_00355_),
    .Q_N(_13021_),
    .Q(\top_ihp.oisc.op_b[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1107),
    .D(_00356_),
    .Q_N(_13020_),
    .Q(\top_ihp.oisc.op_b[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1108),
    .D(_00357_),
    .Q_N(_13019_),
    .Q(\top_ihp.oisc.op_b[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1235),
    .D(_00358_),
    .Q_N(_13018_),
    .Q(\top_ihp.oisc.regs[0][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1171),
    .D(_00359_),
    .Q_N(_00117_),
    .Q(\top_ihp.oisc.regs[0][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1171),
    .D(_00360_),
    .Q_N(_00118_),
    .Q(\top_ihp.oisc.regs[0][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1172),
    .D(_00361_),
    .Q_N(_00119_),
    .Q(\top_ihp.oisc.regs[0][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1223),
    .D(_00362_),
    .Q_N(_00120_),
    .Q(\top_ihp.oisc.regs[0][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1181),
    .D(_00363_),
    .Q_N(_00121_),
    .Q(\top_ihp.oisc.regs[0][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1170),
    .D(_00364_),
    .Q_N(_00122_),
    .Q(\top_ihp.oisc.regs[0][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1224),
    .D(_00365_),
    .Q_N(_00123_),
    .Q(\top_ihp.oisc.regs[0][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1181),
    .D(_00366_),
    .Q_N(_00124_),
    .Q(\top_ihp.oisc.regs[0][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1182),
    .D(_00367_),
    .Q_N(_00125_),
    .Q(\top_ihp.oisc.regs[0][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1183),
    .D(_00368_),
    .Q_N(_00126_),
    .Q(\top_ihp.oisc.regs[0][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1224),
    .D(_00369_),
    .Q_N(_00108_),
    .Q(\top_ihp.oisc.regs[0][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1235),
    .D(_00370_),
    .Q_N(_00127_),
    .Q(\top_ihp.oisc.regs[0][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1225),
    .D(_00371_),
    .Q_N(_00128_),
    .Q(\top_ihp.oisc.regs[0][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1233),
    .D(_00372_),
    .Q_N(_00129_),
    .Q(\top_ihp.oisc.regs[0][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1236),
    .D(_00373_),
    .Q_N(_00130_),
    .Q(\top_ihp.oisc.regs[0][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1233),
    .D(_00374_),
    .Q_N(_00131_),
    .Q(\top_ihp.oisc.regs[0][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1233),
    .D(_00375_),
    .Q_N(_00132_),
    .Q(\top_ihp.oisc.regs[0][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1225),
    .D(_00376_),
    .Q_N(_00133_),
    .Q(\top_ihp.oisc.regs[0][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1233),
    .D(_00377_),
    .Q_N(_00134_),
    .Q(\top_ihp.oisc.regs[0][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1233),
    .D(_00378_),
    .Q_N(_00135_),
    .Q(\top_ihp.oisc.regs[0][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1225),
    .D(_00379_),
    .Q_N(_00136_),
    .Q(\top_ihp.oisc.regs[0][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1224),
    .D(_00380_),
    .Q_N(_00109_),
    .Q(\top_ihp.oisc.regs[0][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1224),
    .D(_00381_),
    .Q_N(_00137_),
    .Q(\top_ihp.oisc.regs[0][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1183),
    .D(_00382_),
    .Q_N(_00068_),
    .Q(\top_ihp.oisc.regs[0][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1183),
    .D(_00383_),
    .Q_N(_00110_),
    .Q(\top_ihp.oisc.regs[0][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1181),
    .D(_00384_),
    .Q_N(_00111_),
    .Q(\top_ihp.oisc.regs[0][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1181),
    .D(_00385_),
    .Q_N(_00112_),
    .Q(\top_ihp.oisc.regs[0][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1172),
    .D(_00386_),
    .Q_N(_00113_),
    .Q(\top_ihp.oisc.regs[0][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1172),
    .D(_00387_),
    .Q_N(_00114_),
    .Q(\top_ihp.oisc.regs[0][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1172),
    .D(_00388_),
    .Q_N(_00115_),
    .Q(\top_ihp.oisc.regs[0][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1172),
    .D(_00389_),
    .Q_N(_00116_),
    .Q(\top_ihp.oisc.regs[0][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1159),
    .D(_00390_),
    .Q_N(\top_ihp.oisc.regs[10][0] ),
    .Q(_00141_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1121),
    .D(_00391_),
    .Q_N(_13017_),
    .Q(\top_ihp.oisc.regs[10][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1124),
    .D(_00392_),
    .Q_N(_13016_),
    .Q(\top_ihp.oisc.regs[10][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1126),
    .D(_00393_),
    .Q_N(_13015_),
    .Q(\top_ihp.oisc.regs[10][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1235),
    .D(_00394_),
    .Q_N(_13014_),
    .Q(\top_ihp.oisc.regs[10][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1133),
    .D(_00395_),
    .Q_N(_13013_),
    .Q(\top_ihp.oisc.regs[10][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1125),
    .D(_00396_),
    .Q_N(_13012_),
    .Q(\top_ihp.oisc.regs[10][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1235),
    .D(_00397_),
    .Q_N(_13011_),
    .Q(\top_ihp.oisc.regs[10][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1133),
    .D(_00398_),
    .Q_N(_13010_),
    .Q(\top_ihp.oisc.regs[10][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1135),
    .D(_00399_),
    .Q_N(_13009_),
    .Q(\top_ihp.oisc.regs[10][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1130),
    .D(_00400_),
    .Q_N(_13008_),
    .Q(\top_ihp.oisc.regs[10][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1130),
    .D(_00401_),
    .Q_N(_13007_),
    .Q(\top_ihp.oisc.regs[10][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1164),
    .D(_00402_),
    .Q_N(_13006_),
    .Q(\top_ihp.oisc.regs[10][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1155),
    .D(_00403_),
    .Q_N(_13005_),
    .Q(\top_ihp.oisc.regs[10][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1165),
    .D(_00404_),
    .Q_N(_13004_),
    .Q(\top_ihp.oisc.regs[10][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1164),
    .D(_00405_),
    .Q_N(_13003_),
    .Q(\top_ihp.oisc.regs[10][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1159),
    .D(_00406_),
    .Q_N(_13002_),
    .Q(\top_ihp.oisc.regs[10][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1158),
    .D(_00407_),
    .Q_N(_13001_),
    .Q(\top_ihp.oisc.regs[10][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1155),
    .D(_00408_),
    .Q_N(_13000_),
    .Q(\top_ihp.oisc.regs[10][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1165),
    .D(_00409_),
    .Q_N(_12999_),
    .Q(\top_ihp.oisc.regs[10][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1162),
    .D(_00410_),
    .Q_N(_12998_),
    .Q(\top_ihp.oisc.regs[10][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1155),
    .D(_00411_),
    .Q_N(_12997_),
    .Q(\top_ihp.oisc.regs[10][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1149),
    .D(_00412_),
    .Q_N(_12996_),
    .Q(\top_ihp.oisc.regs[10][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1149),
    .D(_00413_),
    .Q_N(_12995_),
    .Q(\top_ihp.oisc.regs[10][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1130),
    .D(_00414_),
    .Q_N(_12994_),
    .Q(\top_ihp.oisc.regs[10][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1130),
    .D(_00415_),
    .Q_N(_12993_),
    .Q(\top_ihp.oisc.regs[10][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1130),
    .D(_00416_),
    .Q_N(_12992_),
    .Q(\top_ihp.oisc.regs[10][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1129),
    .D(_00417_),
    .Q_N(_12991_),
    .Q(\top_ihp.oisc.regs[10][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1119),
    .D(_00418_),
    .Q_N(_12990_),
    .Q(\top_ihp.oisc.regs[10][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1119),
    .D(_00419_),
    .Q_N(_12989_),
    .Q(\top_ihp.oisc.regs[10][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1121),
    .D(_00420_),
    .Q_N(_12988_),
    .Q(\top_ihp.oisc.regs[10][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1121),
    .D(_00421_),
    .Q_N(_12987_),
    .Q(\top_ihp.oisc.regs[10][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1130),
    .D(_00422_),
    .Q_N(\top_ihp.oisc.regs[11][0] ),
    .Q(_00142_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1122),
    .D(_00423_),
    .Q_N(_12986_),
    .Q(\top_ihp.oisc.regs[11][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1126),
    .D(_00424_),
    .Q_N(_12985_),
    .Q(\top_ihp.oisc.regs[11][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1126),
    .D(_00425_),
    .Q_N(_12984_),
    .Q(\top_ihp.oisc.regs[11][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1153),
    .D(_00426_),
    .Q_N(_12983_),
    .Q(\top_ihp.oisc.regs[11][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1133),
    .D(_00427_),
    .Q_N(_12982_),
    .Q(\top_ihp.oisc.regs[11][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1126),
    .D(_00428_),
    .Q_N(_12981_),
    .Q(\top_ihp.oisc.regs[11][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1153),
    .D(_00429_),
    .Q_N(_12980_),
    .Q(\top_ihp.oisc.regs[11][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1180),
    .D(_00430_),
    .Q_N(_12979_),
    .Q(\top_ihp.oisc.regs[11][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1182),
    .D(_00431_),
    .Q_N(_12978_),
    .Q(\top_ihp.oisc.regs[11][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1135),
    .D(_00432_),
    .Q_N(_12977_),
    .Q(\top_ihp.oisc.regs[11][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][1]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1115),
    .D(_00433_),
    .Q_N(\top_ihp.oisc.regs[11][1] ),
    .Q(_00143_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1146),
    .D(_00434_),
    .Q_N(_12976_),
    .Q(\top_ihp.oisc.regs[11][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1155),
    .D(_00435_),
    .Q_N(_12975_),
    .Q(\top_ihp.oisc.regs[11][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1162),
    .D(_00436_),
    .Q_N(_12974_),
    .Q(\top_ihp.oisc.regs[11][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1146),
    .D(_00437_),
    .Q_N(_12973_),
    .Q(\top_ihp.oisc.regs[11][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1158),
    .D(_00438_),
    .Q_N(_12972_),
    .Q(\top_ihp.oisc.regs[11][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1158),
    .D(_00439_),
    .Q_N(_12971_),
    .Q(\top_ihp.oisc.regs[11][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1162),
    .D(_00440_),
    .Q_N(_12970_),
    .Q(\top_ihp.oisc.regs[11][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1163),
    .D(_00441_),
    .Q_N(_12969_),
    .Q(\top_ihp.oisc.regs[11][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1234),
    .D(_00442_),
    .Q_N(_12968_),
    .Q(\top_ihp.oisc.regs[11][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1225),
    .D(_00443_),
    .Q_N(_12967_),
    .Q(\top_ihp.oisc.regs[11][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1140),
    .D(_00444_),
    .Q_N(\top_ihp.oisc.regs[11][2] ),
    .Q(_00144_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1153),
    .D(_00445_),
    .Q_N(_12966_),
    .Q(\top_ihp.oisc.regs[11][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1130),
    .D(_00446_),
    .Q_N(_12965_),
    .Q(\top_ihp.oisc.regs[11][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1115),
    .D(_00447_),
    .Q_N(\top_ihp.oisc.regs[11][3] ),
    .Q(_00145_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1114),
    .D(_00448_),
    .Q_N(\top_ihp.oisc.regs[11][4] ),
    .Q(_00146_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1129),
    .D(_00449_),
    .Q_N(_12964_),
    .Q(\top_ihp.oisc.regs[11][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1119),
    .D(_00450_),
    .Q_N(_12963_),
    .Q(\top_ihp.oisc.regs[11][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1119),
    .D(_00451_),
    .Q_N(_12962_),
    .Q(\top_ihp.oisc.regs[11][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1121),
    .D(_00452_),
    .Q_N(_12961_),
    .Q(\top_ihp.oisc.regs[11][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1121),
    .D(_00453_),
    .Q_N(_12960_),
    .Q(\top_ihp.oisc.regs[11][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1147),
    .D(_00454_),
    .Q_N(\top_ihp.oisc.regs[12][0] ),
    .Q(_00147_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][10]$_DFFE_PN1P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1119),
    .D(_00455_),
    .Q_N(\top_ihp.oisc.regs[12][10] ),
    .Q(_00148_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1124),
    .D(_00456_),
    .Q_N(\top_ihp.oisc.regs[12][11] ),
    .Q(_00149_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][12]$_DFFE_PN1P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1124),
    .D(_00457_),
    .Q_N(\top_ihp.oisc.regs[12][12] ),
    .Q(_00150_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][13]$_DFFE_PN1P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1142),
    .D(_00458_),
    .Q_N(\top_ihp.oisc.regs[12][13] ),
    .Q(_00151_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][14]$_DFFE_PN1P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1133),
    .D(_00459_),
    .Q_N(\top_ihp.oisc.regs[12][14] ),
    .Q(_00152_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1127),
    .D(_00460_),
    .Q_N(\top_ihp.oisc.regs[12][15] ),
    .Q(_00153_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][16]$_DFFE_PN1P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1142),
    .D(_00461_),
    .Q_N(\top_ihp.oisc.regs[12][16] ),
    .Q(_00154_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][17]$_DFFE_PN1P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1114),
    .D(_00462_),
    .Q_N(\top_ihp.oisc.regs[12][17] ),
    .Q(_00155_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][18]$_DFFE_PN1P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1136),
    .D(_00463_),
    .Q_N(\top_ihp.oisc.regs[12][18] ),
    .Q(_00156_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][19]$_DFFE_PN1P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1135),
    .D(_00464_),
    .Q_N(\top_ihp.oisc.regs[12][19] ),
    .Q(_00157_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][1]$_DFFE_PN1P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1153),
    .D(_00465_),
    .Q_N(\top_ihp.oisc.regs[12][1] ),
    .Q(_00158_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][20]$_DFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1146),
    .D(_00466_),
    .Q_N(\top_ihp.oisc.regs[12][20] ),
    .Q(_00159_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][21]$_DFFE_PN1P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1151),
    .D(_00467_),
    .Q_N(\top_ihp.oisc.regs[12][21] ),
    .Q(_00160_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][22]$_DFFE_PN1P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1147),
    .D(_00468_),
    .Q_N(\top_ihp.oisc.regs[12][22] ),
    .Q(_00161_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][23]$_DFFE_PN1P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1146),
    .D(_00469_),
    .Q_N(\top_ihp.oisc.regs[12][23] ),
    .Q(_00162_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][24]$_DFFE_PN1P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1150),
    .D(_00470_),
    .Q_N(\top_ihp.oisc.regs[12][24] ),
    .Q(_00163_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][25]$_DFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1146),
    .D(_00471_),
    .Q_N(\top_ihp.oisc.regs[12][25] ),
    .Q(_00164_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][26]$_DFFE_PN1P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1156),
    .D(_00472_),
    .Q_N(\top_ihp.oisc.regs[12][26] ),
    .Q(_00165_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1147),
    .D(_00473_),
    .Q_N(\top_ihp.oisc.regs[12][27] ),
    .Q(_00166_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][28]$_DFFE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1140),
    .D(_00474_),
    .Q_N(\top_ihp.oisc.regs[12][28] ),
    .Q(_00167_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][29]$_DFFE_PN1P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1140),
    .D(_00475_),
    .Q_N(\top_ihp.oisc.regs[12][29] ),
    .Q(_00168_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1142),
    .D(_00476_),
    .Q_N(\top_ihp.oisc.regs[12][2] ),
    .Q(_00169_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1142),
    .D(_00477_),
    .Q_N(\top_ihp.oisc.regs[12][30] ),
    .Q(_00170_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1115),
    .D(_00478_),
    .Q_N(\top_ihp.oisc.regs[12][31] ),
    .Q(_00171_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1115),
    .D(_00479_),
    .Q_N(\top_ihp.oisc.regs[12][3] ),
    .Q(_00172_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1114),
    .D(_00480_),
    .Q_N(\top_ihp.oisc.regs[12][4] ),
    .Q(_00173_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][5]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1114),
    .D(_00481_),
    .Q_N(\top_ihp.oisc.regs[12][5] ),
    .Q(_00174_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][6]$_DFFE_PN1P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1109),
    .D(_00482_),
    .Q_N(\top_ihp.oisc.regs[12][6] ),
    .Q(_00175_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][7]$_DFFE_PN1P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1109),
    .D(_00483_),
    .Q_N(\top_ihp.oisc.regs[12][7] ),
    .Q(_00176_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][8]$_DFFE_PN1P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1114),
    .D(_00484_),
    .Q_N(\top_ihp.oisc.regs[12][8] ),
    .Q(_00177_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][9]$_DFFE_PN1P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1109),
    .D(_00485_),
    .Q_N(\top_ihp.oisc.regs[12][9] ),
    .Q(_00178_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1147),
    .D(_00486_),
    .Q_N(_12959_),
    .Q(\top_ihp.oisc.regs[13][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][10]$_DFFE_PN1P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1108),
    .D(_00487_),
    .Q_N(\top_ihp.oisc.regs[13][10] ),
    .Q(_00179_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1109),
    .D(_00488_),
    .Q_N(\top_ihp.oisc.regs[13][11] ),
    .Q(_00180_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][12]$_DFFE_PN1P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1109),
    .D(_00489_),
    .Q_N(\top_ihp.oisc.regs[13][12] ),
    .Q(_00181_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][13]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1140),
    .D(_00490_),
    .Q_N(\top_ihp.oisc.regs[13][13] ),
    .Q(_00182_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][14]$_DFFE_PN1P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1133),
    .D(_00491_),
    .Q_N(\top_ihp.oisc.regs[13][14] ),
    .Q(_00183_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1171),
    .D(_00492_),
    .Q_N(\top_ihp.oisc.regs[13][15] ),
    .Q(_00184_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][16]$_DFFE_PN1P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1225),
    .D(_00493_),
    .Q_N(\top_ihp.oisc.regs[13][16] ),
    .Q(_00185_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][17]$_DFFE_PN1P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1180),
    .D(_00494_),
    .Q_N(\top_ihp.oisc.regs[13][17] ),
    .Q(_00186_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][18]$_DFFE_PN1P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1180),
    .D(_00495_),
    .Q_N(\top_ihp.oisc.regs[13][18] ),
    .Q(_00187_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][19]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1115),
    .D(_00496_),
    .Q_N(\top_ihp.oisc.regs[13][19] ),
    .Q(_00188_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1115),
    .D(_00497_),
    .Q_N(_12958_),
    .Q(\top_ihp.oisc.regs[13][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][20]$_DFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1150),
    .D(_00498_),
    .Q_N(\top_ihp.oisc.regs[13][20] ),
    .Q(_00189_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][21]$_DFFE_PN1P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1155),
    .D(_00499_),
    .Q_N(\top_ihp.oisc.regs[13][21] ),
    .Q(_00190_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][22]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1147),
    .D(_00500_),
    .Q_N(\top_ihp.oisc.regs[13][22] ),
    .Q(_00191_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][23]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1147),
    .D(_00501_),
    .Q_N(\top_ihp.oisc.regs[13][23] ),
    .Q(_00192_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][24]$_DFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1145),
    .D(_00502_),
    .Q_N(\top_ihp.oisc.regs[13][24] ),
    .Q(_00193_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][25]$_DFFE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1147),
    .D(_00503_),
    .Q_N(\top_ihp.oisc.regs[13][25] ),
    .Q(_00194_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][26]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1140),
    .D(_00504_),
    .Q_N(\top_ihp.oisc.regs[13][26] ),
    .Q(_00195_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1146),
    .D(_00505_),
    .Q_N(\top_ihp.oisc.regs[13][27] ),
    .Q(_00196_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][28]$_DFFE_PN1P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1147),
    .D(_00506_),
    .Q_N(\top_ihp.oisc.regs[13][28] ),
    .Q(_00197_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][29]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1140),
    .D(_00507_),
    .Q_N(\top_ihp.oisc.regs[13][29] ),
    .Q(_00198_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1142),
    .D(_00508_),
    .Q_N(\top_ihp.oisc.regs[13][2] ),
    .Q(_00199_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1142),
    .D(_00509_),
    .Q_N(\top_ihp.oisc.regs[13][30] ),
    .Q(_00200_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1112),
    .D(_00510_),
    .Q_N(\top_ihp.oisc.regs[13][31] ),
    .Q(_00201_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1115),
    .D(_00511_),
    .Q_N(\top_ihp.oisc.regs[13][3] ),
    .Q(_00202_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1118),
    .D(_00512_),
    .Q_N(\top_ihp.oisc.regs[13][4] ),
    .Q(_00203_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][5]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1114),
    .D(_00513_),
    .Q_N(\top_ihp.oisc.regs[13][5] ),
    .Q(_00204_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][6]$_DFFE_PN1P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1109),
    .D(_00514_),
    .Q_N(\top_ihp.oisc.regs[13][6] ),
    .Q(_00205_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][7]$_DFFE_PN1P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1109),
    .D(_00515_),
    .Q_N(\top_ihp.oisc.regs[13][7] ),
    .Q(_00206_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][8]$_DFFE_PN1P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1109),
    .D(_00516_),
    .Q_N(\top_ihp.oisc.regs[13][8] ),
    .Q(_00207_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][9]$_DFFE_PN1P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1108),
    .D(_00517_),
    .Q_N(\top_ihp.oisc.regs[13][9] ),
    .Q(_00208_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1159),
    .D(_00518_),
    .Q_N(_12957_),
    .Q(\top_ihp.oisc.regs[14][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1122),
    .D(_00519_),
    .Q_N(_12956_),
    .Q(\top_ihp.oisc.regs[14][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1126),
    .D(_00520_),
    .Q_N(_12955_),
    .Q(\top_ihp.oisc.regs[14][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1127),
    .D(_00521_),
    .Q_N(_12954_),
    .Q(\top_ihp.oisc.regs[14][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1239),
    .D(_00522_),
    .Q_N(_12953_),
    .Q(\top_ihp.oisc.regs[14][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1133),
    .D(_00523_),
    .Q_N(_12952_),
    .Q(\top_ihp.oisc.regs[14][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1127),
    .D(_00524_),
    .Q_N(_12951_),
    .Q(\top_ihp.oisc.regs[14][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1239),
    .D(_00525_),
    .Q_N(_12950_),
    .Q(\top_ihp.oisc.regs[14][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1180),
    .D(_00526_),
    .Q_N(_12949_),
    .Q(\top_ihp.oisc.regs[14][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1136),
    .D(_00527_),
    .Q_N(_12948_),
    .Q(\top_ihp.oisc.regs[14][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1135),
    .D(_00528_),
    .Q_N(_12947_),
    .Q(\top_ihp.oisc.regs[14][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1135),
    .D(_00529_),
    .Q_N(_12946_),
    .Q(\top_ihp.oisc.regs[14][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1160),
    .D(_00530_),
    .Q_N(_12945_),
    .Q(\top_ihp.oisc.regs[14][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1156),
    .D(_00531_),
    .Q_N(_12944_),
    .Q(\top_ihp.oisc.regs[14][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1239),
    .D(_00532_),
    .Q_N(_12943_),
    .Q(\top_ihp.oisc.regs[14][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1241),
    .D(_00533_),
    .Q_N(_12942_),
    .Q(\top_ihp.oisc.regs[14][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1151),
    .D(_00534_),
    .Q_N(_12941_),
    .Q(\top_ihp.oisc.regs[14][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1162),
    .D(_00535_),
    .Q_N(_12940_),
    .Q(\top_ihp.oisc.regs[14][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1156),
    .D(_00536_),
    .Q_N(_12939_),
    .Q(\top_ihp.oisc.regs[14][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1163),
    .D(_00537_),
    .Q_N(_12938_),
    .Q(\top_ihp.oisc.regs[14][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1234),
    .D(_00538_),
    .Q_N(_12937_),
    .Q(\top_ihp.oisc.regs[14][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1225),
    .D(_00539_),
    .Q_N(_12936_),
    .Q(\top_ihp.oisc.regs[14][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1149),
    .D(_00540_),
    .Q_N(_12935_),
    .Q(\top_ihp.oisc.regs[14][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1154),
    .D(_00541_),
    .Q_N(_12934_),
    .Q(\top_ihp.oisc.regs[14][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1182),
    .D(_00542_),
    .Q_N(_12933_),
    .Q(\top_ihp.oisc.regs[14][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1135),
    .D(_00543_),
    .Q_N(_12932_),
    .Q(\top_ihp.oisc.regs[14][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1129),
    .D(_00544_),
    .Q_N(_12931_),
    .Q(\top_ihp.oisc.regs[14][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1129),
    .D(_00545_),
    .Q_N(_12930_),
    .Q(\top_ihp.oisc.regs[14][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1121),
    .D(_00546_),
    .Q_N(_12929_),
    .Q(\top_ihp.oisc.regs[14][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1121),
    .D(_00547_),
    .Q_N(_12928_),
    .Q(\top_ihp.oisc.regs[14][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1122),
    .D(_00548_),
    .Q_N(_12927_),
    .Q(\top_ihp.oisc.regs[14][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1122),
    .D(_00549_),
    .Q_N(_12926_),
    .Q(\top_ihp.oisc.regs[14][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1160),
    .D(_00550_),
    .Q_N(_12925_),
    .Q(\top_ihp.oisc.regs[15][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1124),
    .D(_00551_),
    .Q_N(_12924_),
    .Q(\top_ihp.oisc.regs[15][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1124),
    .D(_00552_),
    .Q_N(_12923_),
    .Q(\top_ihp.oisc.regs[15][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1171),
    .D(_00553_),
    .Q_N(_12922_),
    .Q(\top_ihp.oisc.regs[15][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1223),
    .D(_00554_),
    .Q_N(_12921_),
    .Q(\top_ihp.oisc.regs[15][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1124),
    .D(_00555_),
    .Q_N(_12920_),
    .Q(\top_ihp.oisc.regs[15][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1125),
    .D(_00556_),
    .Q_N(_12919_),
    .Q(\top_ihp.oisc.regs[15][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1223),
    .D(_00557_),
    .Q_N(_12918_),
    .Q(\top_ihp.oisc.regs[15][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1133),
    .D(_00558_),
    .Q_N(_12917_),
    .Q(\top_ihp.oisc.regs[15][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1136),
    .D(_00559_),
    .Q_N(_12916_),
    .Q(\top_ihp.oisc.regs[15][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1135),
    .D(_00560_),
    .Q_N(_12915_),
    .Q(\top_ihp.oisc.regs[15][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1149),
    .D(_00561_),
    .Q_N(_12914_),
    .Q(\top_ihp.oisc.regs[15][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1150),
    .D(_00562_),
    .Q_N(_12913_),
    .Q(\top_ihp.oisc.regs[15][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1153),
    .D(_00563_),
    .Q_N(_12912_),
    .Q(\top_ihp.oisc.regs[15][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1163),
    .D(_00564_),
    .Q_N(_12911_),
    .Q(\top_ihp.oisc.regs[15][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1160),
    .D(_00565_),
    .Q_N(_12910_),
    .Q(\top_ihp.oisc.regs[15][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1158),
    .D(_00566_),
    .Q_N(_12909_),
    .Q(\top_ihp.oisc.regs[15][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1158),
    .D(_00567_),
    .Q_N(_12908_),
    .Q(\top_ihp.oisc.regs[15][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1155),
    .D(_00568_),
    .Q_N(_12907_),
    .Q(\top_ihp.oisc.regs[15][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1163),
    .D(_00569_),
    .Q_N(_12906_),
    .Q(\top_ihp.oisc.regs[15][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1162),
    .D(_00570_),
    .Q_N(_12905_),
    .Q(\top_ihp.oisc.regs[15][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1156),
    .D(_00571_),
    .Q_N(_12904_),
    .Q(\top_ihp.oisc.regs[15][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1149),
    .D(_00572_),
    .Q_N(_12903_),
    .Q(\top_ihp.oisc.regs[15][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1149),
    .D(_00573_),
    .Q_N(_12902_),
    .Q(\top_ihp.oisc.regs[15][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1130),
    .D(_00574_),
    .Q_N(_12901_),
    .Q(\top_ihp.oisc.regs[15][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1131),
    .D(_00575_),
    .Q_N(_12900_),
    .Q(\top_ihp.oisc.regs[15][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1117),
    .D(_00576_),
    .Q_N(_12899_),
    .Q(\top_ihp.oisc.regs[15][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1129),
    .D(_00577_),
    .Q_N(_12898_),
    .Q(\top_ihp.oisc.regs[15][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1110),
    .D(_00578_),
    .Q_N(_12897_),
    .Q(\top_ihp.oisc.regs[15][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1121),
    .D(_00579_),
    .Q_N(_12896_),
    .Q(\top_ihp.oisc.regs[15][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1129),
    .D(_00580_),
    .Q_N(_12895_),
    .Q(\top_ihp.oisc.regs[15][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1122),
    .D(_00581_),
    .Q_N(_12894_),
    .Q(\top_ihp.oisc.regs[15][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1413),
    .D(_00582_),
    .Q_N(_12893_),
    .Q(\top_ihp.oisc.regs[16][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1414),
    .D(_00583_),
    .Q_N(_12892_),
    .Q(\top_ihp.oisc.regs[16][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1415),
    .D(_00584_),
    .Q_N(_12891_),
    .Q(\top_ihp.oisc.regs[16][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1416),
    .D(_00585_),
    .Q_N(_12890_),
    .Q(\top_ihp.oisc.regs[16][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1417),
    .D(_00586_),
    .Q_N(_12889_),
    .Q(\top_ihp.oisc.regs[16][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1418),
    .D(_00587_),
    .Q_N(_12888_),
    .Q(\top_ihp.oisc.regs[16][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1419),
    .D(_00588_),
    .Q_N(_12887_),
    .Q(\top_ihp.oisc.regs[16][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1420),
    .D(_00589_),
    .Q_N(_12886_),
    .Q(\top_ihp.oisc.regs[16][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1421),
    .D(_00590_),
    .Q_N(_12885_),
    .Q(\top_ihp.oisc.regs[16][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1422),
    .D(_00591_),
    .Q_N(_12884_),
    .Q(\top_ihp.oisc.regs[16][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1423),
    .D(_00592_),
    .Q_N(_12883_),
    .Q(\top_ihp.oisc.regs[16][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1424),
    .D(_00593_),
    .Q_N(_12882_),
    .Q(\top_ihp.oisc.regs[16][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1425),
    .D(_00594_),
    .Q_N(_12881_),
    .Q(\top_ihp.oisc.regs[16][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1426),
    .D(_00595_),
    .Q_N(_12880_),
    .Q(\top_ihp.oisc.regs[16][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1427),
    .D(_00596_),
    .Q_N(_12879_),
    .Q(\top_ihp.oisc.regs[16][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1428),
    .D(_00597_),
    .Q_N(_12878_),
    .Q(\top_ihp.oisc.regs[16][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1429),
    .D(_00598_),
    .Q_N(_12877_),
    .Q(\top_ihp.oisc.regs[16][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1430),
    .D(_00599_),
    .Q_N(_12876_),
    .Q(\top_ihp.oisc.regs[16][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1431),
    .D(_00600_),
    .Q_N(_12875_),
    .Q(\top_ihp.oisc.regs[16][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1432),
    .D(_00601_),
    .Q_N(_12874_),
    .Q(\top_ihp.oisc.regs[16][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1433),
    .D(_00602_),
    .Q_N(_12873_),
    .Q(\top_ihp.oisc.regs[16][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1434),
    .D(_00603_),
    .Q_N(_12872_),
    .Q(\top_ihp.oisc.regs[16][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1435),
    .D(_00604_),
    .Q_N(_12871_),
    .Q(\top_ihp.oisc.regs[16][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1436),
    .D(_00605_),
    .Q_N(_12870_),
    .Q(\top_ihp.oisc.regs[16][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1437),
    .D(_00606_),
    .Q_N(_12869_),
    .Q(\top_ihp.oisc.regs[16][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1438),
    .D(_00607_),
    .Q_N(_12868_),
    .Q(\top_ihp.oisc.regs[16][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1439),
    .D(_00608_),
    .Q_N(_12867_),
    .Q(\top_ihp.oisc.regs[16][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1440),
    .D(_00609_),
    .Q_N(_12866_),
    .Q(\top_ihp.oisc.regs[16][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1441),
    .D(_00610_),
    .Q_N(_12865_),
    .Q(\top_ihp.oisc.regs[16][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1442),
    .D(_00611_),
    .Q_N(_12864_),
    .Q(\top_ihp.oisc.regs[16][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1443),
    .D(_00612_),
    .Q_N(_12863_),
    .Q(\top_ihp.oisc.regs[16][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1444),
    .D(_00613_),
    .Q_N(_12862_),
    .Q(\top_ihp.oisc.regs[16][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1445),
    .D(_00614_),
    .Q_N(_12861_),
    .Q(\top_ihp.oisc.regs[17][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1446),
    .D(_00615_),
    .Q_N(_12860_),
    .Q(\top_ihp.oisc.regs[17][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1447),
    .D(_00616_),
    .Q_N(_12859_),
    .Q(\top_ihp.oisc.regs[17][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1448),
    .D(_00617_),
    .Q_N(_12858_),
    .Q(\top_ihp.oisc.regs[17][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1449),
    .D(_00618_),
    .Q_N(_12857_),
    .Q(\top_ihp.oisc.regs[17][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][14]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1450),
    .D(_00619_),
    .Q_N(_12856_),
    .Q(\top_ihp.oisc.regs[17][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1451),
    .D(_00620_),
    .Q_N(_12855_),
    .Q(\top_ihp.oisc.regs[17][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1452),
    .D(_00621_),
    .Q_N(_12854_),
    .Q(\top_ihp.oisc.regs[17][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1453),
    .D(_00622_),
    .Q_N(_12853_),
    .Q(\top_ihp.oisc.regs[17][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1454),
    .D(_00623_),
    .Q_N(_12852_),
    .Q(\top_ihp.oisc.regs[17][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1455),
    .D(_00624_),
    .Q_N(_12851_),
    .Q(\top_ihp.oisc.regs[17][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1456),
    .D(_00625_),
    .Q_N(_12850_),
    .Q(\top_ihp.oisc.regs[17][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1457),
    .D(_00626_),
    .Q_N(_12849_),
    .Q(\top_ihp.oisc.regs[17][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1458),
    .D(_00627_),
    .Q_N(_12848_),
    .Q(\top_ihp.oisc.regs[17][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1459),
    .D(_00628_),
    .Q_N(_12847_),
    .Q(\top_ihp.oisc.regs[17][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1460),
    .D(_00629_),
    .Q_N(_12846_),
    .Q(\top_ihp.oisc.regs[17][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1461),
    .D(_00630_),
    .Q_N(_12845_),
    .Q(\top_ihp.oisc.regs[17][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][25]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1462),
    .D(_00631_),
    .Q_N(_12844_),
    .Q(\top_ihp.oisc.regs[17][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1463),
    .D(_00632_),
    .Q_N(_12843_),
    .Q(\top_ihp.oisc.regs[17][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1464),
    .D(_00633_),
    .Q_N(_12842_),
    .Q(\top_ihp.oisc.regs[17][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1465),
    .D(_00634_),
    .Q_N(_12841_),
    .Q(\top_ihp.oisc.regs[17][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1466),
    .D(_00635_),
    .Q_N(_12840_),
    .Q(\top_ihp.oisc.regs[17][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1467),
    .D(_00636_),
    .Q_N(_12839_),
    .Q(\top_ihp.oisc.regs[17][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1468),
    .D(_00637_),
    .Q_N(_12838_),
    .Q(\top_ihp.oisc.regs[17][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1469),
    .D(_00638_),
    .Q_N(_12837_),
    .Q(\top_ihp.oisc.regs[17][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1470),
    .D(_00639_),
    .Q_N(_12836_),
    .Q(\top_ihp.oisc.regs[17][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1471),
    .D(_00640_),
    .Q_N(_12835_),
    .Q(\top_ihp.oisc.regs[17][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1472),
    .D(_00641_),
    .Q_N(_12834_),
    .Q(\top_ihp.oisc.regs[17][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1473),
    .D(_00642_),
    .Q_N(_12833_),
    .Q(\top_ihp.oisc.regs[17][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1474),
    .D(_00643_),
    .Q_N(_12832_),
    .Q(\top_ihp.oisc.regs[17][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1475),
    .D(_00644_),
    .Q_N(_12831_),
    .Q(\top_ihp.oisc.regs[17][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1476),
    .D(_00645_),
    .Q_N(_12830_),
    .Q(\top_ihp.oisc.regs[17][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1477),
    .D(_00646_),
    .Q_N(_12829_),
    .Q(\top_ihp.oisc.regs[18][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1478),
    .D(_00647_),
    .Q_N(_12828_),
    .Q(\top_ihp.oisc.regs[18][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1479),
    .D(_00648_),
    .Q_N(_12827_),
    .Q(\top_ihp.oisc.regs[18][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][12]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1480),
    .D(_00649_),
    .Q_N(_12826_),
    .Q(\top_ihp.oisc.regs[18][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1481),
    .D(_00650_),
    .Q_N(_12825_),
    .Q(\top_ihp.oisc.regs[18][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1482),
    .D(_00651_),
    .Q_N(_12824_),
    .Q(\top_ihp.oisc.regs[18][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1483),
    .D(_00652_),
    .Q_N(_12823_),
    .Q(\top_ihp.oisc.regs[18][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1484),
    .D(_00653_),
    .Q_N(_12822_),
    .Q(\top_ihp.oisc.regs[18][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1485),
    .D(_00654_),
    .Q_N(_12821_),
    .Q(\top_ihp.oisc.regs[18][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1486),
    .D(_00655_),
    .Q_N(_12820_),
    .Q(\top_ihp.oisc.regs[18][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][19]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1487),
    .D(_00656_),
    .Q_N(_12819_),
    .Q(\top_ihp.oisc.regs[18][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1488),
    .D(_00657_),
    .Q_N(_12818_),
    .Q(\top_ihp.oisc.regs[18][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][20]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1489),
    .D(_00658_),
    .Q_N(_12817_),
    .Q(\top_ihp.oisc.regs[18][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1490),
    .D(_00659_),
    .Q_N(_12816_),
    .Q(\top_ihp.oisc.regs[18][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1491),
    .D(_00660_),
    .Q_N(_12815_),
    .Q(\top_ihp.oisc.regs[18][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1492),
    .D(_00661_),
    .Q_N(_12814_),
    .Q(\top_ihp.oisc.regs[18][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1493),
    .D(_00662_),
    .Q_N(_12813_),
    .Q(\top_ihp.oisc.regs[18][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1494),
    .D(_00663_),
    .Q_N(_12812_),
    .Q(\top_ihp.oisc.regs[18][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1495),
    .D(_00664_),
    .Q_N(_12811_),
    .Q(\top_ihp.oisc.regs[18][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1496),
    .D(_00665_),
    .Q_N(_12810_),
    .Q(\top_ihp.oisc.regs[18][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][28]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1497),
    .D(_00666_),
    .Q_N(_12809_),
    .Q(\top_ihp.oisc.regs[18][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1498),
    .D(_00667_),
    .Q_N(_12808_),
    .Q(\top_ihp.oisc.regs[18][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1499),
    .D(_00668_),
    .Q_N(_12807_),
    .Q(\top_ihp.oisc.regs[18][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1500),
    .D(_00669_),
    .Q_N(_12806_),
    .Q(\top_ihp.oisc.regs[18][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1501),
    .D(_00670_),
    .Q_N(_12805_),
    .Q(\top_ihp.oisc.regs[18][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1502),
    .D(_00671_),
    .Q_N(_12804_),
    .Q(\top_ihp.oisc.regs[18][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1503),
    .D(_00672_),
    .Q_N(_12803_),
    .Q(\top_ihp.oisc.regs[18][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1504),
    .D(_00673_),
    .Q_N(_12802_),
    .Q(\top_ihp.oisc.regs[18][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1505),
    .D(_00674_),
    .Q_N(_12801_),
    .Q(\top_ihp.oisc.regs[18][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1506),
    .D(_00675_),
    .Q_N(_12800_),
    .Q(\top_ihp.oisc.regs[18][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1507),
    .D(_00676_),
    .Q_N(_12799_),
    .Q(\top_ihp.oisc.regs[18][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1508),
    .D(_00677_),
    .Q_N(_12798_),
    .Q(\top_ihp.oisc.regs[18][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1509),
    .D(_00678_),
    .Q_N(_12797_),
    .Q(\top_ihp.oisc.regs[19][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1510),
    .D(_00679_),
    .Q_N(_12796_),
    .Q(\top_ihp.oisc.regs[19][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1511),
    .D(_00680_),
    .Q_N(_12795_),
    .Q(\top_ihp.oisc.regs[19][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1512),
    .D(_00681_),
    .Q_N(_12794_),
    .Q(\top_ihp.oisc.regs[19][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1513),
    .D(_00682_),
    .Q_N(_12793_),
    .Q(\top_ihp.oisc.regs[19][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1514),
    .D(_00683_),
    .Q_N(_12792_),
    .Q(\top_ihp.oisc.regs[19][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1515),
    .D(_00684_),
    .Q_N(_12791_),
    .Q(\top_ihp.oisc.regs[19][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][16]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1516),
    .D(_00685_),
    .Q_N(_12790_),
    .Q(\top_ihp.oisc.regs[19][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1517),
    .D(_00686_),
    .Q_N(_12789_),
    .Q(\top_ihp.oisc.regs[19][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1518),
    .D(_00687_),
    .Q_N(_12788_),
    .Q(\top_ihp.oisc.regs[19][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1519),
    .D(_00688_),
    .Q_N(_12787_),
    .Q(\top_ihp.oisc.regs[19][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1520),
    .D(_00689_),
    .Q_N(_12786_),
    .Q(\top_ihp.oisc.regs[19][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1521),
    .D(_00690_),
    .Q_N(_12785_),
    .Q(\top_ihp.oisc.regs[19][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1522),
    .D(_00691_),
    .Q_N(_12784_),
    .Q(\top_ihp.oisc.regs[19][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][22]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1523),
    .D(_00692_),
    .Q_N(_12783_),
    .Q(\top_ihp.oisc.regs[19][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1524),
    .D(_00693_),
    .Q_N(_12782_),
    .Q(\top_ihp.oisc.regs[19][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][24]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1525),
    .D(_00694_),
    .Q_N(_12781_),
    .Q(\top_ihp.oisc.regs[19][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1526),
    .D(_00695_),
    .Q_N(_12780_),
    .Q(\top_ihp.oisc.regs[19][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1527),
    .D(_00696_),
    .Q_N(_12779_),
    .Q(\top_ihp.oisc.regs[19][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1528),
    .D(_00697_),
    .Q_N(_12778_),
    .Q(\top_ihp.oisc.regs[19][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1529),
    .D(_00698_),
    .Q_N(_12777_),
    .Q(\top_ihp.oisc.regs[19][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1530),
    .D(_00699_),
    .Q_N(_12776_),
    .Q(\top_ihp.oisc.regs[19][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1531),
    .D(_00700_),
    .Q_N(_12775_),
    .Q(\top_ihp.oisc.regs[19][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1532),
    .D(_00701_),
    .Q_N(_12774_),
    .Q(\top_ihp.oisc.regs[19][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1533),
    .D(_00702_),
    .Q_N(_12773_),
    .Q(\top_ihp.oisc.regs[19][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1534),
    .D(_00703_),
    .Q_N(_12772_),
    .Q(\top_ihp.oisc.regs[19][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1535),
    .D(_00704_),
    .Q_N(_12771_),
    .Q(\top_ihp.oisc.regs[19][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1536),
    .D(_00705_),
    .Q_N(_12770_),
    .Q(\top_ihp.oisc.regs[19][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1537),
    .D(_00706_),
    .Q_N(_12769_),
    .Q(\top_ihp.oisc.regs[19][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1538),
    .D(_00707_),
    .Q_N(_12768_),
    .Q(\top_ihp.oisc.regs[19][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1539),
    .D(_00708_),
    .Q_N(_12767_),
    .Q(\top_ihp.oisc.regs[19][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1540),
    .D(_00709_),
    .Q_N(_12766_),
    .Q(\top_ihp.oisc.regs[19][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1161),
    .D(_00710_),
    .Q_N(_12765_),
    .Q(\top_ihp.oisc.regs[1][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1170),
    .D(_00711_),
    .Q_N(_12764_),
    .Q(\top_ihp.oisc.regs[1][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1124),
    .D(_00712_),
    .Q_N(_12763_),
    .Q(\top_ihp.oisc.regs[1][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1170),
    .D(_00713_),
    .Q_N(_12762_),
    .Q(\top_ihp.oisc.regs[1][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1223),
    .D(_00714_),
    .Q_N(_12761_),
    .Q(\top_ihp.oisc.regs[1][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1125),
    .D(_00715_),
    .Q_N(_12760_),
    .Q(\top_ihp.oisc.regs[1][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1170),
    .D(_00716_),
    .Q_N(_12759_),
    .Q(\top_ihp.oisc.regs[1][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1223),
    .D(_00717_),
    .Q_N(_12758_),
    .Q(\top_ihp.oisc.regs[1][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1134),
    .D(_00718_),
    .Q_N(_12757_),
    .Q(\top_ihp.oisc.regs[1][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1182),
    .D(_00719_),
    .Q_N(_12756_),
    .Q(\top_ihp.oisc.regs[1][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1136),
    .D(_00720_),
    .Q_N(_12755_),
    .Q(\top_ihp.oisc.regs[1][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1153),
    .D(_00721_),
    .Q_N(_12754_),
    .Q(\top_ihp.oisc.regs[1][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1162),
    .D(_00722_),
    .Q_N(_12753_),
    .Q(\top_ihp.oisc.regs[1][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1225),
    .D(_00723_),
    .Q_N(_12752_),
    .Q(\top_ihp.oisc.regs[1][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1234),
    .D(_00724_),
    .Q_N(_12751_),
    .Q(\top_ihp.oisc.regs[1][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1162),
    .D(_00725_),
    .Q_N(_12750_),
    .Q(\top_ihp.oisc.regs[1][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1151),
    .D(_00726_),
    .Q_N(_12749_),
    .Q(\top_ihp.oisc.regs[1][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1161),
    .D(_00727_),
    .Q_N(_12748_),
    .Q(\top_ihp.oisc.regs[1][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1155),
    .D(_00728_),
    .Q_N(_12747_),
    .Q(\top_ihp.oisc.regs[1][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1234),
    .D(_00729_),
    .Q_N(_12746_),
    .Q(\top_ihp.oisc.regs[1][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1234),
    .D(_00730_),
    .Q_N(_12745_),
    .Q(\top_ihp.oisc.regs[1][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1225),
    .D(_00731_),
    .Q_N(_12744_),
    .Q(\top_ihp.oisc.regs[1][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1152),
    .D(_00732_),
    .Q_N(_12743_),
    .Q(\top_ihp.oisc.regs[1][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1153),
    .D(_00733_),
    .Q_N(\top_ihp.oisc.regs[1][30] ),
    .Q(_00209_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1182),
    .D(_00734_),
    .Q_N(_12742_),
    .Q(\top_ihp.oisc.regs[1][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1131),
    .D(_00735_),
    .Q_N(_12741_),
    .Q(\top_ihp.oisc.regs[1][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1129),
    .D(_00736_),
    .Q_N(_12740_),
    .Q(\top_ihp.oisc.regs[1][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1132),
    .D(_00737_),
    .Q_N(_12739_),
    .Q(\top_ihp.oisc.regs[1][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1119),
    .D(_00738_),
    .Q_N(_12738_),
    .Q(\top_ihp.oisc.regs[1][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1120),
    .D(_00739_),
    .Q_N(_12737_),
    .Q(\top_ihp.oisc.regs[1][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1122),
    .D(_00740_),
    .Q_N(_12736_),
    .Q(\top_ihp.oisc.regs[1][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1126),
    .D(_00741_),
    .Q_N(_12735_),
    .Q(\top_ihp.oisc.regs[1][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1541),
    .D(_00742_),
    .Q_N(_12734_),
    .Q(\top_ihp.oisc.regs[20][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1542),
    .D(_00743_),
    .Q_N(_12733_),
    .Q(\top_ihp.oisc.regs[20][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1543),
    .D(_00744_),
    .Q_N(_12732_),
    .Q(\top_ihp.oisc.regs[20][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1544),
    .D(_00745_),
    .Q_N(_12731_),
    .Q(\top_ihp.oisc.regs[20][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1545),
    .D(_00746_),
    .Q_N(_12730_),
    .Q(\top_ihp.oisc.regs[20][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1546),
    .D(_00747_),
    .Q_N(_12729_),
    .Q(\top_ihp.oisc.regs[20][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][15]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1547),
    .D(_00748_),
    .Q_N(_12728_),
    .Q(\top_ihp.oisc.regs[20][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1548),
    .D(_00749_),
    .Q_N(_12727_),
    .Q(\top_ihp.oisc.regs[20][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1549),
    .D(_00750_),
    .Q_N(_12726_),
    .Q(\top_ihp.oisc.regs[20][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1550),
    .D(_00751_),
    .Q_N(_12725_),
    .Q(\top_ihp.oisc.regs[20][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1551),
    .D(_00752_),
    .Q_N(_12724_),
    .Q(\top_ihp.oisc.regs[20][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1552),
    .D(_00753_),
    .Q_N(_12723_),
    .Q(\top_ihp.oisc.regs[20][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1553),
    .D(_00754_),
    .Q_N(_12722_),
    .Q(\top_ihp.oisc.regs[20][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][21]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1554),
    .D(_00755_),
    .Q_N(_12721_),
    .Q(\top_ihp.oisc.regs[20][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1555),
    .D(_00756_),
    .Q_N(_12720_),
    .Q(\top_ihp.oisc.regs[20][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1556),
    .D(_00757_),
    .Q_N(_12719_),
    .Q(\top_ihp.oisc.regs[20][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1557),
    .D(_00758_),
    .Q_N(_12718_),
    .Q(\top_ihp.oisc.regs[20][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1558),
    .D(_00759_),
    .Q_N(_12717_),
    .Q(\top_ihp.oisc.regs[20][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1559),
    .D(_00760_),
    .Q_N(_12716_),
    .Q(\top_ihp.oisc.regs[20][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1560),
    .D(_00761_),
    .Q_N(_12715_),
    .Q(\top_ihp.oisc.regs[20][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][28]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1561),
    .D(_00762_),
    .Q_N(_12714_),
    .Q(\top_ihp.oisc.regs[20][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1562),
    .D(_00763_),
    .Q_N(_12713_),
    .Q(\top_ihp.oisc.regs[20][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1563),
    .D(_00764_),
    .Q_N(_12712_),
    .Q(\top_ihp.oisc.regs[20][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1564),
    .D(_00765_),
    .Q_N(_12711_),
    .Q(\top_ihp.oisc.regs[20][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1565),
    .D(_00766_),
    .Q_N(_12710_),
    .Q(\top_ihp.oisc.regs[20][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1566),
    .D(_00767_),
    .Q_N(_12709_),
    .Q(\top_ihp.oisc.regs[20][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1567),
    .D(_00768_),
    .Q_N(_12708_),
    .Q(\top_ihp.oisc.regs[20][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1568),
    .D(_00769_),
    .Q_N(_12707_),
    .Q(\top_ihp.oisc.regs[20][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1569),
    .D(_00770_),
    .Q_N(_12706_),
    .Q(\top_ihp.oisc.regs[20][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1570),
    .D(_00771_),
    .Q_N(_12705_),
    .Q(\top_ihp.oisc.regs[20][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1571),
    .D(_00772_),
    .Q_N(_12704_),
    .Q(\top_ihp.oisc.regs[20][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1572),
    .D(_00773_),
    .Q_N(_12703_),
    .Q(\top_ihp.oisc.regs[20][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1573),
    .D(_00774_),
    .Q_N(_12702_),
    .Q(\top_ihp.oisc.regs[21][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1574),
    .D(_00775_),
    .Q_N(_12701_),
    .Q(\top_ihp.oisc.regs[21][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1575),
    .D(_00776_),
    .Q_N(_12700_),
    .Q(\top_ihp.oisc.regs[21][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1576),
    .D(_00777_),
    .Q_N(_12699_),
    .Q(\top_ihp.oisc.regs[21][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1577),
    .D(_00778_),
    .Q_N(_12698_),
    .Q(\top_ihp.oisc.regs[21][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1578),
    .D(_00779_),
    .Q_N(_12697_),
    .Q(\top_ihp.oisc.regs[21][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1579),
    .D(_00780_),
    .Q_N(_12696_),
    .Q(\top_ihp.oisc.regs[21][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1580),
    .D(_00781_),
    .Q_N(_12695_),
    .Q(\top_ihp.oisc.regs[21][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][17]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1581),
    .D(_00782_),
    .Q_N(_12694_),
    .Q(\top_ihp.oisc.regs[21][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1582),
    .D(_00783_),
    .Q_N(_12693_),
    .Q(\top_ihp.oisc.regs[21][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1583),
    .D(_00784_),
    .Q_N(_12692_),
    .Q(\top_ihp.oisc.regs[21][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1584),
    .D(_00785_),
    .Q_N(_12691_),
    .Q(\top_ihp.oisc.regs[21][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1585),
    .D(_00786_),
    .Q_N(_12690_),
    .Q(\top_ihp.oisc.regs[21][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1586),
    .D(_00787_),
    .Q_N(_12689_),
    .Q(\top_ihp.oisc.regs[21][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1587),
    .D(_00788_),
    .Q_N(_12688_),
    .Q(\top_ihp.oisc.regs[21][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1588),
    .D(_00789_),
    .Q_N(_12687_),
    .Q(\top_ihp.oisc.regs[21][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1589),
    .D(_00790_),
    .Q_N(_12686_),
    .Q(\top_ihp.oisc.regs[21][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1590),
    .D(_00791_),
    .Q_N(_12685_),
    .Q(\top_ihp.oisc.regs[21][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][26]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1591),
    .D(_00792_),
    .Q_N(_12684_),
    .Q(\top_ihp.oisc.regs[21][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1592),
    .D(_00793_),
    .Q_N(_12683_),
    .Q(\top_ihp.oisc.regs[21][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1593),
    .D(_00794_),
    .Q_N(_12682_),
    .Q(\top_ihp.oisc.regs[21][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][29]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1594),
    .D(_00795_),
    .Q_N(_12681_),
    .Q(\top_ihp.oisc.regs[21][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1595),
    .D(_00796_),
    .Q_N(_12680_),
    .Q(\top_ihp.oisc.regs[21][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1596),
    .D(_00797_),
    .Q_N(_12679_),
    .Q(\top_ihp.oisc.regs[21][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1597),
    .D(_00798_),
    .Q_N(_12678_),
    .Q(\top_ihp.oisc.regs[21][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1598),
    .D(_00799_),
    .Q_N(_12677_),
    .Q(\top_ihp.oisc.regs[21][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1599),
    .D(_00800_),
    .Q_N(_12676_),
    .Q(\top_ihp.oisc.regs[21][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1600),
    .D(_00801_),
    .Q_N(_12675_),
    .Q(\top_ihp.oisc.regs[21][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1601),
    .D(_00802_),
    .Q_N(_12674_),
    .Q(\top_ihp.oisc.regs[21][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1602),
    .D(_00803_),
    .Q_N(_12673_),
    .Q(\top_ihp.oisc.regs[21][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1603),
    .D(_00804_),
    .Q_N(_12672_),
    .Q(\top_ihp.oisc.regs[21][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1604),
    .D(_00805_),
    .Q_N(_12671_),
    .Q(\top_ihp.oisc.regs[21][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1605),
    .D(_00806_),
    .Q_N(_12670_),
    .Q(\top_ihp.oisc.regs[22][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1606),
    .D(_00807_),
    .Q_N(_12669_),
    .Q(\top_ihp.oisc.regs[22][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1607),
    .D(_00808_),
    .Q_N(_12668_),
    .Q(\top_ihp.oisc.regs[22][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1608),
    .D(_00809_),
    .Q_N(_12667_),
    .Q(\top_ihp.oisc.regs[22][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1609),
    .D(_00810_),
    .Q_N(_12666_),
    .Q(\top_ihp.oisc.regs[22][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1610),
    .D(_00811_),
    .Q_N(_12665_),
    .Q(\top_ihp.oisc.regs[22][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][15]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1611),
    .D(_00812_),
    .Q_N(_12664_),
    .Q(\top_ihp.oisc.regs[22][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][16]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1612),
    .D(_00813_),
    .Q_N(_12663_),
    .Q(\top_ihp.oisc.regs[22][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1613),
    .D(_00814_),
    .Q_N(_12662_),
    .Q(\top_ihp.oisc.regs[22][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1614),
    .D(_00815_),
    .Q_N(_12661_),
    .Q(\top_ihp.oisc.regs[22][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1615),
    .D(_00816_),
    .Q_N(_12660_),
    .Q(\top_ihp.oisc.regs[22][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1616),
    .D(_00817_),
    .Q_N(_12659_),
    .Q(\top_ihp.oisc.regs[22][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1617),
    .D(_00818_),
    .Q_N(_12658_),
    .Q(\top_ihp.oisc.regs[22][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1618),
    .D(_00819_),
    .Q_N(_12657_),
    .Q(\top_ihp.oisc.regs[22][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1619),
    .D(_00820_),
    .Q_N(_12656_),
    .Q(\top_ihp.oisc.regs[22][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1620),
    .D(_00821_),
    .Q_N(_12655_),
    .Q(\top_ihp.oisc.regs[22][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1621),
    .D(_00822_),
    .Q_N(_12654_),
    .Q(\top_ihp.oisc.regs[22][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1622),
    .D(_00823_),
    .Q_N(_12653_),
    .Q(\top_ihp.oisc.regs[22][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1623),
    .D(_00824_),
    .Q_N(_12652_),
    .Q(\top_ihp.oisc.regs[22][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1624),
    .D(_00825_),
    .Q_N(_12651_),
    .Q(\top_ihp.oisc.regs[22][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1625),
    .D(_00826_),
    .Q_N(_12650_),
    .Q(\top_ihp.oisc.regs[22][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1626),
    .D(_00827_),
    .Q_N(_12649_),
    .Q(\top_ihp.oisc.regs[22][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1627),
    .D(_00828_),
    .Q_N(_12648_),
    .Q(\top_ihp.oisc.regs[22][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1628),
    .D(_00829_),
    .Q_N(_12647_),
    .Q(\top_ihp.oisc.regs[22][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1629),
    .D(_00830_),
    .Q_N(_12646_),
    .Q(\top_ihp.oisc.regs[22][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1630),
    .D(_00831_),
    .Q_N(_12645_),
    .Q(\top_ihp.oisc.regs[22][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1631),
    .D(_00832_),
    .Q_N(_12644_),
    .Q(\top_ihp.oisc.regs[22][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1632),
    .D(_00833_),
    .Q_N(_12643_),
    .Q(\top_ihp.oisc.regs[22][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1633),
    .D(_00834_),
    .Q_N(_12642_),
    .Q(\top_ihp.oisc.regs[22][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1634),
    .D(_00835_),
    .Q_N(_12641_),
    .Q(\top_ihp.oisc.regs[22][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1635),
    .D(_00836_),
    .Q_N(_12640_),
    .Q(\top_ihp.oisc.regs[22][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1636),
    .D(_00837_),
    .Q_N(_12639_),
    .Q(\top_ihp.oisc.regs[22][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1637),
    .D(_00838_),
    .Q_N(_12638_),
    .Q(\top_ihp.oisc.regs[23][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1638),
    .D(_00839_),
    .Q_N(_12637_),
    .Q(\top_ihp.oisc.regs[23][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1639),
    .D(_00840_),
    .Q_N(_12636_),
    .Q(\top_ihp.oisc.regs[23][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1640),
    .D(_00841_),
    .Q_N(_12635_),
    .Q(\top_ihp.oisc.regs[23][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1641),
    .D(_00842_),
    .Q_N(_12634_),
    .Q(\top_ihp.oisc.regs[23][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1642),
    .D(_00843_),
    .Q_N(_12633_),
    .Q(\top_ihp.oisc.regs[23][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1643),
    .D(_00844_),
    .Q_N(_12632_),
    .Q(\top_ihp.oisc.regs[23][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1644),
    .D(_00845_),
    .Q_N(_12631_),
    .Q(\top_ihp.oisc.regs[23][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1645),
    .D(_00846_),
    .Q_N(_12630_),
    .Q(\top_ihp.oisc.regs[23][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1646),
    .D(_00847_),
    .Q_N(_12629_),
    .Q(\top_ihp.oisc.regs[23][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1647),
    .D(_00848_),
    .Q_N(_12628_),
    .Q(\top_ihp.oisc.regs[23][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1648),
    .D(_00849_),
    .Q_N(_12627_),
    .Q(\top_ihp.oisc.regs[23][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1649),
    .D(_00850_),
    .Q_N(_12626_),
    .Q(\top_ihp.oisc.regs[23][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1650),
    .D(_00851_),
    .Q_N(_12625_),
    .Q(\top_ihp.oisc.regs[23][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1651),
    .D(_00852_),
    .Q_N(_12624_),
    .Q(\top_ihp.oisc.regs[23][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][23]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1652),
    .D(_00853_),
    .Q_N(_12623_),
    .Q(\top_ihp.oisc.regs[23][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1653),
    .D(_00854_),
    .Q_N(_12622_),
    .Q(\top_ihp.oisc.regs[23][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1654),
    .D(_00855_),
    .Q_N(_12621_),
    .Q(\top_ihp.oisc.regs[23][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1655),
    .D(_00856_),
    .Q_N(_12620_),
    .Q(\top_ihp.oisc.regs[23][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][27]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1656),
    .D(_00857_),
    .Q_N(_12619_),
    .Q(\top_ihp.oisc.regs[23][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1657),
    .D(_00858_),
    .Q_N(_12618_),
    .Q(\top_ihp.oisc.regs[23][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1658),
    .D(_00859_),
    .Q_N(_12617_),
    .Q(\top_ihp.oisc.regs[23][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1659),
    .D(_00860_),
    .Q_N(_12616_),
    .Q(\top_ihp.oisc.regs[23][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][30]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1660),
    .D(_00861_),
    .Q_N(_12615_),
    .Q(\top_ihp.oisc.regs[23][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1661),
    .D(_00862_),
    .Q_N(_12614_),
    .Q(\top_ihp.oisc.regs[23][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1662),
    .D(_00863_),
    .Q_N(_12613_),
    .Q(\top_ihp.oisc.regs[23][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1663),
    .D(_00864_),
    .Q_N(_12612_),
    .Q(\top_ihp.oisc.regs[23][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1664),
    .D(_00865_),
    .Q_N(_12611_),
    .Q(\top_ihp.oisc.regs[23][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1665),
    .D(_00866_),
    .Q_N(_12610_),
    .Q(\top_ihp.oisc.regs[23][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1666),
    .D(_00867_),
    .Q_N(_12609_),
    .Q(\top_ihp.oisc.regs[23][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1667),
    .D(_00868_),
    .Q_N(_12608_),
    .Q(\top_ihp.oisc.regs[23][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1668),
    .D(_00869_),
    .Q_N(_12607_),
    .Q(\top_ihp.oisc.regs[23][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1669),
    .D(_00870_),
    .Q_N(_12606_),
    .Q(\top_ihp.oisc.regs[24][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1670),
    .D(_00871_),
    .Q_N(_12605_),
    .Q(\top_ihp.oisc.regs[24][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1671),
    .D(_00872_),
    .Q_N(_12604_),
    .Q(\top_ihp.oisc.regs[24][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1672),
    .D(_00873_),
    .Q_N(_12603_),
    .Q(\top_ihp.oisc.regs[24][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][13]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1673),
    .D(_00874_),
    .Q_N(_12602_),
    .Q(\top_ihp.oisc.regs[24][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1674),
    .D(_00875_),
    .Q_N(_12601_),
    .Q(\top_ihp.oisc.regs[24][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1675),
    .D(_00876_),
    .Q_N(_12600_),
    .Q(\top_ihp.oisc.regs[24][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1676),
    .D(_00877_),
    .Q_N(_12599_),
    .Q(\top_ihp.oisc.regs[24][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][17]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1677),
    .D(_00878_),
    .Q_N(_12598_),
    .Q(\top_ihp.oisc.regs[24][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][18]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1678),
    .D(_00879_),
    .Q_N(_12597_),
    .Q(\top_ihp.oisc.regs[24][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][19]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1679),
    .D(_00880_),
    .Q_N(_12596_),
    .Q(\top_ihp.oisc.regs[24][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1680),
    .D(_00881_),
    .Q_N(_12595_),
    .Q(\top_ihp.oisc.regs[24][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1681),
    .D(_00882_),
    .Q_N(_12594_),
    .Q(\top_ihp.oisc.regs[24][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1682),
    .D(_00883_),
    .Q_N(_12593_),
    .Q(\top_ihp.oisc.regs[24][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1683),
    .D(_00884_),
    .Q_N(_12592_),
    .Q(\top_ihp.oisc.regs[24][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1684),
    .D(_00885_),
    .Q_N(_12591_),
    .Q(\top_ihp.oisc.regs[24][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1685),
    .D(_00886_),
    .Q_N(_12590_),
    .Q(\top_ihp.oisc.regs[24][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][25]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1686),
    .D(_00887_),
    .Q_N(_12589_),
    .Q(\top_ihp.oisc.regs[24][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1687),
    .D(_00888_),
    .Q_N(_12588_),
    .Q(\top_ihp.oisc.regs[24][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1688),
    .D(_00889_),
    .Q_N(_12587_),
    .Q(\top_ihp.oisc.regs[24][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1689),
    .D(_00890_),
    .Q_N(_12586_),
    .Q(\top_ihp.oisc.regs[24][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1690),
    .D(_00891_),
    .Q_N(_12585_),
    .Q(\top_ihp.oisc.regs[24][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1691),
    .D(_00892_),
    .Q_N(_12584_),
    .Q(\top_ihp.oisc.regs[24][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1692),
    .D(_00893_),
    .Q_N(_12583_),
    .Q(\top_ihp.oisc.regs[24][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1693),
    .D(_00894_),
    .Q_N(_12582_),
    .Q(\top_ihp.oisc.regs[24][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1694),
    .D(_00895_),
    .Q_N(_12581_),
    .Q(\top_ihp.oisc.regs[24][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1695),
    .D(_00896_),
    .Q_N(_12580_),
    .Q(\top_ihp.oisc.regs[24][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1696),
    .D(_00897_),
    .Q_N(_12579_),
    .Q(\top_ihp.oisc.regs[24][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1697),
    .D(_00898_),
    .Q_N(_12578_),
    .Q(\top_ihp.oisc.regs[24][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1698),
    .D(_00899_),
    .Q_N(_12577_),
    .Q(\top_ihp.oisc.regs[24][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1699),
    .D(_00900_),
    .Q_N(_12576_),
    .Q(\top_ihp.oisc.regs[24][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1700),
    .D(_00901_),
    .Q_N(_12575_),
    .Q(\top_ihp.oisc.regs[24][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1701),
    .D(_00902_),
    .Q_N(_12574_),
    .Q(\top_ihp.oisc.regs[25][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1702),
    .D(_00903_),
    .Q_N(_12573_),
    .Q(\top_ihp.oisc.regs[25][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1703),
    .D(_00904_),
    .Q_N(_12572_),
    .Q(\top_ihp.oisc.regs[25][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1704),
    .D(_00905_),
    .Q_N(_12571_),
    .Q(\top_ihp.oisc.regs[25][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1705),
    .D(_00906_),
    .Q_N(_12570_),
    .Q(\top_ihp.oisc.regs[25][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1706),
    .D(_00907_),
    .Q_N(_12569_),
    .Q(\top_ihp.oisc.regs[25][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1707),
    .D(_00908_),
    .Q_N(_12568_),
    .Q(\top_ihp.oisc.regs[25][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1708),
    .D(_00909_),
    .Q_N(_12567_),
    .Q(\top_ihp.oisc.regs[25][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1709),
    .D(_00910_),
    .Q_N(_12566_),
    .Q(\top_ihp.oisc.regs[25][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1710),
    .D(_00911_),
    .Q_N(_12565_),
    .Q(\top_ihp.oisc.regs[25][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1711),
    .D(_00912_),
    .Q_N(_12564_),
    .Q(\top_ihp.oisc.regs[25][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1712),
    .D(_00913_),
    .Q_N(_12563_),
    .Q(\top_ihp.oisc.regs[25][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1713),
    .D(_00914_),
    .Q_N(_12562_),
    .Q(\top_ihp.oisc.regs[25][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1714),
    .D(_00915_),
    .Q_N(_12561_),
    .Q(\top_ihp.oisc.regs[25][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1715),
    .D(_00916_),
    .Q_N(_12560_),
    .Q(\top_ihp.oisc.regs[25][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1716),
    .D(_00917_),
    .Q_N(_12559_),
    .Q(\top_ihp.oisc.regs[25][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1717),
    .D(_00918_),
    .Q_N(_12558_),
    .Q(\top_ihp.oisc.regs[25][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][25]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1718),
    .D(_00919_),
    .Q_N(_12557_),
    .Q(\top_ihp.oisc.regs[25][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1719),
    .D(_00920_),
    .Q_N(_12556_),
    .Q(\top_ihp.oisc.regs[25][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1720),
    .D(_00921_),
    .Q_N(_12555_),
    .Q(\top_ihp.oisc.regs[25][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1721),
    .D(_00922_),
    .Q_N(_12554_),
    .Q(\top_ihp.oisc.regs[25][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1722),
    .D(_00923_),
    .Q_N(_12553_),
    .Q(\top_ihp.oisc.regs[25][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1723),
    .D(_00924_),
    .Q_N(_12552_),
    .Q(\top_ihp.oisc.regs[25][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1724),
    .D(_00925_),
    .Q_N(_12551_),
    .Q(\top_ihp.oisc.regs[25][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1725),
    .D(_00926_),
    .Q_N(_12550_),
    .Q(\top_ihp.oisc.regs[25][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1726),
    .D(_00927_),
    .Q_N(_12549_),
    .Q(\top_ihp.oisc.regs[25][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1727),
    .D(_00928_),
    .Q_N(_12548_),
    .Q(\top_ihp.oisc.regs[25][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1728),
    .D(_00929_),
    .Q_N(_12547_),
    .Q(\top_ihp.oisc.regs[25][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1729),
    .D(_00930_),
    .Q_N(_12546_),
    .Q(\top_ihp.oisc.regs[25][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1730),
    .D(_00931_),
    .Q_N(_12545_),
    .Q(\top_ihp.oisc.regs[25][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1731),
    .D(_00932_),
    .Q_N(_12544_),
    .Q(\top_ihp.oisc.regs[25][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1732),
    .D(_00933_),
    .Q_N(_12543_),
    .Q(\top_ihp.oisc.regs[25][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1733),
    .D(_00934_),
    .Q_N(_12542_),
    .Q(\top_ihp.oisc.regs[26][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1734),
    .D(_00935_),
    .Q_N(_12541_),
    .Q(\top_ihp.oisc.regs[26][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1735),
    .D(_00936_),
    .Q_N(_12540_),
    .Q(\top_ihp.oisc.regs[26][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1736),
    .D(_00937_),
    .Q_N(_12539_),
    .Q(\top_ihp.oisc.regs[26][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1737),
    .D(_00938_),
    .Q_N(_12538_),
    .Q(\top_ihp.oisc.regs[26][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1738),
    .D(_00939_),
    .Q_N(_12537_),
    .Q(\top_ihp.oisc.regs[26][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1739),
    .D(_00940_),
    .Q_N(_12536_),
    .Q(\top_ihp.oisc.regs[26][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1740),
    .D(_00941_),
    .Q_N(_12535_),
    .Q(\top_ihp.oisc.regs[26][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1741),
    .D(_00942_),
    .Q_N(_12534_),
    .Q(\top_ihp.oisc.regs[26][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][18]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1742),
    .D(_00943_),
    .Q_N(_12533_),
    .Q(\top_ihp.oisc.regs[26][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1743),
    .D(_00944_),
    .Q_N(_12532_),
    .Q(\top_ihp.oisc.regs[26][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1744),
    .D(_00945_),
    .Q_N(_12531_),
    .Q(\top_ihp.oisc.regs[26][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1745),
    .D(_00946_),
    .Q_N(_12530_),
    .Q(\top_ihp.oisc.regs[26][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1746),
    .D(_00947_),
    .Q_N(_12529_),
    .Q(\top_ihp.oisc.regs[26][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][22]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1747),
    .D(_00948_),
    .Q_N(_12528_),
    .Q(\top_ihp.oisc.regs[26][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1748),
    .D(_00949_),
    .Q_N(_12527_),
    .Q(\top_ihp.oisc.regs[26][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][24]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1749),
    .D(_00950_),
    .Q_N(_12526_),
    .Q(\top_ihp.oisc.regs[26][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1750),
    .D(_00951_),
    .Q_N(_12525_),
    .Q(\top_ihp.oisc.regs[26][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1751),
    .D(_00952_),
    .Q_N(_12524_),
    .Q(\top_ihp.oisc.regs[26][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1752),
    .D(_00953_),
    .Q_N(_12523_),
    .Q(\top_ihp.oisc.regs[26][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1753),
    .D(_00954_),
    .Q_N(_12522_),
    .Q(\top_ihp.oisc.regs[26][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1754),
    .D(_00955_),
    .Q_N(_12521_),
    .Q(\top_ihp.oisc.regs[26][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1755),
    .D(_00956_),
    .Q_N(_12520_),
    .Q(\top_ihp.oisc.regs[26][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][30]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1756),
    .D(_00957_),
    .Q_N(_12519_),
    .Q(\top_ihp.oisc.regs[26][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1757),
    .D(_00958_),
    .Q_N(_12518_),
    .Q(\top_ihp.oisc.regs[26][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1758),
    .D(_00959_),
    .Q_N(_12517_),
    .Q(\top_ihp.oisc.regs[26][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1759),
    .D(_00960_),
    .Q_N(_12516_),
    .Q(\top_ihp.oisc.regs[26][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1760),
    .D(_00961_),
    .Q_N(_12515_),
    .Q(\top_ihp.oisc.regs[26][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1761),
    .D(_00962_),
    .Q_N(_12514_),
    .Q(\top_ihp.oisc.regs[26][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1762),
    .D(_00963_),
    .Q_N(_12513_),
    .Q(\top_ihp.oisc.regs[26][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1763),
    .D(_00964_),
    .Q_N(_12512_),
    .Q(\top_ihp.oisc.regs[26][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1764),
    .D(_00965_),
    .Q_N(_12511_),
    .Q(\top_ihp.oisc.regs[26][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1765),
    .D(_00966_),
    .Q_N(_12510_),
    .Q(\top_ihp.oisc.regs[27][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1766),
    .D(_00967_),
    .Q_N(_12509_),
    .Q(\top_ihp.oisc.regs[27][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1767),
    .D(_00968_),
    .Q_N(_12508_),
    .Q(\top_ihp.oisc.regs[27][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1768),
    .D(_00969_),
    .Q_N(_12507_),
    .Q(\top_ihp.oisc.regs[27][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1769),
    .D(_00970_),
    .Q_N(_12506_),
    .Q(\top_ihp.oisc.regs[27][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1770),
    .D(_00971_),
    .Q_N(_12505_),
    .Q(\top_ihp.oisc.regs[27][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1771),
    .D(_00972_),
    .Q_N(_12504_),
    .Q(\top_ihp.oisc.regs[27][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1772),
    .D(_00973_),
    .Q_N(_12503_),
    .Q(\top_ihp.oisc.regs[27][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][17]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1773),
    .D(_00974_),
    .Q_N(_12502_),
    .Q(\top_ihp.oisc.regs[27][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1774),
    .D(_00975_),
    .Q_N(_12501_),
    .Q(\top_ihp.oisc.regs[27][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1775),
    .D(_00976_),
    .Q_N(_12500_),
    .Q(\top_ihp.oisc.regs[27][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1776),
    .D(_00977_),
    .Q_N(_12499_),
    .Q(\top_ihp.oisc.regs[27][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1777),
    .D(_00978_),
    .Q_N(_12498_),
    .Q(\top_ihp.oisc.regs[27][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][21]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1778),
    .D(_00979_),
    .Q_N(_12497_),
    .Q(\top_ihp.oisc.regs[27][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1779),
    .D(_00980_),
    .Q_N(_12496_),
    .Q(\top_ihp.oisc.regs[27][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1780),
    .D(_00981_),
    .Q_N(_12495_),
    .Q(\top_ihp.oisc.regs[27][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1781),
    .D(_00982_),
    .Q_N(_12494_),
    .Q(\top_ihp.oisc.regs[27][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][25]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1782),
    .D(_00983_),
    .Q_N(_12493_),
    .Q(\top_ihp.oisc.regs[27][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1783),
    .D(_00984_),
    .Q_N(_12492_),
    .Q(\top_ihp.oisc.regs[27][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1784),
    .D(_00985_),
    .Q_N(_12491_),
    .Q(\top_ihp.oisc.regs[27][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1785),
    .D(_00986_),
    .Q_N(_12490_),
    .Q(\top_ihp.oisc.regs[27][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1786),
    .D(_00987_),
    .Q_N(_12489_),
    .Q(\top_ihp.oisc.regs[27][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1787),
    .D(_00988_),
    .Q_N(_12488_),
    .Q(\top_ihp.oisc.regs[27][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1788),
    .D(_00989_),
    .Q_N(_12487_),
    .Q(\top_ihp.oisc.regs[27][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1789),
    .D(_00990_),
    .Q_N(_12486_),
    .Q(\top_ihp.oisc.regs[27][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1790),
    .D(_00991_),
    .Q_N(_12485_),
    .Q(\top_ihp.oisc.regs[27][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1791),
    .D(_00992_),
    .Q_N(_12484_),
    .Q(\top_ihp.oisc.regs[27][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1792),
    .D(_00993_),
    .Q_N(_12483_),
    .Q(\top_ihp.oisc.regs[27][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1793),
    .D(_00994_),
    .Q_N(_12482_),
    .Q(\top_ihp.oisc.regs[27][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1794),
    .D(_00995_),
    .Q_N(_12481_),
    .Q(\top_ihp.oisc.regs[27][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1795),
    .D(_00996_),
    .Q_N(_12480_),
    .Q(\top_ihp.oisc.regs[27][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1796),
    .D(_00997_),
    .Q_N(_12479_),
    .Q(\top_ihp.oisc.regs[27][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1797),
    .D(_00998_),
    .Q_N(_12478_),
    .Q(\top_ihp.oisc.regs[28][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1798),
    .D(_00999_),
    .Q_N(_12477_),
    .Q(\top_ihp.oisc.regs[28][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1799),
    .D(_01000_),
    .Q_N(_12476_),
    .Q(\top_ihp.oisc.regs[28][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1800),
    .D(_01001_),
    .Q_N(_12475_),
    .Q(\top_ihp.oisc.regs[28][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][13]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1801),
    .D(_01002_),
    .Q_N(_12474_),
    .Q(\top_ihp.oisc.regs[28][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1802),
    .D(_01003_),
    .Q_N(_12473_),
    .Q(\top_ihp.oisc.regs[28][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1803),
    .D(_01004_),
    .Q_N(_12472_),
    .Q(\top_ihp.oisc.regs[28][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][16]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1804),
    .D(_01005_),
    .Q_N(_12471_),
    .Q(\top_ihp.oisc.regs[28][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][17]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1805),
    .D(_01006_),
    .Q_N(_12470_),
    .Q(\top_ihp.oisc.regs[28][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1806),
    .D(_01007_),
    .Q_N(_12469_),
    .Q(\top_ihp.oisc.regs[28][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1807),
    .D(_01008_),
    .Q_N(_12468_),
    .Q(\top_ihp.oisc.regs[28][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1808),
    .D(_01009_),
    .Q_N(_12467_),
    .Q(\top_ihp.oisc.regs[28][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1809),
    .D(_01010_),
    .Q_N(_12466_),
    .Q(\top_ihp.oisc.regs[28][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1810),
    .D(_01011_),
    .Q_N(_12465_),
    .Q(\top_ihp.oisc.regs[28][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1811),
    .D(_01012_),
    .Q_N(_12464_),
    .Q(\top_ihp.oisc.regs[28][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1812),
    .D(_01013_),
    .Q_N(_12463_),
    .Q(\top_ihp.oisc.regs[28][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][24]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1813),
    .D(_01014_),
    .Q_N(_12462_),
    .Q(\top_ihp.oisc.regs[28][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1814),
    .D(_01015_),
    .Q_N(_12461_),
    .Q(\top_ihp.oisc.regs[28][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1815),
    .D(_01016_),
    .Q_N(_12460_),
    .Q(\top_ihp.oisc.regs[28][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1816),
    .D(_01017_),
    .Q_N(_12459_),
    .Q(\top_ihp.oisc.regs[28][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1817),
    .D(_01018_),
    .Q_N(_12458_),
    .Q(\top_ihp.oisc.regs[28][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1818),
    .D(_01019_),
    .Q_N(_12457_),
    .Q(\top_ihp.oisc.regs[28][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1819),
    .D(_01020_),
    .Q_N(_12456_),
    .Q(\top_ihp.oisc.regs[28][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1820),
    .D(_01021_),
    .Q_N(_12455_),
    .Q(\top_ihp.oisc.regs[28][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1821),
    .D(_01022_),
    .Q_N(_12454_),
    .Q(\top_ihp.oisc.regs[28][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1822),
    .D(_01023_),
    .Q_N(_12453_),
    .Q(\top_ihp.oisc.regs[28][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1823),
    .D(_01024_),
    .Q_N(_12452_),
    .Q(\top_ihp.oisc.regs[28][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1824),
    .D(_01025_),
    .Q_N(_12451_),
    .Q(\top_ihp.oisc.regs[28][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1825),
    .D(_01026_),
    .Q_N(_12450_),
    .Q(\top_ihp.oisc.regs[28][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1826),
    .D(_01027_),
    .Q_N(_12449_),
    .Q(\top_ihp.oisc.regs[28][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1827),
    .D(_01028_),
    .Q_N(_12448_),
    .Q(\top_ihp.oisc.regs[28][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1828),
    .D(_01029_),
    .Q_N(_12447_),
    .Q(\top_ihp.oisc.regs[28][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1829),
    .D(_01030_),
    .Q_N(_12446_),
    .Q(\top_ihp.oisc.regs[29][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1830),
    .D(_01031_),
    .Q_N(_12445_),
    .Q(\top_ihp.oisc.regs[29][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1831),
    .D(_01032_),
    .Q_N(_12444_),
    .Q(\top_ihp.oisc.regs[29][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1832),
    .D(_01033_),
    .Q_N(_12443_),
    .Q(\top_ihp.oisc.regs[29][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1833),
    .D(_01034_),
    .Q_N(_12442_),
    .Q(\top_ihp.oisc.regs[29][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1834),
    .D(_01035_),
    .Q_N(_12441_),
    .Q(\top_ihp.oisc.regs[29][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1835),
    .D(_01036_),
    .Q_N(_12440_),
    .Q(\top_ihp.oisc.regs[29][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1836),
    .D(_01037_),
    .Q_N(_12439_),
    .Q(\top_ihp.oisc.regs[29][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][17]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1837),
    .D(_01038_),
    .Q_N(_12438_),
    .Q(\top_ihp.oisc.regs[29][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1838),
    .D(_01039_),
    .Q_N(_12437_),
    .Q(\top_ihp.oisc.regs[29][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1839),
    .D(_01040_),
    .Q_N(_12436_),
    .Q(\top_ihp.oisc.regs[29][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1840),
    .D(_01041_),
    .Q_N(_12435_),
    .Q(\top_ihp.oisc.regs[29][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1841),
    .D(_01042_),
    .Q_N(_12434_),
    .Q(\top_ihp.oisc.regs[29][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1842),
    .D(_01043_),
    .Q_N(_12433_),
    .Q(\top_ihp.oisc.regs[29][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1843),
    .D(_01044_),
    .Q_N(_12432_),
    .Q(\top_ihp.oisc.regs[29][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1844),
    .D(_01045_),
    .Q_N(_12431_),
    .Q(\top_ihp.oisc.regs[29][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1845),
    .D(_01046_),
    .Q_N(_12430_),
    .Q(\top_ihp.oisc.regs[29][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1846),
    .D(_01047_),
    .Q_N(_12429_),
    .Q(\top_ihp.oisc.regs[29][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1847),
    .D(_01048_),
    .Q_N(_12428_),
    .Q(\top_ihp.oisc.regs[29][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1848),
    .D(_01049_),
    .Q_N(_12427_),
    .Q(\top_ihp.oisc.regs[29][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][28]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1849),
    .D(_01050_),
    .Q_N(_12426_),
    .Q(\top_ihp.oisc.regs[29][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1850),
    .D(_01051_),
    .Q_N(_12425_),
    .Q(\top_ihp.oisc.regs[29][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1851),
    .D(_01052_),
    .Q_N(_12424_),
    .Q(\top_ihp.oisc.regs[29][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1852),
    .D(_01053_),
    .Q_N(_12423_),
    .Q(\top_ihp.oisc.regs[29][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1853),
    .D(_01054_),
    .Q_N(_12422_),
    .Q(\top_ihp.oisc.regs[29][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1854),
    .D(_01055_),
    .Q_N(_12421_),
    .Q(\top_ihp.oisc.regs[29][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1855),
    .D(_01056_),
    .Q_N(_12420_),
    .Q(\top_ihp.oisc.regs[29][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1856),
    .D(_01057_),
    .Q_N(_12419_),
    .Q(\top_ihp.oisc.regs[29][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1857),
    .D(_01058_),
    .Q_N(_12418_),
    .Q(\top_ihp.oisc.regs[29][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1858),
    .D(_01059_),
    .Q_N(_12417_),
    .Q(\top_ihp.oisc.regs[29][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1859),
    .D(_01060_),
    .Q_N(_12416_),
    .Q(\top_ihp.oisc.regs[29][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1860),
    .D(_01061_),
    .Q_N(_12415_),
    .Q(\top_ihp.oisc.regs[29][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1164),
    .D(_01062_),
    .Q_N(_12414_),
    .Q(\top_ihp.oisc.regs[2][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1176),
    .D(_01063_),
    .Q_N(_12413_),
    .Q(\top_ihp.oisc.regs[2][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1178),
    .D(_01064_),
    .Q_N(_12412_),
    .Q(\top_ihp.oisc.regs[2][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1176),
    .D(_01065_),
    .Q_N(_12411_),
    .Q(\top_ihp.oisc.regs[2][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1228),
    .D(_01066_),
    .Q_N(_12410_),
    .Q(\top_ihp.oisc.regs[2][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1186),
    .D(_01067_),
    .Q_N(_12409_),
    .Q(\top_ihp.oisc.regs[2][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1177),
    .D(_01068_),
    .Q_N(_12408_),
    .Q(\top_ihp.oisc.regs[2][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1228),
    .D(_01069_),
    .Q_N(_12407_),
    .Q(\top_ihp.oisc.regs[2][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1185),
    .D(_01070_),
    .Q_N(_12406_),
    .Q(\top_ihp.oisc.regs[2][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1188),
    .D(_01071_),
    .Q_N(_12405_),
    .Q(\top_ihp.oisc.regs[2][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1187),
    .D(_01072_),
    .Q_N(_12404_),
    .Q(\top_ihp.oisc.regs[2][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1187),
    .D(_01073_),
    .Q_N(_12403_),
    .Q(\top_ihp.oisc.regs[2][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1165),
    .D(_01074_),
    .Q_N(_12402_),
    .Q(\top_ihp.oisc.regs[2][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1230),
    .D(_01075_),
    .Q_N(_12401_),
    .Q(\top_ihp.oisc.regs[2][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1237),
    .D(_01076_),
    .Q_N(_12400_),
    .Q(\top_ihp.oisc.regs[2][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1165),
    .D(_01077_),
    .Q_N(_12399_),
    .Q(\top_ihp.oisc.regs[2][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1237),
    .D(_01078_),
    .Q_N(_12398_),
    .Q(\top_ihp.oisc.regs[2][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1237),
    .D(_01079_),
    .Q_N(_12397_),
    .Q(\top_ihp.oisc.regs[2][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1231),
    .D(_01080_),
    .Q_N(_12396_),
    .Q(\top_ihp.oisc.regs[2][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1238),
    .D(_01081_),
    .Q_N(_12395_),
    .Q(\top_ihp.oisc.regs[2][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1238),
    .D(_01082_),
    .Q_N(_12394_),
    .Q(\top_ihp.oisc.regs[2][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1231),
    .D(_01083_),
    .Q_N(_12393_),
    .Q(\top_ihp.oisc.regs[2][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1231),
    .D(_01084_),
    .Q_N(_12392_),
    .Q(\top_ihp.oisc.regs[2][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1228),
    .D(_01085_),
    .Q_N(_12391_),
    .Q(\top_ihp.oisc.regs[2][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1187),
    .D(_01086_),
    .Q_N(_12390_),
    .Q(\top_ihp.oisc.regs[2][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1187),
    .D(_01087_),
    .Q_N(_12389_),
    .Q(\top_ihp.oisc.regs[2][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1186),
    .D(_01088_),
    .Q_N(_12388_),
    .Q(\top_ihp.oisc.regs[2][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1186),
    .D(_01089_),
    .Q_N(_12387_),
    .Q(\top_ihp.oisc.regs[2][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1178),
    .D(_01090_),
    .Q_N(_12386_),
    .Q(\top_ihp.oisc.regs[2][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1178),
    .D(_01091_),
    .Q_N(_12385_),
    .Q(\top_ihp.oisc.regs[2][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1178),
    .D(_01092_),
    .Q_N(_12384_),
    .Q(\top_ihp.oisc.regs[2][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1178),
    .D(_01093_),
    .Q_N(_12383_),
    .Q(\top_ihp.oisc.regs[2][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1861),
    .D(_01094_),
    .Q_N(_12382_),
    .Q(\top_ihp.oisc.regs[30][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1862),
    .D(_01095_),
    .Q_N(_12381_),
    .Q(\top_ihp.oisc.regs[30][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1863),
    .D(_01096_),
    .Q_N(_12380_),
    .Q(\top_ihp.oisc.regs[30][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1864),
    .D(_01097_),
    .Q_N(_12379_),
    .Q(\top_ihp.oisc.regs[30][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1865),
    .D(_01098_),
    .Q_N(_12378_),
    .Q(\top_ihp.oisc.regs[30][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1866),
    .D(_01099_),
    .Q_N(_12377_),
    .Q(\top_ihp.oisc.regs[30][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][15]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1867),
    .D(_01100_),
    .Q_N(_12376_),
    .Q(\top_ihp.oisc.regs[30][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1868),
    .D(_01101_),
    .Q_N(_12375_),
    .Q(\top_ihp.oisc.regs[30][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][17]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1869),
    .D(_01102_),
    .Q_N(_12374_),
    .Q(\top_ihp.oisc.regs[30][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1870),
    .D(_01103_),
    .Q_N(_12373_),
    .Q(\top_ihp.oisc.regs[30][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1871),
    .D(_01104_),
    .Q_N(_12372_),
    .Q(\top_ihp.oisc.regs[30][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1872),
    .D(_01105_),
    .Q_N(_12371_),
    .Q(\top_ihp.oisc.regs[30][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][20]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1873),
    .D(_01106_),
    .Q_N(_12370_),
    .Q(\top_ihp.oisc.regs[30][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1874),
    .D(_01107_),
    .Q_N(_12369_),
    .Q(\top_ihp.oisc.regs[30][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][22]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1875),
    .D(_01108_),
    .Q_N(_12368_),
    .Q(\top_ihp.oisc.regs[30][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1876),
    .D(_01109_),
    .Q_N(_12367_),
    .Q(\top_ihp.oisc.regs[30][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1877),
    .D(_01110_),
    .Q_N(_12366_),
    .Q(\top_ihp.oisc.regs[30][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1878),
    .D(_01111_),
    .Q_N(_12365_),
    .Q(\top_ihp.oisc.regs[30][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][26]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1879),
    .D(_01112_),
    .Q_N(_12364_),
    .Q(\top_ihp.oisc.regs[30][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1880),
    .D(_01113_),
    .Q_N(_12363_),
    .Q(\top_ihp.oisc.regs[30][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][28]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1881),
    .D(_01114_),
    .Q_N(_12362_),
    .Q(\top_ihp.oisc.regs[30][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1882),
    .D(_01115_),
    .Q_N(_12361_),
    .Q(\top_ihp.oisc.regs[30][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1883),
    .D(_01116_),
    .Q_N(_12360_),
    .Q(\top_ihp.oisc.regs[30][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1884),
    .D(_01117_),
    .Q_N(_12359_),
    .Q(\top_ihp.oisc.regs[30][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1885),
    .D(_01118_),
    .Q_N(_12358_),
    .Q(\top_ihp.oisc.regs[30][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1886),
    .D(_01119_),
    .Q_N(_12357_),
    .Q(\top_ihp.oisc.regs[30][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1887),
    .D(_01120_),
    .Q_N(_12356_),
    .Q(\top_ihp.oisc.regs[30][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1888),
    .D(_01121_),
    .Q_N(_12355_),
    .Q(\top_ihp.oisc.regs[30][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1889),
    .D(_01122_),
    .Q_N(_12354_),
    .Q(\top_ihp.oisc.regs[30][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1890),
    .D(_01123_),
    .Q_N(_12353_),
    .Q(\top_ihp.oisc.regs[30][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1891),
    .D(_01124_),
    .Q_N(_12352_),
    .Q(\top_ihp.oisc.regs[30][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1892),
    .D(_01125_),
    .Q_N(_12351_),
    .Q(\top_ihp.oisc.regs[30][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1893),
    .D(_01126_),
    .Q_N(_12350_),
    .Q(\top_ihp.oisc.regs[31][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1894),
    .D(_01127_),
    .Q_N(_12349_),
    .Q(\top_ihp.oisc.regs[31][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1895),
    .D(_01128_),
    .Q_N(_12348_),
    .Q(\top_ihp.oisc.regs[31][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1896),
    .D(_01129_),
    .Q_N(_12347_),
    .Q(\top_ihp.oisc.regs[31][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][13]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1897),
    .D(_01130_),
    .Q_N(_12346_),
    .Q(\top_ihp.oisc.regs[31][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1898),
    .D(_01131_),
    .Q_N(_12345_),
    .Q(\top_ihp.oisc.regs[31][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1899),
    .D(_01132_),
    .Q_N(_12344_),
    .Q(\top_ihp.oisc.regs[31][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1900),
    .D(_01133_),
    .Q_N(_12343_),
    .Q(\top_ihp.oisc.regs[31][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1901),
    .D(_01134_),
    .Q_N(_12342_),
    .Q(\top_ihp.oisc.regs[31][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1902),
    .D(_01135_),
    .Q_N(_12341_),
    .Q(\top_ihp.oisc.regs[31][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1903),
    .D(_01136_),
    .Q_N(_12340_),
    .Q(\top_ihp.oisc.regs[31][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1904),
    .D(_01137_),
    .Q_N(_12339_),
    .Q(\top_ihp.oisc.regs[31][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][20]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1905),
    .D(_01138_),
    .Q_N(_12338_),
    .Q(\top_ihp.oisc.regs[31][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][21]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1906),
    .D(_01139_),
    .Q_N(_12337_),
    .Q(\top_ihp.oisc.regs[31][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1907),
    .D(_01140_),
    .Q_N(_12336_),
    .Q(\top_ihp.oisc.regs[31][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1908),
    .D(_01141_),
    .Q_N(_12335_),
    .Q(\top_ihp.oisc.regs[31][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][24]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1909),
    .D(_01142_),
    .Q_N(_12334_),
    .Q(\top_ihp.oisc.regs[31][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1910),
    .D(_01143_),
    .Q_N(_12333_),
    .Q(\top_ihp.oisc.regs[31][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1911),
    .D(_01144_),
    .Q_N(_12332_),
    .Q(\top_ihp.oisc.regs[31][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1912),
    .D(_01145_),
    .Q_N(_12331_),
    .Q(\top_ihp.oisc.regs[31][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1913),
    .D(_01146_),
    .Q_N(_12330_),
    .Q(\top_ihp.oisc.regs[31][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][29]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1914),
    .D(_01147_),
    .Q_N(_12329_),
    .Q(\top_ihp.oisc.regs[31][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1915),
    .D(_01148_),
    .Q_N(_12328_),
    .Q(\top_ihp.oisc.regs[31][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1916),
    .D(_01149_),
    .Q_N(_12327_),
    .Q(\top_ihp.oisc.regs[31][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1917),
    .D(_01150_),
    .Q_N(_12326_),
    .Q(\top_ihp.oisc.regs[31][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1918),
    .D(_01151_),
    .Q_N(_12325_),
    .Q(\top_ihp.oisc.regs[31][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1919),
    .D(_01152_),
    .Q_N(_12324_),
    .Q(\top_ihp.oisc.regs[31][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1920),
    .D(_01153_),
    .Q_N(_12323_),
    .Q(\top_ihp.oisc.regs[31][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1921),
    .D(_01154_),
    .Q_N(_12322_),
    .Q(\top_ihp.oisc.regs[31][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1922),
    .D(_01155_),
    .Q_N(_12321_),
    .Q(\top_ihp.oisc.regs[31][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1923),
    .D(_01156_),
    .Q_N(_12320_),
    .Q(\top_ihp.oisc.regs[31][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1924),
    .D(_01157_),
    .Q_N(_12319_),
    .Q(\top_ihp.oisc.regs[31][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1925),
    .D(_01158_),
    .Q_N(_12318_),
    .Q(\top_ihp.oisc.regs[32][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1926),
    .D(_01159_),
    .Q_N(_12317_),
    .Q(\top_ihp.oisc.regs[32][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][11]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1927),
    .D(_01160_),
    .Q_N(_12316_),
    .Q(\top_ihp.oisc.regs[32][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][12]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1928),
    .D(_01161_),
    .Q_N(_12315_),
    .Q(\top_ihp.oisc.regs[32][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][13]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1929),
    .D(_01162_),
    .Q_N(_12314_),
    .Q(\top_ihp.oisc.regs[32][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][14]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1930),
    .D(_01163_),
    .Q_N(_12313_),
    .Q(\top_ihp.oisc.regs[32][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][15]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1931),
    .D(_01164_),
    .Q_N(_12312_),
    .Q(\top_ihp.oisc.regs[32][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1932),
    .D(_01165_),
    .Q_N(_12311_),
    .Q(\top_ihp.oisc.regs[32][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][17]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1933),
    .D(_01166_),
    .Q_N(_12310_),
    .Q(\top_ihp.oisc.regs[32][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][18]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1934),
    .D(_01167_),
    .Q_N(_12309_),
    .Q(\top_ihp.oisc.regs[32][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][19]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1935),
    .D(_01168_),
    .Q_N(_12308_),
    .Q(\top_ihp.oisc.regs[32][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][1]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1936),
    .D(_01169_),
    .Q_N(_12307_),
    .Q(\top_ihp.oisc.regs[32][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][20]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1937),
    .D(_01170_),
    .Q_N(_12306_),
    .Q(\top_ihp.oisc.regs[32][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][21]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1938),
    .D(_01171_),
    .Q_N(_12305_),
    .Q(\top_ihp.oisc.regs[32][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][22]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1939),
    .D(_01172_),
    .Q_N(_12304_),
    .Q(\top_ihp.oisc.regs[32][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][23]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1940),
    .D(_01173_),
    .Q_N(_12303_),
    .Q(\top_ihp.oisc.regs[32][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][24]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1941),
    .D(_01174_),
    .Q_N(_12302_),
    .Q(\top_ihp.oisc.regs[32][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][25]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1942),
    .D(_01175_),
    .Q_N(_12301_),
    .Q(\top_ihp.oisc.regs[32][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][26]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1943),
    .D(_01176_),
    .Q_N(_12300_),
    .Q(\top_ihp.oisc.regs[32][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][27]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1944),
    .D(_01177_),
    .Q_N(_12299_),
    .Q(\top_ihp.oisc.regs[32][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][28]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1945),
    .D(_01178_),
    .Q_N(_12298_),
    .Q(\top_ihp.oisc.regs[32][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][29]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1946),
    .D(_01179_),
    .Q_N(_12297_),
    .Q(\top_ihp.oisc.regs[32][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][2]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1947),
    .D(_01180_),
    .Q_N(_12296_),
    .Q(\top_ihp.oisc.regs[32][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][30]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1948),
    .D(_01181_),
    .Q_N(_12295_),
    .Q(\top_ihp.oisc.regs[32][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][31]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1949),
    .D(_01182_),
    .Q_N(_12294_),
    .Q(\top_ihp.oisc.regs[32][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][3]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1950),
    .D(_01183_),
    .Q_N(_12293_),
    .Q(\top_ihp.oisc.regs[32][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1951),
    .D(_01184_),
    .Q_N(_12292_),
    .Q(\top_ihp.oisc.regs[32][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][5]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1952),
    .D(_01185_),
    .Q_N(_12291_),
    .Q(\top_ihp.oisc.regs[32][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1953),
    .D(_01186_),
    .Q_N(_12290_),
    .Q(\top_ihp.oisc.regs[32][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][7]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1954),
    .D(_01187_),
    .Q_N(_12289_),
    .Q(\top_ihp.oisc.regs[32][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][8]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1955),
    .D(_01188_),
    .Q_N(_12288_),
    .Q(\top_ihp.oisc.regs[32][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1956),
    .D(_01189_),
    .Q_N(_12287_),
    .Q(\top_ihp.oisc.regs[32][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1240),
    .D(_01190_),
    .Q_N(_12286_),
    .Q(\top_ihp.oisc.regs[33][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1274),
    .D(_01191_),
    .Q_N(_12285_),
    .Q(\top_ihp.oisc.regs[33][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1272),
    .D(_01192_),
    .Q_N(_12284_),
    .Q(\top_ihp.oisc.regs[33][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1275),
    .D(_01193_),
    .Q_N(_12283_),
    .Q(\top_ihp.oisc.regs[33][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1240),
    .D(_01194_),
    .Q_N(_12282_),
    .Q(\top_ihp.oisc.regs[33][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1201),
    .D(_01195_),
    .Q_N(_12281_),
    .Q(\top_ihp.oisc.regs[33][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1193),
    .D(_01196_),
    .Q_N(_12280_),
    .Q(\top_ihp.oisc.regs[33][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1260),
    .D(_01197_),
    .Q_N(_12279_),
    .Q(\top_ihp.oisc.regs[33][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1210),
    .D(_01198_),
    .Q_N(_12278_),
    .Q(\top_ihp.oisc.regs[33][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1220),
    .D(_01199_),
    .Q_N(_12277_),
    .Q(\top_ihp.oisc.regs[33][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1220),
    .D(_01200_),
    .Q_N(_12276_),
    .Q(\top_ihp.oisc.regs[33][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1291),
    .D(_01201_),
    .Q_N(_12275_),
    .Q(\top_ihp.oisc.regs[33][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1258),
    .D(_01202_),
    .Q_N(_12274_),
    .Q(\top_ihp.oisc.regs[33][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1337),
    .D(_01203_),
    .Q_N(_12273_),
    .Q(\top_ihp.oisc.regs[33][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1357),
    .D(_01204_),
    .Q_N(_12272_),
    .Q(\top_ihp.oisc.regs[33][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1258),
    .D(_01205_),
    .Q_N(_12271_),
    .Q(\top_ihp.oisc.regs[33][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1354),
    .D(_01206_),
    .Q_N(_12270_),
    .Q(\top_ihp.oisc.regs[33][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1354),
    .D(_01207_),
    .Q_N(_12269_),
    .Q(\top_ihp.oisc.regs[33][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1354),
    .D(_01208_),
    .Q_N(_12268_),
    .Q(\top_ihp.oisc.regs[33][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1256),
    .D(_01209_),
    .Q_N(_12267_),
    .Q(\top_ihp.oisc.regs[33][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1367),
    .D(_01210_),
    .Q_N(_12266_),
    .Q(\top_ihp.oisc.regs[33][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1367),
    .D(_01211_),
    .Q_N(_12265_),
    .Q(\top_ihp.oisc.regs[33][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1363),
    .D(_01212_),
    .Q_N(_12264_),
    .Q(\top_ihp.oisc.regs[33][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1364),
    .D(_01213_),
    .Q_N(_12263_),
    .Q(\top_ihp.oisc.regs[33][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1297),
    .D(_01214_),
    .Q_N(_12262_),
    .Q(\top_ihp.oisc.regs[33][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1324),
    .D(_01215_),
    .Q_N(_12261_),
    .Q(\top_ihp.oisc.regs[33][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1294),
    .D(_01216_),
    .Q_N(_12260_),
    .Q(\top_ihp.oisc.regs[33][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1321),
    .D(_01217_),
    .Q_N(_12259_),
    .Q(\top_ihp.oisc.regs[33][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1302),
    .D(_01218_),
    .Q_N(_12258_),
    .Q(\top_ihp.oisc.regs[33][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1304),
    .D(_01219_),
    .Q_N(_12257_),
    .Q(\top_ihp.oisc.regs[33][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1285),
    .D(_01220_),
    .Q_N(_12256_),
    .Q(\top_ihp.oisc.regs[33][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1293),
    .D(_01221_),
    .Q_N(_12255_),
    .Q(\top_ihp.oisc.regs[33][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1345),
    .D(_01222_),
    .Q_N(_12254_),
    .Q(\top_ihp.oisc.regs[34][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1284),
    .D(_01223_),
    .Q_N(_12253_),
    .Q(\top_ihp.oisc.regs[34][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1277),
    .D(_01224_),
    .Q_N(_12252_),
    .Q(\top_ihp.oisc.regs[34][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1277),
    .D(_01225_),
    .Q_N(_12251_),
    .Q(\top_ihp.oisc.regs[34][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1244),
    .D(_01226_),
    .Q_N(_12250_),
    .Q(\top_ihp.oisc.regs[34][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1196),
    .D(_01227_),
    .Q_N(_12249_),
    .Q(\top_ihp.oisc.regs[34][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1197),
    .D(_01228_),
    .Q_N(\top_ihp.oisc.regs[34][15] ),
    .Q(_00210_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1247),
    .D(_01229_),
    .Q_N(_12248_),
    .Q(\top_ihp.oisc.regs[34][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1210),
    .D(_01230_),
    .Q_N(_12247_),
    .Q(\top_ihp.oisc.regs[34][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1251),
    .D(_01231_),
    .Q_N(_12246_),
    .Q(\top_ihp.oisc.regs[34][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1210),
    .D(_01232_),
    .Q_N(_12245_),
    .Q(\top_ihp.oisc.regs[34][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1290),
    .D(_01233_),
    .Q_N(_12244_),
    .Q(\top_ihp.oisc.regs[34][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1260),
    .D(_01234_),
    .Q_N(_12243_),
    .Q(\top_ihp.oisc.regs[34][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1253),
    .D(_01235_),
    .Q_N(_12242_),
    .Q(\top_ihp.oisc.regs[34][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1351),
    .D(_01236_),
    .Q_N(_12241_),
    .Q(\top_ihp.oisc.regs[34][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1266),
    .D(_01237_),
    .Q_N(_12240_),
    .Q(\top_ihp.oisc.regs[34][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1353),
    .D(_01238_),
    .Q_N(_12239_),
    .Q(\top_ihp.oisc.regs[34][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1355),
    .D(_01239_),
    .Q_N(_12238_),
    .Q(\top_ihp.oisc.regs[34][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1378),
    .D(_01240_),
    .Q_N(_12237_),
    .Q(\top_ihp.oisc.regs[34][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1379),
    .D(_01241_),
    .Q_N(_12236_),
    .Q(\top_ihp.oisc.regs[34][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1379),
    .D(_01242_),
    .Q_N(_12235_),
    .Q(\top_ihp.oisc.regs[34][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1337),
    .D(_01243_),
    .Q_N(_12234_),
    .Q(\top_ihp.oisc.regs[34][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1335),
    .D(_01244_),
    .Q_N(_12233_),
    .Q(\top_ihp.oisc.regs[34][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1364),
    .D(_01245_),
    .Q_N(_12232_),
    .Q(\top_ihp.oisc.regs[34][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1297),
    .D(_01246_),
    .Q_N(\top_ihp.oisc.regs[34][31] ),
    .Q(_00211_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1291),
    .D(_01247_),
    .Q_N(_12231_),
    .Q(\top_ihp.oisc.regs[34][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1319),
    .D(_01248_),
    .Q_N(_12230_),
    .Q(\top_ihp.oisc.regs[34][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1288),
    .D(_01249_),
    .Q_N(_12229_),
    .Q(\top_ihp.oisc.regs[34][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1306),
    .D(_01250_),
    .Q_N(_12228_),
    .Q(\top_ihp.oisc.regs[34][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1307),
    .D(_01251_),
    .Q_N(_12227_),
    .Q(\top_ihp.oisc.regs[34][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1306),
    .D(_01252_),
    .Q_N(_12226_),
    .Q(\top_ihp.oisc.regs[34][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1293),
    .D(_01253_),
    .Q_N(_12225_),
    .Q(\top_ihp.oisc.regs[34][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1345),
    .D(_01254_),
    .Q_N(_12224_),
    .Q(\top_ihp.oisc.regs[35][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1277),
    .D(_01255_),
    .Q_N(_12223_),
    .Q(\top_ihp.oisc.regs[35][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1220),
    .D(_01256_),
    .Q_N(\top_ihp.oisc.regs[35][11] ),
    .Q(_00212_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1204),
    .D(_01257_),
    .Q_N(_12222_),
    .Q(\top_ihp.oisc.regs[35][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1219),
    .D(_01258_),
    .Q_N(_12221_),
    .Q(\top_ihp.oisc.regs[35][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1287),
    .D(_01259_),
    .Q_N(_12220_),
    .Q(\top_ihp.oisc.regs[35][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1196),
    .D(_01260_),
    .Q_N(_12219_),
    .Q(\top_ihp.oisc.regs[35][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1244),
    .D(_01261_),
    .Q_N(_12218_),
    .Q(\top_ihp.oisc.regs[35][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1210),
    .D(_01262_),
    .Q_N(_12217_),
    .Q(\top_ihp.oisc.regs[35][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1220),
    .D(_01263_),
    .Q_N(_12216_),
    .Q(\top_ihp.oisc.regs[35][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1216),
    .D(_01264_),
    .Q_N(_12215_),
    .Q(\top_ihp.oisc.regs[35][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1290),
    .D(_01265_),
    .Q_N(_12214_),
    .Q(\top_ihp.oisc.regs[35][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1264),
    .D(_01266_),
    .Q_N(_12213_),
    .Q(\top_ihp.oisc.regs[35][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1353),
    .D(_01267_),
    .Q_N(_12212_),
    .Q(\top_ihp.oisc.regs[35][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1353),
    .D(_01268_),
    .Q_N(_12211_),
    .Q(\top_ihp.oisc.regs[35][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1264),
    .D(_01269_),
    .Q_N(_12210_),
    .Q(\top_ihp.oisc.regs[35][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1353),
    .D(_01270_),
    .Q_N(_12209_),
    .Q(\top_ihp.oisc.regs[35][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1355),
    .D(_01271_),
    .Q_N(_12208_),
    .Q(\top_ihp.oisc.regs[35][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1378),
    .D(_01272_),
    .Q_N(_12207_),
    .Q(\top_ihp.oisc.regs[35][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1380),
    .D(_01273_),
    .Q_N(_12206_),
    .Q(\top_ihp.oisc.regs[35][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1367),
    .D(_01274_),
    .Q_N(_12205_),
    .Q(\top_ihp.oisc.regs[35][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1342),
    .D(_01275_),
    .Q_N(_12204_),
    .Q(\top_ihp.oisc.regs[35][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1363),
    .D(_01276_),
    .Q_N(_12203_),
    .Q(\top_ihp.oisc.regs[35][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1363),
    .D(_01277_),
    .Q_N(_12202_),
    .Q(\top_ihp.oisc.regs[35][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1297),
    .D(_01278_),
    .Q_N(\top_ihp.oisc.regs[35][31] ),
    .Q(_00213_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1324),
    .D(_01279_),
    .Q_N(_12201_),
    .Q(\top_ihp.oisc.regs[35][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1320),
    .D(_01280_),
    .Q_N(_12200_),
    .Q(\top_ihp.oisc.regs[35][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1321),
    .D(_01281_),
    .Q_N(_12199_),
    .Q(\top_ihp.oisc.regs[35][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1306),
    .D(_01282_),
    .Q_N(_12198_),
    .Q(\top_ihp.oisc.regs[35][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1307),
    .D(_01283_),
    .Q_N(_12197_),
    .Q(\top_ihp.oisc.regs[35][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1306),
    .D(_01284_),
    .Q_N(_12196_),
    .Q(\top_ihp.oisc.regs[35][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1285),
    .D(_01285_),
    .Q_N(_12195_),
    .Q(\top_ihp.oisc.regs[35][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1260),
    .D(_01286_),
    .Q_N(_12194_),
    .Q(\top_ihp.oisc.regs[36][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1280),
    .D(_01287_),
    .Q_N(_12193_),
    .Q(\top_ihp.oisc.regs[36][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1201),
    .D(_01288_),
    .Q_N(_12192_),
    .Q(\top_ihp.oisc.regs[36][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1273),
    .D(_01289_),
    .Q_N(_12191_),
    .Q(\top_ihp.oisc.regs[36][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1244),
    .D(_01290_),
    .Q_N(_12190_),
    .Q(\top_ihp.oisc.regs[36][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1287),
    .D(_01291_),
    .Q_N(_12189_),
    .Q(\top_ihp.oisc.regs[36][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1191),
    .D(_01292_),
    .Q_N(_12188_),
    .Q(\top_ihp.oisc.regs[36][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1244),
    .D(_01293_),
    .Q_N(_12187_),
    .Q(\top_ihp.oisc.regs[36][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1200),
    .D(_01294_),
    .Q_N(_12186_),
    .Q(\top_ihp.oisc.regs[36][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1334),
    .D(_01295_),
    .Q_N(_12185_),
    .Q(\top_ihp.oisc.regs[36][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1209),
    .D(_01296_),
    .Q_N(_12184_),
    .Q(\top_ihp.oisc.regs[36][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1334),
    .D(_01297_),
    .Q_N(_12183_),
    .Q(\top_ihp.oisc.regs[36][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1260),
    .D(_01298_),
    .Q_N(_12182_),
    .Q(\top_ihp.oisc.regs[36][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1247),
    .D(_01299_),
    .Q_N(_12181_),
    .Q(\top_ihp.oisc.regs[36][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1351),
    .D(_01300_),
    .Q_N(_12180_),
    .Q(\top_ihp.oisc.regs[36][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1266),
    .D(_01301_),
    .Q_N(_12179_),
    .Q(\top_ihp.oisc.regs[36][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1359),
    .D(_01302_),
    .Q_N(_12178_),
    .Q(\top_ihp.oisc.regs[36][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1381),
    .D(_01303_),
    .Q_N(_12177_),
    .Q(\top_ihp.oisc.regs[36][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1381),
    .D(_01304_),
    .Q_N(_12176_),
    .Q(\top_ihp.oisc.regs[36][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1383),
    .D(_01305_),
    .Q_N(_12175_),
    .Q(\top_ihp.oisc.regs[36][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1383),
    .D(_01306_),
    .Q_N(_12174_),
    .Q(\top_ihp.oisc.regs[36][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1336),
    .D(_01307_),
    .Q_N(_12173_),
    .Q(\top_ihp.oisc.regs[36][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1247),
    .D(_01308_),
    .Q_N(_12172_),
    .Q(\top_ihp.oisc.regs[36][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1364),
    .D(_01309_),
    .Q_N(_12171_),
    .Q(\top_ihp.oisc.regs[36][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1297),
    .D(_01310_),
    .Q_N(_12170_),
    .Q(\top_ihp.oisc.regs[36][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1324),
    .D(_01311_),
    .Q_N(_12169_),
    .Q(\top_ihp.oisc.regs[36][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1320),
    .D(_01312_),
    .Q_N(_12168_),
    .Q(\top_ihp.oisc.regs[36][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1307),
    .D(_01313_),
    .Q_N(_12167_),
    .Q(\top_ihp.oisc.regs[36][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1304),
    .D(_01314_),
    .Q_N(_12166_),
    .Q(\top_ihp.oisc.regs[36][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1303),
    .D(_01315_),
    .Q_N(_12165_),
    .Q(\top_ihp.oisc.regs[36][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1303),
    .D(_01316_),
    .Q_N(_12164_),
    .Q(\top_ihp.oisc.regs[36][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1293),
    .D(_01317_),
    .Q_N(_12163_),
    .Q(\top_ihp.oisc.regs[36][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1349),
    .D(_01318_),
    .Q_N(_12162_),
    .Q(\top_ihp.oisc.regs[37][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1284),
    .D(_01319_),
    .Q_N(_12161_),
    .Q(\top_ihp.oisc.regs[37][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1278),
    .D(_01320_),
    .Q_N(_12160_),
    .Q(\top_ihp.oisc.regs[37][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1277),
    .D(_01321_),
    .Q_N(_12159_),
    .Q(\top_ihp.oisc.regs[37][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1267),
    .D(_01322_),
    .Q_N(_12158_),
    .Q(\top_ihp.oisc.regs[37][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1287),
    .D(_01323_),
    .Q_N(_12157_),
    .Q(\top_ihp.oisc.regs[37][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1205),
    .D(_01324_),
    .Q_N(_12156_),
    .Q(\top_ihp.oisc.regs[37][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1266),
    .D(_01325_),
    .Q_N(_12155_),
    .Q(\top_ihp.oisc.regs[37][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1205),
    .D(_01326_),
    .Q_N(_12154_),
    .Q(\top_ihp.oisc.regs[37][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1290),
    .D(_01327_),
    .Q_N(_12153_),
    .Q(\top_ihp.oisc.regs[37][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1287),
    .D(_01328_),
    .Q_N(_12152_),
    .Q(\top_ihp.oisc.regs[37][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1296),
    .D(_01329_),
    .Q_N(_12151_),
    .Q(\top_ihp.oisc.regs[37][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1267),
    .D(_01330_),
    .Q_N(_12150_),
    .Q(\top_ihp.oisc.regs[37][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1337),
    .D(_01331_),
    .Q_N(_12149_),
    .Q(\top_ihp.oisc.regs[37][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1351),
    .D(_01332_),
    .Q_N(_12148_),
    .Q(\top_ihp.oisc.regs[37][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1266),
    .D(_01333_),
    .Q_N(_12147_),
    .Q(\top_ihp.oisc.regs[37][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1389),
    .D(_01334_),
    .Q_N(_12146_),
    .Q(\top_ihp.oisc.regs[37][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1381),
    .D(_01335_),
    .Q_N(_12145_),
    .Q(\top_ihp.oisc.regs[37][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1382),
    .D(_01336_),
    .Q_N(_12144_),
    .Q(\top_ihp.oisc.regs[37][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1389),
    .D(_01337_),
    .Q_N(_12143_),
    .Q(\top_ihp.oisc.regs[37][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1383),
    .D(_01338_),
    .Q_N(_12142_),
    .Q(\top_ihp.oisc.regs[37][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1342),
    .D(_01339_),
    .Q_N(_12141_),
    .Q(\top_ihp.oisc.regs[37][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1364),
    .D(_01340_),
    .Q_N(_12140_),
    .Q(\top_ihp.oisc.regs[37][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1370),
    .D(_01341_),
    .Q_N(_12139_),
    .Q(\top_ihp.oisc.regs[37][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1323),
    .D(_01342_),
    .Q_N(_12138_),
    .Q(\top_ihp.oisc.regs[37][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1329),
    .D(_01343_),
    .Q_N(_12137_),
    .Q(\top_ihp.oisc.regs[37][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1326),
    .D(_01344_),
    .Q_N(_12136_),
    .Q(\top_ihp.oisc.regs[37][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1314),
    .D(_01345_),
    .Q_N(_12135_),
    .Q(\top_ihp.oisc.regs[37][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1314),
    .D(_01346_),
    .Q_N(_12134_),
    .Q(\top_ihp.oisc.regs[37][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1314),
    .D(_01347_),
    .Q_N(_12133_),
    .Q(\top_ihp.oisc.regs[37][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1287),
    .D(_01348_),
    .Q_N(_12132_),
    .Q(\top_ihp.oisc.regs[37][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1294),
    .D(_01349_),
    .Q_N(_12131_),
    .Q(\top_ihp.oisc.regs[37][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1349),
    .D(_01350_),
    .Q_N(_12130_),
    .Q(\top_ihp.oisc.regs[38][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1282),
    .D(_01351_),
    .Q_N(_12129_),
    .Q(\top_ihp.oisc.regs[38][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1273),
    .D(_01352_),
    .Q_N(_12128_),
    .Q(\top_ihp.oisc.regs[38][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1278),
    .D(_01353_),
    .Q_N(_12127_),
    .Q(\top_ihp.oisc.regs[38][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1245),
    .D(_01354_),
    .Q_N(_12126_),
    .Q(\top_ihp.oisc.regs[38][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1196),
    .D(_01355_),
    .Q_N(_12125_),
    .Q(\top_ihp.oisc.regs[38][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1215),
    .D(_01356_),
    .Q_N(_12124_),
    .Q(\top_ihp.oisc.regs[38][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1245),
    .D(_01357_),
    .Q_N(_12123_),
    .Q(\top_ihp.oisc.regs[38][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1200),
    .D(_01358_),
    .Q_N(_12122_),
    .Q(\top_ihp.oisc.regs[38][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1220),
    .D(_01359_),
    .Q_N(_12121_),
    .Q(\top_ihp.oisc.regs[38][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1216),
    .D(_01360_),
    .Q_N(_12120_),
    .Q(\top_ihp.oisc.regs[38][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1334),
    .D(_01361_),
    .Q_N(_12119_),
    .Q(\top_ihp.oisc.regs[38][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1267),
    .D(_01362_),
    .Q_N(_12118_),
    .Q(\top_ihp.oisc.regs[38][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1341),
    .D(_01363_),
    .Q_N(_12117_),
    .Q(\top_ihp.oisc.regs[38][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1357),
    .D(_01364_),
    .Q_N(_12116_),
    .Q(\top_ihp.oisc.regs[38][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1266),
    .D(_01365_),
    .Q_N(_12115_),
    .Q(\top_ihp.oisc.regs[38][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1378),
    .D(_01366_),
    .Q_N(_12114_),
    .Q(\top_ihp.oisc.regs[38][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1382),
    .D(_01367_),
    .Q_N(_12113_),
    .Q(\top_ihp.oisc.regs[38][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1383),
    .D(_01368_),
    .Q_N(_12112_),
    .Q(\top_ihp.oisc.regs[38][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1383),
    .D(_01369_),
    .Q_N(_12111_),
    .Q(\top_ihp.oisc.regs[38][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1367),
    .D(_01370_),
    .Q_N(_12110_),
    .Q(\top_ihp.oisc.regs[38][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1336),
    .D(_01371_),
    .Q_N(_12109_),
    .Q(\top_ihp.oisc.regs[38][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1334),
    .D(_01372_),
    .Q_N(_12108_),
    .Q(\top_ihp.oisc.regs[38][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1364),
    .D(_01373_),
    .Q_N(_12107_),
    .Q(\top_ihp.oisc.regs[38][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1297),
    .D(_01374_),
    .Q_N(_12106_),
    .Q(\top_ihp.oisc.regs[38][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1324),
    .D(_01375_),
    .Q_N(_12105_),
    .Q(\top_ihp.oisc.regs[38][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1321),
    .D(_01376_),
    .Q_N(_12104_),
    .Q(\top_ihp.oisc.regs[38][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1321),
    .D(_01377_),
    .Q_N(_12103_),
    .Q(\top_ihp.oisc.regs[38][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1302),
    .D(_01378_),
    .Q_N(_12102_),
    .Q(\top_ihp.oisc.regs[38][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1304),
    .D(_01379_),
    .Q_N(_12101_),
    .Q(\top_ihp.oisc.regs[38][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1319),
    .D(_01380_),
    .Q_N(_12100_),
    .Q(\top_ihp.oisc.regs[38][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1282),
    .D(_01381_),
    .Q_N(_12099_),
    .Q(\top_ihp.oisc.regs[38][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1350),
    .D(_01382_),
    .Q_N(_12098_),
    .Q(\top_ihp.oisc.regs[39][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1284),
    .D(_01383_),
    .Q_N(_12097_),
    .Q(\top_ihp.oisc.regs[39][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1273),
    .D(_01384_),
    .Q_N(_12096_),
    .Q(\top_ihp.oisc.regs[39][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1273),
    .D(_01385_),
    .Q_N(_12095_),
    .Q(\top_ihp.oisc.regs[39][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1219),
    .D(_01386_),
    .Q_N(_12094_),
    .Q(\top_ihp.oisc.regs[39][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1287),
    .D(_01387_),
    .Q_N(_12093_),
    .Q(\top_ihp.oisc.regs[39][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1193),
    .D(_01388_),
    .Q_N(_12092_),
    .Q(\top_ihp.oisc.regs[39][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1212),
    .D(_01389_),
    .Q_N(_12091_),
    .Q(\top_ihp.oisc.regs[39][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1200),
    .D(_01390_),
    .Q_N(_12090_),
    .Q(\top_ihp.oisc.regs[39][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1212),
    .D(_01391_),
    .Q_N(_12089_),
    .Q(\top_ihp.oisc.regs[39][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1216),
    .D(_01392_),
    .Q_N(_12088_),
    .Q(\top_ihp.oisc.regs[39][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1335),
    .D(_01393_),
    .Q_N(_12087_),
    .Q(\top_ihp.oisc.regs[39][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1268),
    .D(_01394_),
    .Q_N(_12086_),
    .Q(\top_ihp.oisc.regs[39][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1336),
    .D(_01395_),
    .Q_N(_12085_),
    .Q(\top_ihp.oisc.regs[39][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1358),
    .D(_01396_),
    .Q_N(_12084_),
    .Q(\top_ihp.oisc.regs[39][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1268),
    .D(_01397_),
    .Q_N(_12083_),
    .Q(\top_ihp.oisc.regs[39][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1359),
    .D(_01398_),
    .Q_N(_12082_),
    .Q(\top_ihp.oisc.regs[39][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1359),
    .D(_01399_),
    .Q_N(_12081_),
    .Q(\top_ihp.oisc.regs[39][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1360),
    .D(_01400_),
    .Q_N(_12080_),
    .Q(\top_ihp.oisc.regs[39][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1358),
    .D(_01401_),
    .Q_N(_12079_),
    .Q(\top_ihp.oisc.regs[39][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1382),
    .D(_01402_),
    .Q_N(_12078_),
    .Q(\top_ihp.oisc.regs[39][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1336),
    .D(_01403_),
    .Q_N(_12077_),
    .Q(\top_ihp.oisc.regs[39][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1363),
    .D(_01404_),
    .Q_N(_12076_),
    .Q(\top_ihp.oisc.regs[39][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1363),
    .D(_01405_),
    .Q_N(_12075_),
    .Q(\top_ihp.oisc.regs[39][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1324),
    .D(_01406_),
    .Q_N(_12074_),
    .Q(\top_ihp.oisc.regs[39][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1324),
    .D(_01407_),
    .Q_N(_12073_),
    .Q(\top_ihp.oisc.regs[39][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1319),
    .D(_01408_),
    .Q_N(_12072_),
    .Q(\top_ihp.oisc.regs[39][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1321),
    .D(_01409_),
    .Q_N(_12071_),
    .Q(\top_ihp.oisc.regs[39][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1303),
    .D(_01410_),
    .Q_N(_12070_),
    .Q(\top_ihp.oisc.regs[39][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1303),
    .D(_01411_),
    .Q_N(_12069_),
    .Q(\top_ihp.oisc.regs[39][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1303),
    .D(_01412_),
    .Q_N(_12068_),
    .Q(\top_ihp.oisc.regs[39][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1281),
    .D(_01413_),
    .Q_N(_12067_),
    .Q(\top_ihp.oisc.regs[39][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1159),
    .D(_01414_),
    .Q_N(_12066_),
    .Q(\top_ihp.oisc.regs[3][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1176),
    .D(_01415_),
    .Q_N(_12065_),
    .Q(\top_ihp.oisc.regs[3][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1176),
    .D(_01416_),
    .Q_N(_12064_),
    .Q(\top_ihp.oisc.regs[3][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1177),
    .D(_01417_),
    .Q_N(_12063_),
    .Q(\top_ihp.oisc.regs[3][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1188),
    .D(_01418_),
    .Q_N(_12062_),
    .Q(\top_ihp.oisc.regs[3][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1177),
    .D(_01419_),
    .Q_N(_12061_),
    .Q(\top_ihp.oisc.regs[3][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1176),
    .D(_01420_),
    .Q_N(_12060_),
    .Q(\top_ihp.oisc.regs[3][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1228),
    .D(_01421_),
    .Q_N(_12059_),
    .Q(\top_ihp.oisc.regs[3][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1185),
    .D(_01422_),
    .Q_N(_12058_),
    .Q(\top_ihp.oisc.regs[3][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1188),
    .D(_01423_),
    .Q_N(_12057_),
    .Q(\top_ihp.oisc.regs[3][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1185),
    .D(_01424_),
    .Q_N(_12056_),
    .Q(\top_ihp.oisc.regs[3][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1188),
    .D(_01425_),
    .Q_N(_12055_),
    .Q(\top_ihp.oisc.regs[3][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1148),
    .D(_01426_),
    .Q_N(_12054_),
    .Q(\top_ihp.oisc.regs[3][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1230),
    .D(_01427_),
    .Q_N(_12053_),
    .Q(\top_ihp.oisc.regs[3][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1239),
    .D(_01428_),
    .Q_N(_12052_),
    .Q(\top_ihp.oisc.regs[3][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1159),
    .D(_01429_),
    .Q_N(_12051_),
    .Q(\top_ihp.oisc.regs[3][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1239),
    .D(_01430_),
    .Q_N(_12050_),
    .Q(\top_ihp.oisc.regs[3][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1239),
    .D(_01431_),
    .Q_N(_12049_),
    .Q(\top_ihp.oisc.regs[3][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1230),
    .D(_01432_),
    .Q_N(_12048_),
    .Q(\top_ihp.oisc.regs[3][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1239),
    .D(_01433_),
    .Q_N(_12047_),
    .Q(\top_ihp.oisc.regs[3][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1239),
    .D(_01434_),
    .Q_N(_12046_),
    .Q(\top_ihp.oisc.regs[3][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1230),
    .D(_01435_),
    .Q_N(_12045_),
    .Q(\top_ihp.oisc.regs[3][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1229),
    .D(_01436_),
    .Q_N(_12044_),
    .Q(\top_ihp.oisc.regs[3][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1229),
    .D(_01437_),
    .Q_N(_12043_),
    .Q(\top_ihp.oisc.regs[3][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1188),
    .D(_01438_),
    .Q_N(_12042_),
    .Q(\top_ihp.oisc.regs[3][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1188),
    .D(_01439_),
    .Q_N(_12041_),
    .Q(\top_ihp.oisc.regs[3][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1185),
    .D(_01440_),
    .Q_N(_12040_),
    .Q(\top_ihp.oisc.regs[3][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1185),
    .D(_01441_),
    .Q_N(_12039_),
    .Q(\top_ihp.oisc.regs[3][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1174),
    .D(_01442_),
    .Q_N(_12038_),
    .Q(\top_ihp.oisc.regs[3][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1174),
    .D(_01443_),
    .Q_N(_12037_),
    .Q(\top_ihp.oisc.regs[3][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1177),
    .D(_01444_),
    .Q_N(_12036_),
    .Q(\top_ihp.oisc.regs[3][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1176),
    .D(_01445_),
    .Q_N(_12035_),
    .Q(\top_ihp.oisc.regs[3][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1347),
    .D(_01446_),
    .Q_N(_12034_),
    .Q(\top_ihp.oisc.regs[40][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1275),
    .D(_01447_),
    .Q_N(_12033_),
    .Q(\top_ihp.oisc.regs[40][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1275),
    .D(_01448_),
    .Q_N(_12032_),
    .Q(\top_ihp.oisc.regs[40][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1204),
    .D(_01449_),
    .Q_N(_12031_),
    .Q(\top_ihp.oisc.regs[40][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1268),
    .D(_01450_),
    .Q_N(_12030_),
    .Q(\top_ihp.oisc.regs[40][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1287),
    .D(_01451_),
    .Q_N(_12029_),
    .Q(\top_ihp.oisc.regs[40][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1195),
    .D(_01452_),
    .Q_N(_12028_),
    .Q(\top_ihp.oisc.regs[40][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1261),
    .D(_01453_),
    .Q_N(_12027_),
    .Q(\top_ihp.oisc.regs[40][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1202),
    .D(_01454_),
    .Q_N(_12026_),
    .Q(\top_ihp.oisc.regs[40][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1249),
    .D(_01455_),
    .Q_N(_12025_),
    .Q(\top_ihp.oisc.regs[40][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1217),
    .D(_01456_),
    .Q_N(_12024_),
    .Q(\top_ihp.oisc.regs[40][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1213),
    .D(_01457_),
    .Q_N(_12023_),
    .Q(\top_ihp.oisc.regs[40][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1268),
    .D(_01458_),
    .Q_N(_12022_),
    .Q(\top_ihp.oisc.regs[40][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1343),
    .D(_01459_),
    .Q_N(_12021_),
    .Q(\top_ihp.oisc.regs[40][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1358),
    .D(_01460_),
    .Q_N(_12020_),
    .Q(\top_ihp.oisc.regs[40][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1266),
    .D(_01461_),
    .Q_N(_12019_),
    .Q(\top_ihp.oisc.regs[40][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1355),
    .D(_01462_),
    .Q_N(_12018_),
    .Q(\top_ihp.oisc.regs[40][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1253),
    .D(_01463_),
    .Q_N(_12017_),
    .Q(\top_ihp.oisc.regs[40][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1252),
    .D(_01464_),
    .Q_N(_12016_),
    .Q(\top_ihp.oisc.regs[40][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1379),
    .D(_01465_),
    .Q_N(_12015_),
    .Q(\top_ihp.oisc.regs[40][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1373),
    .D(_01466_),
    .Q_N(_12014_),
    .Q(\top_ihp.oisc.regs[40][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1373),
    .D(_01467_),
    .Q_N(_12013_),
    .Q(\top_ihp.oisc.regs[40][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1339),
    .D(_01468_),
    .Q_N(_12012_),
    .Q(\top_ihp.oisc.regs[40][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1370),
    .D(_01469_),
    .Q_N(_12011_),
    .Q(\top_ihp.oisc.regs[40][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1324),
    .D(_01470_),
    .Q_N(_12010_),
    .Q(\top_ihp.oisc.regs[40][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1329),
    .D(_01471_),
    .Q_N(_12009_),
    .Q(\top_ihp.oisc.regs[40][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1326),
    .D(_01472_),
    .Q_N(_12008_),
    .Q(\top_ihp.oisc.regs[40][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1307),
    .D(_01473_),
    .Q_N(_12007_),
    .Q(\top_ihp.oisc.regs[40][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1309),
    .D(_01474_),
    .Q_N(_12006_),
    .Q(\top_ihp.oisc.regs[40][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1310),
    .D(_01475_),
    .Q_N(_12005_),
    .Q(\top_ihp.oisc.regs[40][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1301),
    .D(_01476_),
    .Q_N(_12004_),
    .Q(\top_ihp.oisc.regs[40][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1288),
    .D(_01477_),
    .Q_N(_12003_),
    .Q(\top_ihp.oisc.regs[40][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1345),
    .D(_01478_),
    .Q_N(_12002_),
    .Q(\top_ihp.oisc.regs[41][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1275),
    .D(_01479_),
    .Q_N(_12001_),
    .Q(\top_ihp.oisc.regs[41][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1202),
    .D(_01480_),
    .Q_N(_12000_),
    .Q(\top_ihp.oisc.regs[41][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1278),
    .D(_01481_),
    .Q_N(_11999_),
    .Q(\top_ihp.oisc.regs[41][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1249),
    .D(_01482_),
    .Q_N(_11998_),
    .Q(\top_ihp.oisc.regs[41][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1196),
    .D(_01483_),
    .Q_N(_11997_),
    .Q(\top_ihp.oisc.regs[41][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1193),
    .D(_01484_),
    .Q_N(_11996_),
    .Q(\top_ihp.oisc.regs[41][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1247),
    .D(_01485_),
    .Q_N(_11995_),
    .Q(\top_ihp.oisc.regs[41][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1215),
    .D(_01486_),
    .Q_N(_11994_),
    .Q(\top_ihp.oisc.regs[41][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1220),
    .D(_01487_),
    .Q_N(_11993_),
    .Q(\top_ihp.oisc.regs[41][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1287),
    .D(_01488_),
    .Q_N(_11992_),
    .Q(\top_ihp.oisc.regs[41][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1334),
    .D(_01489_),
    .Q_N(_11991_),
    .Q(\top_ihp.oisc.regs[41][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1345),
    .D(_01490_),
    .Q_N(_11990_),
    .Q(\top_ihp.oisc.regs[41][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1353),
    .D(_01491_),
    .Q_N(_11989_),
    .Q(\top_ihp.oisc.regs[41][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1347),
    .D(_01492_),
    .Q_N(_11988_),
    .Q(\top_ihp.oisc.regs[41][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1264),
    .D(_01493_),
    .Q_N(_11987_),
    .Q(\top_ihp.oisc.regs[41][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1386),
    .D(_01494_),
    .Q_N(_11986_),
    .Q(\top_ihp.oisc.regs[41][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1337),
    .D(_01495_),
    .Q_N(_11985_),
    .Q(\top_ihp.oisc.regs[41][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1366),
    .D(_01496_),
    .Q_N(_11984_),
    .Q(\top_ihp.oisc.regs[41][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1380),
    .D(_01497_),
    .Q_N(_11983_),
    .Q(\top_ihp.oisc.regs[41][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1379),
    .D(_01498_),
    .Q_N(_11982_),
    .Q(\top_ihp.oisc.regs[41][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1336),
    .D(_01499_),
    .Q_N(_11981_),
    .Q(\top_ihp.oisc.regs[41][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1364),
    .D(_01500_),
    .Q_N(_11980_),
    .Q(\top_ihp.oisc.regs[41][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1370),
    .D(_01501_),
    .Q_N(_11979_),
    .Q(\top_ihp.oisc.regs[41][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1323),
    .D(_01502_),
    .Q_N(_11978_),
    .Q(\top_ihp.oisc.regs[41][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1296),
    .D(_01503_),
    .Q_N(_11977_),
    .Q(\top_ihp.oisc.regs[41][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1320),
    .D(_01504_),
    .Q_N(_11976_),
    .Q(\top_ihp.oisc.regs[41][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1326),
    .D(_01505_),
    .Q_N(_11975_),
    .Q(\top_ihp.oisc.regs[41][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1314),
    .D(_01506_),
    .Q_N(_11974_),
    .Q(\top_ihp.oisc.regs[41][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1307),
    .D(_01507_),
    .Q_N(_11973_),
    .Q(\top_ihp.oisc.regs[41][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1288),
    .D(_01508_),
    .Q_N(_11972_),
    .Q(\top_ihp.oisc.regs[41][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1288),
    .D(_01509_),
    .Q_N(_11971_),
    .Q(\top_ihp.oisc.regs[41][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1347),
    .D(_01510_),
    .Q_N(_11970_),
    .Q(\top_ihp.oisc.regs[42][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1280),
    .D(_01511_),
    .Q_N(_11969_),
    .Q(\top_ihp.oisc.regs[42][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1277),
    .D(_01512_),
    .Q_N(_11968_),
    .Q(\top_ihp.oisc.regs[42][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1277),
    .D(_01513_),
    .Q_N(_11967_),
    .Q(\top_ihp.oisc.regs[42][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1268),
    .D(_01514_),
    .Q_N(_11966_),
    .Q(\top_ihp.oisc.regs[42][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1196),
    .D(_01515_),
    .Q_N(_11965_),
    .Q(\top_ihp.oisc.regs[42][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1197),
    .D(_01516_),
    .Q_N(_11964_),
    .Q(\top_ihp.oisc.regs[42][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1247),
    .D(_01517_),
    .Q_N(_11963_),
    .Q(\top_ihp.oisc.regs[42][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1196),
    .D(_01518_),
    .Q_N(_11962_),
    .Q(\top_ihp.oisc.regs[42][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1251),
    .D(_01519_),
    .Q_N(_11961_),
    .Q(\top_ihp.oisc.regs[42][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1212),
    .D(_01520_),
    .Q_N(_11960_),
    .Q(\top_ihp.oisc.regs[42][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1296),
    .D(_01521_),
    .Q_N(_11959_),
    .Q(\top_ihp.oisc.regs[42][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1259),
    .D(_01522_),
    .Q_N(_11958_),
    .Q(\top_ihp.oisc.regs[42][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1343),
    .D(_01523_),
    .Q_N(_11957_),
    .Q(\top_ihp.oisc.regs[42][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1259),
    .D(_01524_),
    .Q_N(_11956_),
    .Q(\top_ihp.oisc.regs[42][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1259),
    .D(_01525_),
    .Q_N(_11955_),
    .Q(\top_ihp.oisc.regs[42][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1386),
    .D(_01526_),
    .Q_N(_11954_),
    .Q(\top_ihp.oisc.regs[42][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1354),
    .D(_01527_),
    .Q_N(_11953_),
    .Q(\top_ihp.oisc.regs[42][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1342),
    .D(_01528_),
    .Q_N(_11952_),
    .Q(\top_ihp.oisc.regs[42][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1386),
    .D(_01529_),
    .Q_N(_11951_),
    .Q(\top_ihp.oisc.regs[42][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1387),
    .D(_01530_),
    .Q_N(_11950_),
    .Q(\top_ihp.oisc.regs[42][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1374),
    .D(_01531_),
    .Q_N(_11949_),
    .Q(\top_ihp.oisc.regs[42][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1363),
    .D(_01532_),
    .Q_N(_11948_),
    .Q(\top_ihp.oisc.regs[42][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1370),
    .D(_01533_),
    .Q_N(_11947_),
    .Q(\top_ihp.oisc.regs[42][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1329),
    .D(_01534_),
    .Q_N(_11946_),
    .Q(\top_ihp.oisc.regs[42][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1324),
    .D(_01535_),
    .Q_N(_11945_),
    .Q(\top_ihp.oisc.regs[42][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1326),
    .D(_01536_),
    .Q_N(_11944_),
    .Q(\top_ihp.oisc.regs[42][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1321),
    .D(_01537_),
    .Q_N(_11943_),
    .Q(\top_ihp.oisc.regs[42][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1310),
    .D(_01538_),
    .Q_N(_11942_),
    .Q(\top_ihp.oisc.regs[42][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1314),
    .D(_01539_),
    .Q_N(_11941_),
    .Q(\top_ihp.oisc.regs[42][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1306),
    .D(_01540_),
    .Q_N(_11940_),
    .Q(\top_ihp.oisc.regs[42][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1294),
    .D(_01541_),
    .Q_N(_11939_),
    .Q(\top_ihp.oisc.regs[42][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1258),
    .D(_01542_),
    .Q_N(_11938_),
    .Q(\top_ihp.oisc.regs[43][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1283),
    .D(_01543_),
    .Q_N(_11937_),
    .Q(\top_ihp.oisc.regs[43][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1205),
    .D(_01544_),
    .Q_N(_11936_),
    .Q(\top_ihp.oisc.regs[43][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1202),
    .D(_01545_),
    .Q_N(_11935_),
    .Q(\top_ihp.oisc.regs[43][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1244),
    .D(_01546_),
    .Q_N(_11934_),
    .Q(\top_ihp.oisc.regs[43][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1196),
    .D(_01547_),
    .Q_N(_11933_),
    .Q(\top_ihp.oisc.regs[43][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1204),
    .D(_01548_),
    .Q_N(_11932_),
    .Q(\top_ihp.oisc.regs[43][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1212),
    .D(_01549_),
    .Q_N(_11931_),
    .Q(\top_ihp.oisc.regs[43][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1200),
    .D(_01550_),
    .Q_N(_11930_),
    .Q(\top_ihp.oisc.regs[43][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1219),
    .D(_01551_),
    .Q_N(_11929_),
    .Q(\top_ihp.oisc.regs[43][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1211),
    .D(_01552_),
    .Q_N(_11928_),
    .Q(\top_ihp.oisc.regs[43][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1334),
    .D(_01553_),
    .Q_N(_11927_),
    .Q(\top_ihp.oisc.regs[43][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1258),
    .D(_01554_),
    .Q_N(_11926_),
    .Q(\top_ihp.oisc.regs[43][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1337),
    .D(_01555_),
    .Q_N(_11925_),
    .Q(\top_ihp.oisc.regs[43][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1351),
    .D(_01556_),
    .Q_N(_11924_),
    .Q(\top_ihp.oisc.regs[43][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1258),
    .D(_01557_),
    .Q_N(_11923_),
    .Q(\top_ihp.oisc.regs[43][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1389),
    .D(_01558_),
    .Q_N(_11922_),
    .Q(\top_ihp.oisc.regs[43][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1360),
    .D(_01559_),
    .Q_N(_11921_),
    .Q(\top_ihp.oisc.regs[43][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1360),
    .D(_01560_),
    .Q_N(_11920_),
    .Q(\top_ihp.oisc.regs[43][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1384),
    .D(_01561_),
    .Q_N(_11919_),
    .Q(\top_ihp.oisc.regs[43][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1384),
    .D(_01562_),
    .Q_N(_11918_),
    .Q(\top_ihp.oisc.regs[43][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1337),
    .D(_01563_),
    .Q_N(_11917_),
    .Q(\top_ihp.oisc.regs[43][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1335),
    .D(_01564_),
    .Q_N(_11916_),
    .Q(\top_ihp.oisc.regs[43][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1370),
    .D(_01565_),
    .Q_N(_11915_),
    .Q(\top_ihp.oisc.regs[43][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1297),
    .D(_01566_),
    .Q_N(_11914_),
    .Q(\top_ihp.oisc.regs[43][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1329),
    .D(_01567_),
    .Q_N(_11913_),
    .Q(\top_ihp.oisc.regs[43][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1319),
    .D(_01568_),
    .Q_N(_11912_),
    .Q(\top_ihp.oisc.regs[43][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1322),
    .D(_01569_),
    .Q_N(_11911_),
    .Q(\top_ihp.oisc.regs[43][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1310),
    .D(_01570_),
    .Q_N(_11910_),
    .Q(\top_ihp.oisc.regs[43][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1310),
    .D(_01571_),
    .Q_N(_11909_),
    .Q(\top_ihp.oisc.regs[43][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1282),
    .D(_01572_),
    .Q_N(_11908_),
    .Q(\top_ihp.oisc.regs[43][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1285),
    .D(_01573_),
    .Q_N(_11907_),
    .Q(\top_ihp.oisc.regs[43][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1350),
    .D(_01574_),
    .Q_N(_11906_),
    .Q(\top_ihp.oisc.regs[44][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1284),
    .D(_01575_),
    .Q_N(_11905_),
    .Q(\top_ihp.oisc.regs[44][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1277),
    .D(_01576_),
    .Q_N(_11904_),
    .Q(\top_ihp.oisc.regs[44][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1204),
    .D(_01577_),
    .Q_N(_11903_),
    .Q(\top_ihp.oisc.regs[44][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1249),
    .D(_01578_),
    .Q_N(_11902_),
    .Q(\top_ihp.oisc.regs[44][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1289),
    .D(_01579_),
    .Q_N(_11901_),
    .Q(\top_ihp.oisc.regs[44][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1204),
    .D(_01580_),
    .Q_N(_11900_),
    .Q(\top_ihp.oisc.regs[44][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1250),
    .D(_01581_),
    .Q_N(_11899_),
    .Q(\top_ihp.oisc.regs[44][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1215),
    .D(_01582_),
    .Q_N(_11898_),
    .Q(\top_ihp.oisc.regs[44][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1249),
    .D(_01583_),
    .Q_N(_11897_),
    .Q(\top_ihp.oisc.regs[44][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1219),
    .D(_01584_),
    .Q_N(_11896_),
    .Q(\top_ihp.oisc.regs[44][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1291),
    .D(_01585_),
    .Q_N(_11895_),
    .Q(\top_ihp.oisc.regs[44][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1350),
    .D(_01586_),
    .Q_N(_11894_),
    .Q(\top_ihp.oisc.regs[44][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1341),
    .D(_01587_),
    .Q_N(_11893_),
    .Q(\top_ihp.oisc.regs[44][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1358),
    .D(_01588_),
    .Q_N(_11892_),
    .Q(\top_ihp.oisc.regs[44][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1350),
    .D(_01589_),
    .Q_N(_11891_),
    .Q(\top_ihp.oisc.regs[44][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1390),
    .D(_01590_),
    .Q_N(_11890_),
    .Q(\top_ihp.oisc.regs[44][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1382),
    .D(_01591_),
    .Q_N(_11889_),
    .Q(\top_ihp.oisc.regs[44][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1360),
    .D(_01592_),
    .Q_N(_11888_),
    .Q(\top_ihp.oisc.regs[44][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1390),
    .D(_01593_),
    .Q_N(_11887_),
    .Q(\top_ihp.oisc.regs[44][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1389),
    .D(_01594_),
    .Q_N(_11886_),
    .Q(\top_ihp.oisc.regs[44][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1341),
    .D(_01595_),
    .Q_N(_11885_),
    .Q(\top_ihp.oisc.regs[44][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1363),
    .D(_01596_),
    .Q_N(_11884_),
    .Q(\top_ihp.oisc.regs[44][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1339),
    .D(_01597_),
    .Q_N(_11883_),
    .Q(\top_ihp.oisc.regs[44][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1329),
    .D(_01598_),
    .Q_N(_11882_),
    .Q(\top_ihp.oisc.regs[44][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1296),
    .D(_01599_),
    .Q_N(_11881_),
    .Q(\top_ihp.oisc.regs[44][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1326),
    .D(_01600_),
    .Q_N(_11880_),
    .Q(\top_ihp.oisc.regs[44][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1326),
    .D(_01601_),
    .Q_N(_11879_),
    .Q(\top_ihp.oisc.regs[44][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1309),
    .D(_01602_),
    .Q_N(_11878_),
    .Q(\top_ihp.oisc.regs[44][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1309),
    .D(_01603_),
    .Q_N(_11877_),
    .Q(\top_ihp.oisc.regs[44][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1301),
    .D(_01604_),
    .Q_N(_11876_),
    .Q(\top_ihp.oisc.regs[44][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1295),
    .D(_01605_),
    .Q_N(_11875_),
    .Q(\top_ihp.oisc.regs[44][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1350),
    .D(_01606_),
    .Q_N(_11874_),
    .Q(\top_ihp.oisc.regs[45][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1274),
    .D(_01607_),
    .Q_N(_11873_),
    .Q(\top_ihp.oisc.regs[45][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1202),
    .D(_01608_),
    .Q_N(_11872_),
    .Q(\top_ihp.oisc.regs[45][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1199),
    .D(_01609_),
    .Q_N(_11871_),
    .Q(\top_ihp.oisc.regs[45][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1261),
    .D(_01610_),
    .Q_N(_11870_),
    .Q(\top_ihp.oisc.regs[45][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1278),
    .D(_01611_),
    .Q_N(_11869_),
    .Q(\top_ihp.oisc.regs[45][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1193),
    .D(_01612_),
    .Q_N(_11868_),
    .Q(\top_ihp.oisc.regs[45][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1269),
    .D(_01613_),
    .Q_N(_11867_),
    .Q(\top_ihp.oisc.regs[45][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1197),
    .D(_01614_),
    .Q_N(_11866_),
    .Q(\top_ihp.oisc.regs[45][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1212),
    .D(_01615_),
    .Q_N(_11865_),
    .Q(\top_ihp.oisc.regs[45][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1219),
    .D(_01616_),
    .Q_N(_11864_),
    .Q(\top_ihp.oisc.regs[45][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1290),
    .D(_01617_),
    .Q_N(_11863_),
    .Q(\top_ihp.oisc.regs[45][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1259),
    .D(_01618_),
    .Q_N(_11862_),
    .Q(\top_ihp.oisc.regs[45][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1252),
    .D(_01619_),
    .Q_N(_11861_),
    .Q(\top_ihp.oisc.regs[45][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1352),
    .D(_01620_),
    .Q_N(_11860_),
    .Q(\top_ihp.oisc.regs[45][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1269),
    .D(_01621_),
    .Q_N(_11859_),
    .Q(\top_ihp.oisc.regs[45][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1354),
    .D(_01622_),
    .Q_N(_11858_),
    .Q(\top_ihp.oisc.regs[45][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1256),
    .D(_01623_),
    .Q_N(_11857_),
    .Q(\top_ihp.oisc.regs[45][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1366),
    .D(_01624_),
    .Q_N(_11856_),
    .Q(\top_ihp.oisc.regs[45][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1256),
    .D(_01625_),
    .Q_N(_11855_),
    .Q(\top_ihp.oisc.regs[45][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1373),
    .D(_01626_),
    .Q_N(_11854_),
    .Q(\top_ihp.oisc.regs[45][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1336),
    .D(_01627_),
    .Q_N(_11853_),
    .Q(\top_ihp.oisc.regs[45][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1365),
    .D(_01628_),
    .Q_N(_11852_),
    .Q(\top_ihp.oisc.regs[45][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1370),
    .D(_01629_),
    .Q_N(_11851_),
    .Q(\top_ihp.oisc.regs[45][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1332),
    .D(_01630_),
    .Q_N(_11850_),
    .Q(\top_ihp.oisc.regs[45][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1290),
    .D(_01631_),
    .Q_N(_11849_),
    .Q(\top_ihp.oisc.regs[45][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1327),
    .D(_01632_),
    .Q_N(_11848_),
    .Q(\top_ihp.oisc.regs[45][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1327),
    .D(_01633_),
    .Q_N(_11847_),
    .Q(\top_ihp.oisc.regs[45][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1311),
    .D(_01634_),
    .Q_N(_11846_),
    .Q(\top_ihp.oisc.regs[45][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1310),
    .D(_01635_),
    .Q_N(_11845_),
    .Q(\top_ihp.oisc.regs[45][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1282),
    .D(_01636_),
    .Q_N(_11844_),
    .Q(\top_ihp.oisc.regs[45][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1294),
    .D(_01637_),
    .Q_N(_11843_),
    .Q(\top_ihp.oisc.regs[45][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1346),
    .D(_01638_),
    .Q_N(_11842_),
    .Q(\top_ihp.oisc.regs[46][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1274),
    .D(_01639_),
    .Q_N(_11841_),
    .Q(\top_ihp.oisc.regs[46][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1201),
    .D(_01640_),
    .Q_N(_11840_),
    .Q(\top_ihp.oisc.regs[46][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1199),
    .D(_01641_),
    .Q_N(_11839_),
    .Q(\top_ihp.oisc.regs[46][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1257),
    .D(_01642_),
    .Q_N(_11838_),
    .Q(\top_ihp.oisc.regs[46][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1191),
    .D(_01643_),
    .Q_N(_11837_),
    .Q(\top_ihp.oisc.regs[46][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1209),
    .D(_01644_),
    .Q_N(_11836_),
    .Q(\top_ihp.oisc.regs[46][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1247),
    .D(_01645_),
    .Q_N(_11835_),
    .Q(\top_ihp.oisc.regs[46][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1215),
    .D(_01646_),
    .Q_N(_11834_),
    .Q(\top_ihp.oisc.regs[46][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1214),
    .D(_01647_),
    .Q_N(_11833_),
    .Q(\top_ihp.oisc.regs[46][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1209),
    .D(_01648_),
    .Q_N(_11832_),
    .Q(\top_ihp.oisc.regs[46][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1291),
    .D(_01649_),
    .Q_N(_11831_),
    .Q(\top_ihp.oisc.regs[46][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1267),
    .D(_01650_),
    .Q_N(_11830_),
    .Q(\top_ihp.oisc.regs[46][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1338),
    .D(_01651_),
    .Q_N(_11829_),
    .Q(\top_ihp.oisc.regs[46][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1351),
    .D(_01652_),
    .Q_N(_11828_),
    .Q(\top_ihp.oisc.regs[46][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1265),
    .D(_01653_),
    .Q_N(_11827_),
    .Q(\top_ihp.oisc.regs[46][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1379),
    .D(_01654_),
    .Q_N(_11826_),
    .Q(\top_ihp.oisc.regs[46][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1378),
    .D(_01655_),
    .Q_N(_11825_),
    .Q(\top_ihp.oisc.regs[46][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1379),
    .D(_01656_),
    .Q_N(_11824_),
    .Q(\top_ihp.oisc.regs[46][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1386),
    .D(_01657_),
    .Q_N(_11823_),
    .Q(\top_ihp.oisc.regs[46][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1374),
    .D(_01658_),
    .Q_N(_11822_),
    .Q(\top_ihp.oisc.regs[46][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1374),
    .D(_01659_),
    .Q_N(_11821_),
    .Q(\top_ihp.oisc.regs[46][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1365),
    .D(_01660_),
    .Q_N(_11820_),
    .Q(\top_ihp.oisc.regs[46][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1371),
    .D(_01661_),
    .Q_N(_11819_),
    .Q(\top_ihp.oisc.regs[46][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1332),
    .D(_01662_),
    .Q_N(_11818_),
    .Q(\top_ihp.oisc.regs[46][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1331),
    .D(_01663_),
    .Q_N(_11817_),
    .Q(\top_ihp.oisc.regs[46][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1328),
    .D(_01664_),
    .Q_N(_11816_),
    .Q(\top_ihp.oisc.regs[46][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1326),
    .D(_01665_),
    .Q_N(_11815_),
    .Q(\top_ihp.oisc.regs[46][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1311),
    .D(_01666_),
    .Q_N(_11814_),
    .Q(\top_ihp.oisc.regs[46][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1315),
    .D(_01667_),
    .Q_N(_11813_),
    .Q(\top_ihp.oisc.regs[46][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1301),
    .D(_01668_),
    .Q_N(_11812_),
    .Q(\top_ihp.oisc.regs[46][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1288),
    .D(_01669_),
    .Q_N(_11811_),
    .Q(\top_ihp.oisc.regs[46][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1241),
    .D(_01670_),
    .Q_N(_11810_),
    .Q(\top_ihp.oisc.regs[47][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1274),
    .D(_01671_),
    .Q_N(_11809_),
    .Q(\top_ihp.oisc.regs[47][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1272),
    .D(_01672_),
    .Q_N(_11808_),
    .Q(\top_ihp.oisc.regs[47][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1274),
    .D(_01673_),
    .Q_N(_11807_),
    .Q(\top_ihp.oisc.regs[47][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1250),
    .D(_01674_),
    .Q_N(_11806_),
    .Q(\top_ihp.oisc.regs[47][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1192),
    .D(_01675_),
    .Q_N(_11805_),
    .Q(\top_ihp.oisc.regs[47][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1192),
    .D(_01676_),
    .Q_N(_11804_),
    .Q(\top_ihp.oisc.regs[47][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1245),
    .D(_01677_),
    .Q_N(_11803_),
    .Q(\top_ihp.oisc.regs[47][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1199),
    .D(_01678_),
    .Q_N(_11802_),
    .Q(\top_ihp.oisc.regs[47][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1221),
    .D(_01679_),
    .Q_N(_11801_),
    .Q(\top_ihp.oisc.regs[47][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1211),
    .D(_01680_),
    .Q_N(_11800_),
    .Q(\top_ihp.oisc.regs[47][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1334),
    .D(_01681_),
    .Q_N(_11799_),
    .Q(\top_ihp.oisc.regs[47][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1240),
    .D(_01682_),
    .Q_N(_11798_),
    .Q(\top_ihp.oisc.regs[47][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1343),
    .D(_01683_),
    .Q_N(_11797_),
    .Q(\top_ihp.oisc.regs[47][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1352),
    .D(_01684_),
    .Q_N(_11796_),
    .Q(\top_ihp.oisc.regs[47][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1240),
    .D(_01685_),
    .Q_N(_11795_),
    .Q(\top_ihp.oisc.regs[47][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1389),
    .D(_01686_),
    .Q_N(_11794_),
    .Q(\top_ihp.oisc.regs[47][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1347),
    .D(_01687_),
    .Q_N(_11793_),
    .Q(\top_ihp.oisc.regs[47][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1359),
    .D(_01688_),
    .Q_N(_11792_),
    .Q(\top_ihp.oisc.regs[47][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1390),
    .D(_01689_),
    .Q_N(_11791_),
    .Q(\top_ihp.oisc.regs[47][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1384),
    .D(_01690_),
    .Q_N(_11790_),
    .Q(\top_ihp.oisc.regs[47][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1374),
    .D(_01691_),
    .Q_N(_11789_),
    .Q(\top_ihp.oisc.regs[47][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1339),
    .D(_01692_),
    .Q_N(_11788_),
    .Q(\top_ihp.oisc.regs[47][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1371),
    .D(_01693_),
    .Q_N(_11787_),
    .Q(\top_ihp.oisc.regs[47][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1297),
    .D(_01694_),
    .Q_N(_11786_),
    .Q(\top_ihp.oisc.regs[47][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1292),
    .D(_01695_),
    .Q_N(_11785_),
    .Q(\top_ihp.oisc.regs[47][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1326),
    .D(_01696_),
    .Q_N(_11784_),
    .Q(\top_ihp.oisc.regs[47][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1314),
    .D(_01697_),
    .Q_N(_11783_),
    .Q(\top_ihp.oisc.regs[47][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1309),
    .D(_01698_),
    .Q_N(_11782_),
    .Q(\top_ihp.oisc.regs[47][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1307),
    .D(_01699_),
    .Q_N(_11781_),
    .Q(\top_ihp.oisc.regs[47][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1301),
    .D(_01700_),
    .Q_N(_11780_),
    .Q(\top_ihp.oisc.regs[47][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1294),
    .D(_01701_),
    .Q_N(_11779_),
    .Q(\top_ihp.oisc.regs[47][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1258),
    .D(_01702_),
    .Q_N(_11778_),
    .Q(\top_ihp.oisc.regs[48][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1280),
    .D(_01703_),
    .Q_N(_11777_),
    .Q(\top_ihp.oisc.regs[48][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1274),
    .D(_01704_),
    .Q_N(_11776_),
    .Q(\top_ihp.oisc.regs[48][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1272),
    .D(_01705_),
    .Q_N(_11775_),
    .Q(\top_ihp.oisc.regs[48][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1247),
    .D(_01706_),
    .Q_N(_11774_),
    .Q(\top_ihp.oisc.regs[48][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1272),
    .D(_01707_),
    .Q_N(_11773_),
    .Q(\top_ihp.oisc.regs[48][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1192),
    .D(_01708_),
    .Q_N(_11772_),
    .Q(\top_ihp.oisc.regs[48][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1247),
    .D(_01709_),
    .Q_N(_11771_),
    .Q(\top_ihp.oisc.regs[48][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1199),
    .D(_01710_),
    .Q_N(_11770_),
    .Q(\top_ihp.oisc.regs[48][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1251),
    .D(_01711_),
    .Q_N(_11769_),
    .Q(\top_ihp.oisc.regs[48][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1211),
    .D(_01712_),
    .Q_N(_11768_),
    .Q(\top_ihp.oisc.regs[48][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1249),
    .D(_01713_),
    .Q_N(_11767_),
    .Q(\top_ihp.oisc.regs[48][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1258),
    .D(_01714_),
    .Q_N(_11766_),
    .Q(\top_ihp.oisc.regs[48][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1253),
    .D(_01715_),
    .Q_N(_11765_),
    .Q(\top_ihp.oisc.regs[48][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1351),
    .D(_01716_),
    .Q_N(_11764_),
    .Q(\top_ihp.oisc.regs[48][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1266),
    .D(_01717_),
    .Q_N(_11763_),
    .Q(\top_ihp.oisc.regs[48][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1384),
    .D(_01718_),
    .Q_N(_11762_),
    .Q(\top_ihp.oisc.regs[48][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1378),
    .D(_01719_),
    .Q_N(_11761_),
    .Q(\top_ihp.oisc.regs[48][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1383),
    .D(_01720_),
    .Q_N(_11760_),
    .Q(\top_ihp.oisc.regs[48][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1383),
    .D(_01721_),
    .Q_N(_11759_),
    .Q(\top_ihp.oisc.regs[48][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1368),
    .D(_01722_),
    .Q_N(_11758_),
    .Q(\top_ihp.oisc.regs[48][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1367),
    .D(_01723_),
    .Q_N(_11757_),
    .Q(\top_ihp.oisc.regs[48][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1365),
    .D(_01724_),
    .Q_N(_11756_),
    .Q(\top_ihp.oisc.regs[48][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1364),
    .D(_01725_),
    .Q_N(_11755_),
    .Q(\top_ihp.oisc.regs[48][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1325),
    .D(_01726_),
    .Q_N(_11754_),
    .Q(\top_ihp.oisc.regs[48][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1323),
    .D(_01727_),
    .Q_N(_11753_),
    .Q(\top_ihp.oisc.regs[48][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1303),
    .D(_01728_),
    .Q_N(_11752_),
    .Q(\top_ihp.oisc.regs[48][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1308),
    .D(_01729_),
    .Q_N(_11751_),
    .Q(\top_ihp.oisc.regs[48][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1303),
    .D(_01730_),
    .Q_N(_11750_),
    .Q(\top_ihp.oisc.regs[48][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1303),
    .D(_01731_),
    .Q_N(_11749_),
    .Q(\top_ihp.oisc.regs[48][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1302),
    .D(_01732_),
    .Q_N(_11748_),
    .Q(\top_ihp.oisc.regs[48][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1285),
    .D(_01733_),
    .Q_N(_11747_),
    .Q(\top_ihp.oisc.regs[48][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1264),
    .D(_01734_),
    .Q_N(_11746_),
    .Q(\top_ihp.oisc.regs[49][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1280),
    .D(_01735_),
    .Q_N(_11745_),
    .Q(\top_ihp.oisc.regs[49][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1201),
    .D(_01736_),
    .Q_N(_11744_),
    .Q(\top_ihp.oisc.regs[49][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1201),
    .D(_01737_),
    .Q_N(_11743_),
    .Q(\top_ihp.oisc.regs[49][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1221),
    .D(_01738_),
    .Q_N(_11742_),
    .Q(\top_ihp.oisc.regs[49][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1278),
    .D(_01739_),
    .Q_N(_11741_),
    .Q(\top_ihp.oisc.regs[49][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1199),
    .D(_01740_),
    .Q_N(_11740_),
    .Q(\top_ihp.oisc.regs[49][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1249),
    .D(_01741_),
    .Q_N(_11739_),
    .Q(\top_ihp.oisc.regs[49][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1207),
    .D(_01742_),
    .Q_N(_11738_),
    .Q(\top_ihp.oisc.regs[49][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1219),
    .D(_01743_),
    .Q_N(_11737_),
    .Q(\top_ihp.oisc.regs[49][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1215),
    .D(_01744_),
    .Q_N(_11736_),
    .Q(\top_ihp.oisc.regs[49][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1292),
    .D(_01745_),
    .Q_N(_11735_),
    .Q(\top_ihp.oisc.regs[49][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1267),
    .D(_01746_),
    .Q_N(_11734_),
    .Q(\top_ihp.oisc.regs[49][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1366),
    .D(_01747_),
    .Q_N(_11733_),
    .Q(\top_ihp.oisc.regs[49][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1357),
    .D(_01748_),
    .Q_N(_11732_),
    .Q(\top_ihp.oisc.regs[49][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1267),
    .D(_01749_),
    .Q_N(_11731_),
    .Q(\top_ihp.oisc.regs[49][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1389),
    .D(_01750_),
    .Q_N(_11730_),
    .Q(\top_ihp.oisc.regs[49][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1347),
    .D(_01751_),
    .Q_N(_11729_),
    .Q(\top_ihp.oisc.regs[49][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1359),
    .D(_01752_),
    .Q_N(_11728_),
    .Q(\top_ihp.oisc.regs[49][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1383),
    .D(_01753_),
    .Q_N(_11727_),
    .Q(\top_ihp.oisc.regs[49][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1390),
    .D(_01754_),
    .Q_N(_11726_),
    .Q(\top_ihp.oisc.regs[49][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1373),
    .D(_01755_),
    .Q_N(_11725_),
    .Q(\top_ihp.oisc.regs[49][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1339),
    .D(_01756_),
    .Q_N(_11724_),
    .Q(\top_ihp.oisc.regs[49][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1339),
    .D(_01757_),
    .Q_N(_11723_),
    .Q(\top_ihp.oisc.regs[49][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1323),
    .D(_01758_),
    .Q_N(_11722_),
    .Q(\top_ihp.oisc.regs[49][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1329),
    .D(_01759_),
    .Q_N(_11721_),
    .Q(\top_ihp.oisc.regs[49][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1309),
    .D(_01760_),
    .Q_N(_11720_),
    .Q(\top_ihp.oisc.regs[49][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1314),
    .D(_01761_),
    .Q_N(_11719_),
    .Q(\top_ihp.oisc.regs[49][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1309),
    .D(_01762_),
    .Q_N(_11718_),
    .Q(\top_ihp.oisc.regs[49][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1309),
    .D(_01763_),
    .Q_N(_11717_),
    .Q(\top_ihp.oisc.regs[49][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1301),
    .D(_01764_),
    .Q_N(_11716_),
    .Q(\top_ihp.oisc.regs[49][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1281),
    .D(_01765_),
    .Q_N(_11715_),
    .Q(\top_ihp.oisc.regs[49][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1164),
    .D(_01766_),
    .Q_N(_11714_),
    .Q(\top_ihp.oisc.regs[4][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1175),
    .D(_01767_),
    .Q_N(_11713_),
    .Q(\top_ihp.oisc.regs[4][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1175),
    .D(_01768_),
    .Q_N(_11712_),
    .Q(\top_ihp.oisc.regs[4][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1175),
    .D(_01769_),
    .Q_N(_11711_),
    .Q(\top_ihp.oisc.regs[4][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1229),
    .D(_01770_),
    .Q_N(_11710_),
    .Q(\top_ihp.oisc.regs[4][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1177),
    .D(_01771_),
    .Q_N(_11709_),
    .Q(\top_ihp.oisc.regs[4][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1191),
    .D(_01772_),
    .Q_N(_11708_),
    .Q(\top_ihp.oisc.regs[4][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1229),
    .D(_01773_),
    .Q_N(_11707_),
    .Q(\top_ihp.oisc.regs[4][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1209),
    .D(_01774_),
    .Q_N(_11706_),
    .Q(\top_ihp.oisc.regs[4][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1189),
    .D(_01775_),
    .Q_N(_11705_),
    .Q(\top_ihp.oisc.regs[4][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1209),
    .D(_01776_),
    .Q_N(_11704_),
    .Q(\top_ihp.oisc.regs[4][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1246),
    .D(_01777_),
    .Q_N(_11703_),
    .Q(\top_ihp.oisc.regs[4][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1164),
    .D(_01778_),
    .Q_N(_11702_),
    .Q(\top_ihp.oisc.regs[4][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1230),
    .D(_01779_),
    .Q_N(_11701_),
    .Q(\top_ihp.oisc.regs[4][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1237),
    .D(_01780_),
    .Q_N(_11700_),
    .Q(\top_ihp.oisc.regs[4][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1164),
    .D(_01781_),
    .Q_N(_11699_),
    .Q(\top_ihp.oisc.regs[4][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1237),
    .D(_01782_),
    .Q_N(_11698_),
    .Q(\top_ihp.oisc.regs[4][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1237),
    .D(_01783_),
    .Q_N(_11697_),
    .Q(\top_ihp.oisc.regs[4][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1232),
    .D(_01784_),
    .Q_N(_11696_),
    .Q(\top_ihp.oisc.regs[4][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1242),
    .D(_01785_),
    .Q_N(_11695_),
    .Q(\top_ihp.oisc.regs[4][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1242),
    .D(_01786_),
    .Q_N(_11694_),
    .Q(\top_ihp.oisc.regs[4][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1230),
    .D(_01787_),
    .Q_N(_11693_),
    .Q(\top_ihp.oisc.regs[4][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1230),
    .D(_01788_),
    .Q_N(_11692_),
    .Q(\top_ihp.oisc.regs[4][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1229),
    .D(_01789_),
    .Q_N(_11691_),
    .Q(\top_ihp.oisc.regs[4][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1213),
    .D(_01790_),
    .Q_N(_11690_),
    .Q(\top_ihp.oisc.regs[4][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1189),
    .D(_01791_),
    .Q_N(_11689_),
    .Q(\top_ihp.oisc.regs[4][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1185),
    .D(_01792_),
    .Q_N(_11688_),
    .Q(\top_ihp.oisc.regs[4][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1185),
    .D(_01793_),
    .Q_N(_11687_),
    .Q(\top_ihp.oisc.regs[4][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1174),
    .D(_01794_),
    .Q_N(_11686_),
    .Q(\top_ihp.oisc.regs[4][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1174),
    .D(_01795_),
    .Q_N(_11685_),
    .Q(\top_ihp.oisc.regs[4][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1175),
    .D(_01796_),
    .Q_N(_11684_),
    .Q(\top_ihp.oisc.regs[4][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1175),
    .D(_01797_),
    .Q_N(_11683_),
    .Q(\top_ihp.oisc.regs[4][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1349),
    .D(_01798_),
    .Q_N(_11682_),
    .Q(\top_ihp.oisc.regs[50][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1280),
    .D(_01799_),
    .Q_N(_11681_),
    .Q(\top_ihp.oisc.regs[50][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1274),
    .D(_01800_),
    .Q_N(_11680_),
    .Q(\top_ihp.oisc.regs[50][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1192),
    .D(_01801_),
    .Q_N(_11679_),
    .Q(\top_ihp.oisc.regs[50][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1214),
    .D(_01802_),
    .Q_N(_11678_),
    .Q(\top_ihp.oisc.regs[50][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1201),
    .D(_01803_),
    .Q_N(_11677_),
    .Q(\top_ihp.oisc.regs[50][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1192),
    .D(_01804_),
    .Q_N(_11676_),
    .Q(\top_ihp.oisc.regs[50][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1214),
    .D(_01805_),
    .Q_N(_11675_),
    .Q(\top_ihp.oisc.regs[50][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1200),
    .D(_01806_),
    .Q_N(_11674_),
    .Q(\top_ihp.oisc.regs[50][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1212),
    .D(_01807_),
    .Q_N(_11673_),
    .Q(\top_ihp.oisc.regs[50][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1215),
    .D(_01808_),
    .Q_N(_11672_),
    .Q(\top_ihp.oisc.regs[50][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1292),
    .D(_01809_),
    .Q_N(_11671_),
    .Q(\top_ihp.oisc.regs[50][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1349),
    .D(_01810_),
    .Q_N(_11670_),
    .Q(\top_ihp.oisc.regs[50][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1369),
    .D(_01811_),
    .Q_N(_11669_),
    .Q(\top_ihp.oisc.regs[50][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1353),
    .D(_01812_),
    .Q_N(_11668_),
    .Q(\top_ihp.oisc.regs[50][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1267),
    .D(_01813_),
    .Q_N(_11667_),
    .Q(\top_ihp.oisc.regs[50][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1387),
    .D(_01814_),
    .Q_N(_11666_),
    .Q(\top_ihp.oisc.regs[50][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1378),
    .D(_01815_),
    .Q_N(_11665_),
    .Q(\top_ihp.oisc.regs[50][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1369),
    .D(_01816_),
    .Q_N(_11664_),
    .Q(\top_ihp.oisc.regs[50][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1387),
    .D(_01817_),
    .Q_N(_11663_),
    .Q(\top_ihp.oisc.regs[50][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1375),
    .D(_01818_),
    .Q_N(_11662_),
    .Q(\top_ihp.oisc.regs[50][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1341),
    .D(_01819_),
    .Q_N(_11661_),
    .Q(\top_ihp.oisc.regs[50][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1370),
    .D(_01820_),
    .Q_N(_11660_),
    .Q(\top_ihp.oisc.regs[50][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1371),
    .D(_01821_),
    .Q_N(_11659_),
    .Q(\top_ihp.oisc.regs[50][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1331),
    .D(_01822_),
    .Q_N(_11658_),
    .Q(\top_ihp.oisc.regs[50][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1323),
    .D(_01823_),
    .Q_N(_11657_),
    .Q(\top_ihp.oisc.regs[50][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1320),
    .D(_01824_),
    .Q_N(_11656_),
    .Q(\top_ihp.oisc.regs[50][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1294),
    .D(_01825_),
    .Q_N(_11655_),
    .Q(\top_ihp.oisc.regs[50][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1311),
    .D(_01826_),
    .Q_N(_11654_),
    .Q(\top_ihp.oisc.regs[50][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1315),
    .D(_01827_),
    .Q_N(_11653_),
    .Q(\top_ihp.oisc.regs[50][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1301),
    .D(_01828_),
    .Q_N(_11652_),
    .Q(\top_ihp.oisc.regs[50][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1281),
    .D(_01829_),
    .Q_N(_11651_),
    .Q(\top_ihp.oisc.regs[50][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1257),
    .D(_01830_),
    .Q_N(_11650_),
    .Q(\top_ihp.oisc.regs[51][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1281),
    .D(_01831_),
    .Q_N(_11649_),
    .Q(\top_ihp.oisc.regs[51][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1201),
    .D(_01832_),
    .Q_N(_11648_),
    .Q(\top_ihp.oisc.regs[51][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1191),
    .D(_01833_),
    .Q_N(_11647_),
    .Q(\top_ihp.oisc.regs[51][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1250),
    .D(_01834_),
    .Q_N(_11646_),
    .Q(\top_ihp.oisc.regs[51][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1195),
    .D(_01835_),
    .Q_N(_11645_),
    .Q(\top_ihp.oisc.regs[51][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1191),
    .D(_01836_),
    .Q_N(_11644_),
    .Q(\top_ihp.oisc.regs[51][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1245),
    .D(_01837_),
    .Q_N(_11643_),
    .Q(\top_ihp.oisc.regs[51][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1192),
    .D(_01838_),
    .Q_N(_11642_),
    .Q(\top_ihp.oisc.regs[51][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1213),
    .D(_01839_),
    .Q_N(_11641_),
    .Q(\top_ihp.oisc.regs[51][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1209),
    .D(_01840_),
    .Q_N(_11640_),
    .Q(\top_ihp.oisc.regs[51][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1335),
    .D(_01841_),
    .Q_N(_11639_),
    .Q(\top_ihp.oisc.regs[51][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1257),
    .D(_01842_),
    .Q_N(_11638_),
    .Q(\top_ihp.oisc.regs[51][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1342),
    .D(_01843_),
    .Q_N(_11637_),
    .Q(\top_ihp.oisc.regs[51][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1355),
    .D(_01844_),
    .Q_N(_11636_),
    .Q(\top_ihp.oisc.regs[51][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1256),
    .D(_01845_),
    .Q_N(_11635_),
    .Q(\top_ihp.oisc.regs[51][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1387),
    .D(_01846_),
    .Q_N(_11634_),
    .Q(\top_ihp.oisc.regs[51][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1378),
    .D(_01847_),
    .Q_N(_11633_),
    .Q(\top_ihp.oisc.regs[51][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1368),
    .D(_01848_),
    .Q_N(_11632_),
    .Q(\top_ihp.oisc.regs[51][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1387),
    .D(_01849_),
    .Q_N(_11631_),
    .Q(\top_ihp.oisc.regs[51][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1388),
    .D(_01850_),
    .Q_N(_11630_),
    .Q(\top_ihp.oisc.regs[51][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1374),
    .D(_01851_),
    .Q_N(_11629_),
    .Q(\top_ihp.oisc.regs[51][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1340),
    .D(_01852_),
    .Q_N(_11628_),
    .Q(\top_ihp.oisc.regs[51][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1372),
    .D(_01853_),
    .Q_N(_11627_),
    .Q(\top_ihp.oisc.regs[51][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1330),
    .D(_01854_),
    .Q_N(_11626_),
    .Q(\top_ihp.oisc.regs[51][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1330),
    .D(_01855_),
    .Q_N(_11625_),
    .Q(\top_ihp.oisc.regs[51][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1327),
    .D(_01856_),
    .Q_N(_11624_),
    .Q(\top_ihp.oisc.regs[51][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1315),
    .D(_01857_),
    .Q_N(_11623_),
    .Q(\top_ihp.oisc.regs[51][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1311),
    .D(_01858_),
    .Q_N(_11622_),
    .Q(\top_ihp.oisc.regs[51][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1312),
    .D(_01859_),
    .Q_N(_11621_),
    .Q(\top_ihp.oisc.regs[51][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1302),
    .D(_01860_),
    .Q_N(_11620_),
    .Q(\top_ihp.oisc.regs[51][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1285),
    .D(_01861_),
    .Q_N(_11619_),
    .Q(\top_ihp.oisc.regs[51][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1345),
    .D(_01862_),
    .Q_N(_11618_),
    .Q(\top_ihp.oisc.regs[52][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1281),
    .D(_01863_),
    .Q_N(_11617_),
    .Q(\top_ihp.oisc.regs[52][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1272),
    .D(_01864_),
    .Q_N(_11616_),
    .Q(\top_ihp.oisc.regs[52][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1201),
    .D(_01865_),
    .Q_N(_11615_),
    .Q(\top_ihp.oisc.regs[52][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1250),
    .D(_01866_),
    .Q_N(_11614_),
    .Q(\top_ihp.oisc.regs[52][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1192),
    .D(_01867_),
    .Q_N(_11613_),
    .Q(\top_ihp.oisc.regs[52][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1192),
    .D(_01868_),
    .Q_N(_11612_),
    .Q(\top_ihp.oisc.regs[52][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1244),
    .D(_01869_),
    .Q_N(_11611_),
    .Q(\top_ihp.oisc.regs[52][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1199),
    .D(_01870_),
    .Q_N(_11610_),
    .Q(\top_ihp.oisc.regs[52][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1251),
    .D(_01871_),
    .Q_N(_11609_),
    .Q(\top_ihp.oisc.regs[52][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1212),
    .D(_01872_),
    .Q_N(_11608_),
    .Q(\top_ihp.oisc.regs[52][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1335),
    .D(_01873_),
    .Q_N(_11607_),
    .Q(\top_ihp.oisc.regs[52][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1265),
    .D(_01874_),
    .Q_N(_11606_),
    .Q(\top_ihp.oisc.regs[52][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1342),
    .D(_01875_),
    .Q_N(_11605_),
    .Q(\top_ihp.oisc.regs[52][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1347),
    .D(_01876_),
    .Q_N(_11604_),
    .Q(\top_ihp.oisc.regs[52][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1265),
    .D(_01877_),
    .Q_N(_11603_),
    .Q(\top_ihp.oisc.regs[52][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1387),
    .D(_01878_),
    .Q_N(_11602_),
    .Q(\top_ihp.oisc.regs[52][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1345),
    .D(_01879_),
    .Q_N(_11601_),
    .Q(\top_ihp.oisc.regs[52][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1345),
    .D(_01880_),
    .Q_N(_11600_),
    .Q(\top_ihp.oisc.regs[52][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1387),
    .D(_01881_),
    .Q_N(_11599_),
    .Q(\top_ihp.oisc.regs[52][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1375),
    .D(_01882_),
    .Q_N(_11598_),
    .Q(\top_ihp.oisc.regs[52][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1338),
    .D(_01883_),
    .Q_N(_11597_),
    .Q(\top_ihp.oisc.regs[52][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1335),
    .D(_01884_),
    .Q_N(_11596_),
    .Q(\top_ihp.oisc.regs[52][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1371),
    .D(_01885_),
    .Q_N(_11595_),
    .Q(\top_ihp.oisc.regs[52][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1325),
    .D(_01886_),
    .Q_N(_11594_),
    .Q(\top_ihp.oisc.regs[52][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1296),
    .D(_01887_),
    .Q_N(_11593_),
    .Q(\top_ihp.oisc.regs[52][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1327),
    .D(_01888_),
    .Q_N(_11592_),
    .Q(\top_ihp.oisc.regs[52][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1311),
    .D(_01889_),
    .Q_N(_11591_),
    .Q(\top_ihp.oisc.regs[52][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1311),
    .D(_01890_),
    .Q_N(_11590_),
    .Q(\top_ihp.oisc.regs[52][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1280),
    .D(_01891_),
    .Q_N(_11589_),
    .Q(\top_ihp.oisc.regs[52][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1301),
    .D(_01892_),
    .Q_N(_11588_),
    .Q(\top_ihp.oisc.regs[52][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1293),
    .D(_01893_),
    .Q_N(_11587_),
    .Q(\top_ihp.oisc.regs[52][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1260),
    .D(_01894_),
    .Q_N(_11586_),
    .Q(\top_ihp.oisc.regs[53][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1281),
    .D(_01895_),
    .Q_N(_11585_),
    .Q(\top_ihp.oisc.regs[53][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1272),
    .D(_01896_),
    .Q_N(_11584_),
    .Q(\top_ihp.oisc.regs[53][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1274),
    .D(_01897_),
    .Q_N(_11583_),
    .Q(\top_ihp.oisc.regs[53][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1261),
    .D(_01898_),
    .Q_N(_11582_),
    .Q(\top_ihp.oisc.regs[53][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1272),
    .D(_01899_),
    .Q_N(_11581_),
    .Q(\top_ihp.oisc.regs[53][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1199),
    .D(_01900_),
    .Q_N(_11580_),
    .Q(\top_ihp.oisc.regs[53][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1261),
    .D(_01901_),
    .Q_N(_11579_),
    .Q(\top_ihp.oisc.regs[53][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1199),
    .D(_01902_),
    .Q_N(_11578_),
    .Q(\top_ihp.oisc.regs[53][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1221),
    .D(_01903_),
    .Q_N(_11577_),
    .Q(\top_ihp.oisc.regs[53][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1218),
    .D(_01904_),
    .Q_N(_11576_),
    .Q(\top_ihp.oisc.regs[53][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1290),
    .D(_01905_),
    .Q_N(_11575_),
    .Q(\top_ihp.oisc.regs[53][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1349),
    .D(_01906_),
    .Q_N(_11574_),
    .Q(\top_ihp.oisc.regs[53][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1342),
    .D(_01907_),
    .Q_N(_11573_),
    .Q(\top_ihp.oisc.regs[53][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1352),
    .D(_01908_),
    .Q_N(_11572_),
    .Q(\top_ihp.oisc.regs[53][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1266),
    .D(_01909_),
    .Q_N(_11571_),
    .Q(\top_ihp.oisc.regs[53][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1390),
    .D(_01910_),
    .Q_N(_11570_),
    .Q(\top_ihp.oisc.regs[53][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1381),
    .D(_01911_),
    .Q_N(_11569_),
    .Q(\top_ihp.oisc.regs[53][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1381),
    .D(_01912_),
    .Q_N(_11568_),
    .Q(\top_ihp.oisc.regs[53][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1390),
    .D(_01913_),
    .Q_N(_11567_),
    .Q(\top_ihp.oisc.regs[53][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1375),
    .D(_01914_),
    .Q_N(_11566_),
    .Q(\top_ihp.oisc.regs[53][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1366),
    .D(_01915_),
    .Q_N(_11565_),
    .Q(\top_ihp.oisc.regs[53][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1373),
    .D(_01916_),
    .Q_N(_11564_),
    .Q(\top_ihp.oisc.regs[53][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1363),
    .D(_01917_),
    .Q_N(_11563_),
    .Q(\top_ihp.oisc.regs[53][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1330),
    .D(_01918_),
    .Q_N(_11562_),
    .Q(\top_ihp.oisc.regs[53][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1329),
    .D(_01919_),
    .Q_N(_11561_),
    .Q(\top_ihp.oisc.regs[53][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1309),
    .D(_01920_),
    .Q_N(_11560_),
    .Q(\top_ihp.oisc.regs[53][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1311),
    .D(_01921_),
    .Q_N(_11559_),
    .Q(\top_ihp.oisc.regs[53][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1311),
    .D(_01922_),
    .Q_N(_11558_),
    .Q(\top_ihp.oisc.regs[53][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1281),
    .D(_01923_),
    .Q_N(_11557_),
    .Q(\top_ihp.oisc.regs[53][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1301),
    .D(_01924_),
    .Q_N(_11556_),
    .Q(\top_ihp.oisc.regs[53][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1281),
    .D(_01925_),
    .Q_N(_11555_),
    .Q(\top_ihp.oisc.regs[53][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1256),
    .D(_01926_),
    .Q_N(_11554_),
    .Q(\top_ihp.oisc.regs[54][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1280),
    .D(_01927_),
    .Q_N(_11553_),
    .Q(\top_ihp.oisc.regs[54][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1272),
    .D(_01928_),
    .Q_N(_11552_),
    .Q(\top_ihp.oisc.regs[54][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1293),
    .D(_01929_),
    .Q_N(_11551_),
    .Q(\top_ihp.oisc.regs[54][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1244),
    .D(_01930_),
    .Q_N(_11550_),
    .Q(\top_ihp.oisc.regs[54][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1191),
    .D(_01931_),
    .Q_N(_11549_),
    .Q(\top_ihp.oisc.regs[54][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1191),
    .D(_01932_),
    .Q_N(_11548_),
    .Q(\top_ihp.oisc.regs[54][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1257),
    .D(_01933_),
    .Q_N(_11547_),
    .Q(\top_ihp.oisc.regs[54][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1216),
    .D(_01934_),
    .Q_N(_11546_),
    .Q(\top_ihp.oisc.regs[54][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1291),
    .D(_01935_),
    .Q_N(_11545_),
    .Q(\top_ihp.oisc.regs[54][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1210),
    .D(_01936_),
    .Q_N(_11544_),
    .Q(\top_ihp.oisc.regs[54][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1339),
    .D(_01937_),
    .Q_N(_11543_),
    .Q(\top_ihp.oisc.regs[54][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1256),
    .D(_01938_),
    .Q_N(_11542_),
    .Q(\top_ihp.oisc.regs[54][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1253),
    .D(_01939_),
    .Q_N(_11541_),
    .Q(\top_ihp.oisc.regs[54][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1347),
    .D(_01940_),
    .Q_N(_11540_),
    .Q(\top_ihp.oisc.regs[54][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1264),
    .D(_01941_),
    .Q_N(_11539_),
    .Q(\top_ihp.oisc.regs[54][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1354),
    .D(_01942_),
    .Q_N(_11538_),
    .Q(\top_ihp.oisc.regs[54][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1336),
    .D(_01943_),
    .Q_N(_11537_),
    .Q(\top_ihp.oisc.regs[54][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1338),
    .D(_01944_),
    .Q_N(_11536_),
    .Q(\top_ihp.oisc.regs[54][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1373),
    .D(_01945_),
    .Q_N(_11535_),
    .Q(\top_ihp.oisc.regs[54][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1386),
    .D(_01946_),
    .Q_N(_11534_),
    .Q(\top_ihp.oisc.regs[54][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1376),
    .D(_01947_),
    .Q_N(_11533_),
    .Q(\top_ihp.oisc.regs[54][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1366),
    .D(_01948_),
    .Q_N(_11532_),
    .Q(\top_ihp.oisc.regs[54][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1364),
    .D(_01949_),
    .Q_N(_11531_),
    .Q(\top_ihp.oisc.regs[54][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1325),
    .D(_01950_),
    .Q_N(_11530_),
    .Q(\top_ihp.oisc.regs[54][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1325),
    .D(_01951_),
    .Q_N(_11529_),
    .Q(\top_ihp.oisc.regs[54][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1295),
    .D(_01952_),
    .Q_N(_11528_),
    .Q(\top_ihp.oisc.regs[54][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1317),
    .D(_01953_),
    .Q_N(_11527_),
    .Q(\top_ihp.oisc.regs[54][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1310),
    .D(_01954_),
    .Q_N(_11526_),
    .Q(\top_ihp.oisc.regs[54][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1317),
    .D(_01955_),
    .Q_N(_11525_),
    .Q(\top_ihp.oisc.regs[54][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1308),
    .D(_01956_),
    .Q_N(_11524_),
    .Q(\top_ihp.oisc.regs[54][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1295),
    .D(_01957_),
    .Q_N(_11523_),
    .Q(\top_ihp.oisc.regs[54][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1260),
    .D(_01958_),
    .Q_N(_11522_),
    .Q(\top_ihp.oisc.regs[55][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1283),
    .D(_01959_),
    .Q_N(_11521_),
    .Q(\top_ihp.oisc.regs[55][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1273),
    .D(_01960_),
    .Q_N(_11520_),
    .Q(\top_ihp.oisc.regs[55][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1278),
    .D(_01961_),
    .Q_N(_11519_),
    .Q(\top_ihp.oisc.regs[55][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1252),
    .D(_01962_),
    .Q_N(_11518_),
    .Q(\top_ihp.oisc.regs[55][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1289),
    .D(_01963_),
    .Q_N(_11517_),
    .Q(\top_ihp.oisc.regs[55][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1216),
    .D(_01964_),
    .Q_N(_11516_),
    .Q(\top_ihp.oisc.regs[55][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1260),
    .D(_01965_),
    .Q_N(_11515_),
    .Q(\top_ihp.oisc.regs[55][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1205),
    .D(_01966_),
    .Q_N(_11514_),
    .Q(\top_ihp.oisc.regs[55][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1251),
    .D(_01967_),
    .Q_N(_11513_),
    .Q(\top_ihp.oisc.regs[55][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1220),
    .D(_01968_),
    .Q_N(_11512_),
    .Q(\top_ihp.oisc.regs[55][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1292),
    .D(_01969_),
    .Q_N(_11511_),
    .Q(\top_ihp.oisc.regs[55][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1267),
    .D(_01970_),
    .Q_N(_11510_),
    .Q(\top_ihp.oisc.regs[55][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1341),
    .D(_01971_),
    .Q_N(_11509_),
    .Q(\top_ihp.oisc.regs[55][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1357),
    .D(_01972_),
    .Q_N(_11508_),
    .Q(\top_ihp.oisc.regs[55][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1256),
    .D(_01973_),
    .Q_N(_11507_),
    .Q(\top_ihp.oisc.regs[55][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1343),
    .D(_01974_),
    .Q_N(_11506_),
    .Q(\top_ihp.oisc.regs[55][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1337),
    .D(_01975_),
    .Q_N(_11505_),
    .Q(\top_ihp.oisc.regs[55][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1366),
    .D(_01976_),
    .Q_N(_11504_),
    .Q(\top_ihp.oisc.regs[55][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1368),
    .D(_01977_),
    .Q_N(_11503_),
    .Q(\top_ihp.oisc.regs[55][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1374),
    .D(_01978_),
    .Q_N(_11502_),
    .Q(\top_ihp.oisc.regs[55][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1337),
    .D(_01979_),
    .Q_N(_11501_),
    .Q(\top_ihp.oisc.regs[55][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1335),
    .D(_01980_),
    .Q_N(_11500_),
    .Q(\top_ihp.oisc.regs[55][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1371),
    .D(_01981_),
    .Q_N(_11499_),
    .Q(\top_ihp.oisc.regs[55][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1325),
    .D(_01982_),
    .Q_N(_11498_),
    .Q(\top_ihp.oisc.regs[55][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1331),
    .D(_01983_),
    .Q_N(_11497_),
    .Q(\top_ihp.oisc.regs[55][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1319),
    .D(_01984_),
    .Q_N(_11496_),
    .Q(\top_ihp.oisc.regs[55][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1288),
    .D(_01985_),
    .Q_N(_11495_),
    .Q(\top_ihp.oisc.regs[55][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1315),
    .D(_01986_),
    .Q_N(_11494_),
    .Q(\top_ihp.oisc.regs[55][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1315),
    .D(_01987_),
    .Q_N(_11493_),
    .Q(\top_ihp.oisc.regs[55][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1319),
    .D(_01988_),
    .Q_N(_11492_),
    .Q(\top_ihp.oisc.regs[55][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1293),
    .D(_01989_),
    .Q_N(_11491_),
    .Q(\top_ihp.oisc.regs[55][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1351),
    .D(_01990_),
    .Q_N(_11490_),
    .Q(\top_ihp.oisc.regs[56][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1284),
    .D(_01991_),
    .Q_N(_11489_),
    .Q(\top_ihp.oisc.regs[56][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1205),
    .D(_01992_),
    .Q_N(_11488_),
    .Q(\top_ihp.oisc.regs[56][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1204),
    .D(_01993_),
    .Q_N(_11487_),
    .Q(\top_ihp.oisc.regs[56][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1252),
    .D(_01994_),
    .Q_N(_11486_),
    .Q(\top_ihp.oisc.regs[56][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1288),
    .D(_01995_),
    .Q_N(_11485_),
    .Q(\top_ihp.oisc.regs[56][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1206),
    .D(_01996_),
    .Q_N(_11484_),
    .Q(\top_ihp.oisc.regs[56][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1260),
    .D(_01997_),
    .Q_N(_11483_),
    .Q(\top_ihp.oisc.regs[56][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1205),
    .D(_01998_),
    .Q_N(_11482_),
    .Q(\top_ihp.oisc.regs[56][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1290),
    .D(_01999_),
    .Q_N(_11481_),
    .Q(\top_ihp.oisc.regs[56][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1217),
    .D(_02000_),
    .Q_N(_11480_),
    .Q(\top_ihp.oisc.regs[56][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1296),
    .D(_02001_),
    .Q_N(_11479_),
    .Q(\top_ihp.oisc.regs[56][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1265),
    .D(_02002_),
    .Q_N(_11478_),
    .Q(\top_ihp.oisc.regs[56][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1253),
    .D(_02003_),
    .Q_N(_11477_),
    .Q(\top_ihp.oisc.regs[56][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1351),
    .D(_02004_),
    .Q_N(_11476_),
    .Q(\top_ihp.oisc.regs[56][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1264),
    .D(_02005_),
    .Q_N(_11475_),
    .Q(\top_ihp.oisc.regs[56][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1253),
    .D(_02006_),
    .Q_N(_11474_),
    .Q(\top_ihp.oisc.regs[56][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1341),
    .D(_02007_),
    .Q_N(_11473_),
    .Q(\top_ihp.oisc.regs[56][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1354),
    .D(_02008_),
    .Q_N(_11472_),
    .Q(\top_ihp.oisc.regs[56][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1368),
    .D(_02009_),
    .Q_N(_11471_),
    .Q(\top_ihp.oisc.regs[56][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1386),
    .D(_02010_),
    .Q_N(_11470_),
    .Q(\top_ihp.oisc.regs[56][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1341),
    .D(_02011_),
    .Q_N(_11469_),
    .Q(\top_ihp.oisc.regs[56][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1365),
    .D(_02012_),
    .Q_N(_11468_),
    .Q(\top_ihp.oisc.regs[56][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1370),
    .D(_02013_),
    .Q_N(_11467_),
    .Q(\top_ihp.oisc.regs[56][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1323),
    .D(_02014_),
    .Q_N(_11466_),
    .Q(\top_ihp.oisc.regs[56][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1329),
    .D(_02015_),
    .Q_N(_11465_),
    .Q(\top_ihp.oisc.regs[56][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1320),
    .D(_02016_),
    .Q_N(_11464_),
    .Q(\top_ihp.oisc.regs[56][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1321),
    .D(_02017_),
    .Q_N(_11463_),
    .Q(\top_ihp.oisc.regs[56][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1307),
    .D(_02018_),
    .Q_N(_11462_),
    .Q(\top_ihp.oisc.regs[56][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1314),
    .D(_02019_),
    .Q_N(_11461_),
    .Q(\top_ihp.oisc.regs[56][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1308),
    .D(_02020_),
    .Q_N(_11460_),
    .Q(\top_ihp.oisc.regs[56][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1285),
    .D(_02021_),
    .Q_N(_11459_),
    .Q(\top_ihp.oisc.regs[56][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1346),
    .D(_02022_),
    .Q_N(_11458_),
    .Q(\top_ihp.oisc.regs[57][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1284),
    .D(_02023_),
    .Q_N(_11457_),
    .Q(\top_ihp.oisc.regs[57][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1206),
    .D(_02024_),
    .Q_N(_11456_),
    .Q(\top_ihp.oisc.regs[57][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1277),
    .D(_02025_),
    .Q_N(_11455_),
    .Q(\top_ihp.oisc.regs[57][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1221),
    .D(_02026_),
    .Q_N(_11454_),
    .Q(\top_ihp.oisc.regs[57][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1289),
    .D(_02027_),
    .Q_N(_11453_),
    .Q(\top_ihp.oisc.regs[57][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1216),
    .D(_02028_),
    .Q_N(_11452_),
    .Q(\top_ihp.oisc.regs[57][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1249),
    .D(_02029_),
    .Q_N(_11451_),
    .Q(\top_ihp.oisc.regs[57][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1215),
    .D(_02030_),
    .Q_N(_11450_),
    .Q(\top_ihp.oisc.regs[57][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1290),
    .D(_02031_),
    .Q_N(_11449_),
    .Q(\top_ihp.oisc.regs[57][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1218),
    .D(_02032_),
    .Q_N(_11448_),
    .Q(\top_ihp.oisc.regs[57][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1296),
    .D(_02033_),
    .Q_N(_11447_),
    .Q(\top_ihp.oisc.regs[57][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1265),
    .D(_02034_),
    .Q_N(_11446_),
    .Q(\top_ihp.oisc.regs[57][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1343),
    .D(_02035_),
    .Q_N(_11445_),
    .Q(\top_ihp.oisc.regs[57][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1353),
    .D(_02036_),
    .Q_N(_11444_),
    .Q(\top_ihp.oisc.regs[57][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1270),
    .D(_02037_),
    .Q_N(_11443_),
    .Q(\top_ihp.oisc.regs[57][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1388),
    .D(_02038_),
    .Q_N(_11442_),
    .Q(\top_ihp.oisc.regs[57][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1355),
    .D(_02039_),
    .Q_N(_11441_),
    .Q(\top_ihp.oisc.regs[57][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1381),
    .D(_02040_),
    .Q_N(_11440_),
    .Q(\top_ihp.oisc.regs[57][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1388),
    .D(_02041_),
    .Q_N(_11439_),
    .Q(\top_ihp.oisc.regs[57][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1390),
    .D(_02042_),
    .Q_N(_11438_),
    .Q(\top_ihp.oisc.regs[57][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1339),
    .D(_02043_),
    .Q_N(_11437_),
    .Q(\top_ihp.oisc.regs[57][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1373),
    .D(_02044_),
    .Q_N(_11436_),
    .Q(\top_ihp.oisc.regs[57][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1371),
    .D(_02045_),
    .Q_N(_11435_),
    .Q(\top_ihp.oisc.regs[57][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1331),
    .D(_02046_),
    .Q_N(_11434_),
    .Q(\top_ihp.oisc.regs[57][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1330),
    .D(_02047_),
    .Q_N(_11433_),
    .Q(\top_ihp.oisc.regs[57][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1327),
    .D(_02048_),
    .Q_N(_11432_),
    .Q(\top_ihp.oisc.regs[57][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1316),
    .D(_02049_),
    .Q_N(_11431_),
    .Q(\top_ihp.oisc.regs[57][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1315),
    .D(_02050_),
    .Q_N(_11430_),
    .Q(\top_ihp.oisc.regs[57][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1316),
    .D(_02051_),
    .Q_N(_11429_),
    .Q(\top_ihp.oisc.regs[57][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1294),
    .D(_02052_),
    .Q_N(_11428_),
    .Q(\top_ihp.oisc.regs[57][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1294),
    .D(_02053_),
    .Q_N(_11427_),
    .Q(\top_ihp.oisc.regs[57][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1263),
    .D(_02054_),
    .Q_N(_11426_),
    .Q(\top_ihp.oisc.regs[58][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1283),
    .D(_02055_),
    .Q_N(_11425_),
    .Q(\top_ihp.oisc.regs[58][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1205),
    .D(_02056_),
    .Q_N(_11424_),
    .Q(\top_ihp.oisc.regs[58][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1204),
    .D(_02057_),
    .Q_N(_11423_),
    .Q(\top_ihp.oisc.regs[58][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1249),
    .D(_02058_),
    .Q_N(_11422_),
    .Q(\top_ihp.oisc.regs[58][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1195),
    .D(_02059_),
    .Q_N(_11421_),
    .Q(\top_ihp.oisc.regs[58][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1209),
    .D(_02060_),
    .Q_N(_11420_),
    .Q(\top_ihp.oisc.regs[58][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1244),
    .D(_02061_),
    .Q_N(_11419_),
    .Q(\top_ihp.oisc.regs[58][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1195),
    .D(_02062_),
    .Q_N(_11418_),
    .Q(\top_ihp.oisc.regs[58][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1291),
    .D(_02063_),
    .Q_N(_11417_),
    .Q(\top_ihp.oisc.regs[58][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1210),
    .D(_02064_),
    .Q_N(_11416_),
    .Q(\top_ihp.oisc.regs[58][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1298),
    .D(_02065_),
    .Q_N(_11415_),
    .Q(\top_ihp.oisc.regs[58][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1256),
    .D(_02066_),
    .Q_N(_11414_),
    .Q(\top_ihp.oisc.regs[58][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1353),
    .D(_02067_),
    .Q_N(_11413_),
    .Q(\top_ihp.oisc.regs[58][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1356),
    .D(_02068_),
    .Q_N(_11412_),
    .Q(\top_ihp.oisc.regs[58][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1263),
    .D(_02069_),
    .Q_N(_11411_),
    .Q(\top_ihp.oisc.regs[58][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1386),
    .D(_02070_),
    .Q_N(_11410_),
    .Q(\top_ihp.oisc.regs[58][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1341),
    .D(_02071_),
    .Q_N(_11409_),
    .Q(\top_ihp.oisc.regs[58][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1369),
    .D(_02072_),
    .Q_N(_11408_),
    .Q(\top_ihp.oisc.regs[58][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1376),
    .D(_02073_),
    .Q_N(_11407_),
    .Q(\top_ihp.oisc.regs[58][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1386),
    .D(_02074_),
    .Q_N(_11406_),
    .Q(\top_ihp.oisc.regs[58][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1367),
    .D(_02075_),
    .Q_N(_11405_),
    .Q(\top_ihp.oisc.regs[58][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1372),
    .D(_02076_),
    .Q_N(_11404_),
    .Q(\top_ihp.oisc.regs[58][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1340),
    .D(_02077_),
    .Q_N(_11403_),
    .Q(\top_ihp.oisc.regs[58][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1331),
    .D(_02078_),
    .Q_N(_11402_),
    .Q(\top_ihp.oisc.regs[58][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1330),
    .D(_02079_),
    .Q_N(_11401_),
    .Q(\top_ihp.oisc.regs[58][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1327),
    .D(_02080_),
    .Q_N(_11400_),
    .Q(\top_ihp.oisc.regs[58][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1316),
    .D(_02081_),
    .Q_N(_11399_),
    .Q(\top_ihp.oisc.regs[58][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1312),
    .D(_02082_),
    .Q_N(_11398_),
    .Q(\top_ihp.oisc.regs[58][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1312),
    .D(_02083_),
    .Q_N(_11397_),
    .Q(\top_ihp.oisc.regs[58][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1306),
    .D(_02084_),
    .Q_N(_11396_),
    .Q(\top_ihp.oisc.regs[58][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1280),
    .D(_02085_),
    .Q_N(_11395_),
    .Q(\top_ihp.oisc.regs[58][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1349),
    .D(_02086_),
    .Q_N(_11394_),
    .Q(\top_ihp.oisc.regs[59][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1284),
    .D(_02087_),
    .Q_N(_11393_),
    .Q(\top_ihp.oisc.regs[59][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1206),
    .D(_02088_),
    .Q_N(_11392_),
    .Q(\top_ihp.oisc.regs[59][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1279),
    .D(_02089_),
    .Q_N(_11391_),
    .Q(\top_ihp.oisc.regs[59][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1219),
    .D(_02090_),
    .Q_N(_11390_),
    .Q(\top_ihp.oisc.regs[59][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1278),
    .D(_02091_),
    .Q_N(_11389_),
    .Q(\top_ihp.oisc.regs[59][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1207),
    .D(_02092_),
    .Q_N(_11388_),
    .Q(\top_ihp.oisc.regs[59][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1252),
    .D(_02093_),
    .Q_N(_11387_),
    .Q(\top_ihp.oisc.regs[59][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1215),
    .D(_02094_),
    .Q_N(_11386_),
    .Q(\top_ihp.oisc.regs[59][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1220),
    .D(_02095_),
    .Q_N(_11385_),
    .Q(\top_ihp.oisc.regs[59][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1217),
    .D(_02096_),
    .Q_N(_11384_),
    .Q(\top_ihp.oisc.regs[59][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1334),
    .D(_02097_),
    .Q_N(_11383_),
    .Q(\top_ihp.oisc.regs[59][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1350),
    .D(_02098_),
    .Q_N(_11382_),
    .Q(\top_ihp.oisc.regs[59][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1359),
    .D(_02099_),
    .Q_N(_11381_),
    .Q(\top_ihp.oisc.regs[59][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1357),
    .D(_02100_),
    .Q_N(_11380_),
    .Q(\top_ihp.oisc.regs[59][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1265),
    .D(_02101_),
    .Q_N(_11379_),
    .Q(\top_ihp.oisc.regs[59][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1254),
    .D(_02102_),
    .Q_N(_11378_),
    .Q(\top_ihp.oisc.regs[59][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1354),
    .D(_02103_),
    .Q_N(_11377_),
    .Q(\top_ihp.oisc.regs[59][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1359),
    .D(_02104_),
    .Q_N(_11376_),
    .Q(\top_ihp.oisc.regs[59][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1357),
    .D(_02105_),
    .Q_N(_11375_),
    .Q(\top_ihp.oisc.regs[59][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1367),
    .D(_02106_),
    .Q_N(_11374_),
    .Q(\top_ihp.oisc.regs[59][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1367),
    .D(_02107_),
    .Q_N(_11373_),
    .Q(\top_ihp.oisc.regs[59][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1340),
    .D(_02108_),
    .Q_N(_11372_),
    .Q(\top_ihp.oisc.regs[59][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1371),
    .D(_02109_),
    .Q_N(_11371_),
    .Q(\top_ihp.oisc.regs[59][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1330),
    .D(_02110_),
    .Q_N(_11370_),
    .Q(\top_ihp.oisc.regs[59][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1297),
    .D(_02111_),
    .Q_N(_11369_),
    .Q(\top_ihp.oisc.regs[59][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1327),
    .D(_02112_),
    .Q_N(_11368_),
    .Q(\top_ihp.oisc.regs[59][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1328),
    .D(_02113_),
    .Q_N(_11367_),
    .Q(\top_ihp.oisc.regs[59][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1285),
    .D(_02114_),
    .Q_N(_11366_),
    .Q(\top_ihp.oisc.regs[59][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1315),
    .D(_02115_),
    .Q_N(_11365_),
    .Q(\top_ihp.oisc.regs[59][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1285),
    .D(_02116_),
    .Q_N(_11364_),
    .Q(\top_ihp.oisc.regs[59][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1286),
    .D(_02117_),
    .Q_N(_11363_),
    .Q(\top_ihp.oisc.regs[59][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1164),
    .D(_02118_),
    .Q_N(_11362_),
    .Q(\top_ihp.oisc.regs[5][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1175),
    .D(_02119_),
    .Q_N(_11361_),
    .Q(\top_ihp.oisc.regs[5][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1176),
    .D(_02120_),
    .Q_N(_11360_),
    .Q(\top_ihp.oisc.regs[5][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1186),
    .D(_02121_),
    .Q_N(_11359_),
    .Q(\top_ihp.oisc.regs[5][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1236),
    .D(_02122_),
    .Q_N(_11358_),
    .Q(\top_ihp.oisc.regs[5][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1189),
    .D(_02123_),
    .Q_N(_11357_),
    .Q(\top_ihp.oisc.regs[5][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1195),
    .D(_02124_),
    .Q_N(_11356_),
    .Q(\top_ihp.oisc.regs[5][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1236),
    .D(_02125_),
    .Q_N(_11355_),
    .Q(\top_ihp.oisc.regs[5][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1186),
    .D(_02126_),
    .Q_N(_11354_),
    .Q(\top_ihp.oisc.regs[5][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1187),
    .D(_02127_),
    .Q_N(_11353_),
    .Q(\top_ihp.oisc.regs[5][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1213),
    .D(_02128_),
    .Q_N(_11352_),
    .Q(\top_ihp.oisc.regs[5][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1246),
    .D(_02129_),
    .Q_N(_11351_),
    .Q(\top_ihp.oisc.regs[5][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1226),
    .D(_02130_),
    .Q_N(_11350_),
    .Q(\top_ihp.oisc.regs[5][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1231),
    .D(_02131_),
    .Q_N(_11349_),
    .Q(\top_ihp.oisc.regs[5][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1235),
    .D(_02132_),
    .Q_N(_11348_),
    .Q(\top_ihp.oisc.regs[5][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1164),
    .D(_02133_),
    .Q_N(_11347_),
    .Q(\top_ihp.oisc.regs[5][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1237),
    .D(_02134_),
    .Q_N(_11346_),
    .Q(\top_ihp.oisc.regs[5][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1238),
    .D(_02135_),
    .Q_N(_11345_),
    .Q(\top_ihp.oisc.regs[5][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1231),
    .D(_02136_),
    .Q_N(_11344_),
    .Q(\top_ihp.oisc.regs[5][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1237),
    .D(_02137_),
    .Q_N(_11343_),
    .Q(\top_ihp.oisc.regs[5][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1238),
    .D(_02138_),
    .Q_N(_11342_),
    .Q(\top_ihp.oisc.regs[5][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1231),
    .D(_02139_),
    .Q_N(_11341_),
    .Q(\top_ihp.oisc.regs[5][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1230),
    .D(_02140_),
    .Q_N(_11340_),
    .Q(\top_ihp.oisc.regs[5][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1228),
    .D(_02141_),
    .Q_N(_11339_),
    .Q(\top_ihp.oisc.regs[5][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1188),
    .D(_02142_),
    .Q_N(_11338_),
    .Q(\top_ihp.oisc.regs[5][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1187),
    .D(_02143_),
    .Q_N(_11337_),
    .Q(\top_ihp.oisc.regs[5][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1189),
    .D(_02144_),
    .Q_N(_11336_),
    .Q(\top_ihp.oisc.regs[5][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1185),
    .D(_02145_),
    .Q_N(_11335_),
    .Q(\top_ihp.oisc.regs[5][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1174),
    .D(_02146_),
    .Q_N(_11334_),
    .Q(\top_ihp.oisc.regs[5][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1174),
    .D(_02147_),
    .Q_N(_11333_),
    .Q(\top_ihp.oisc.regs[5][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1178),
    .D(_02148_),
    .Q_N(_11332_),
    .Q(\top_ihp.oisc.regs[5][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1174),
    .D(_02149_),
    .Q_N(_11331_),
    .Q(\top_ihp.oisc.regs[5][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1346),
    .D(_02150_),
    .Q_N(_11330_),
    .Q(\top_ihp.oisc.regs[60][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1284),
    .D(_02151_),
    .Q_N(_11329_),
    .Q(\top_ihp.oisc.regs[60][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1206),
    .D(_02152_),
    .Q_N(_11328_),
    .Q(\top_ihp.oisc.regs[60][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1293),
    .D(_02153_),
    .Q_N(_11327_),
    .Q(\top_ihp.oisc.regs[60][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1248),
    .D(_02154_),
    .Q_N(_11326_),
    .Q(\top_ihp.oisc.regs[60][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1204),
    .D(_02155_),
    .Q_N(_11325_),
    .Q(\top_ihp.oisc.regs[60][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1206),
    .D(_02156_),
    .Q_N(_11324_),
    .Q(\top_ihp.oisc.regs[60][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1252),
    .D(_02157_),
    .Q_N(_11323_),
    .Q(\top_ihp.oisc.regs[60][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1196),
    .D(_02158_),
    .Q_N(_11322_),
    .Q(\top_ihp.oisc.regs[60][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1219),
    .D(_02159_),
    .Q_N(_11321_),
    .Q(\top_ihp.oisc.regs[60][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1211),
    .D(_02160_),
    .Q_N(_11320_),
    .Q(\top_ihp.oisc.regs[60][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1339),
    .D(_02161_),
    .Q_N(_11319_),
    .Q(\top_ihp.oisc.regs[60][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1270),
    .D(_02162_),
    .Q_N(_11318_),
    .Q(\top_ihp.oisc.regs[60][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1359),
    .D(_02163_),
    .Q_N(_11317_),
    .Q(\top_ihp.oisc.regs[60][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1357),
    .D(_02164_),
    .Q_N(_11316_),
    .Q(\top_ihp.oisc.regs[60][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1264),
    .D(_02165_),
    .Q_N(_11315_),
    .Q(\top_ihp.oisc.regs[60][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1389),
    .D(_02166_),
    .Q_N(_11314_),
    .Q(\top_ihp.oisc.regs[60][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1381),
    .D(_02167_),
    .Q_N(_11313_),
    .Q(\top_ihp.oisc.regs[60][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1342),
    .D(_02168_),
    .Q_N(_11312_),
    .Q(\top_ihp.oisc.regs[60][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1389),
    .D(_02169_),
    .Q_N(_11311_),
    .Q(\top_ihp.oisc.regs[60][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1388),
    .D(_02170_),
    .Q_N(_11310_),
    .Q(\top_ihp.oisc.regs[60][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1373),
    .D(_02171_),
    .Q_N(_11309_),
    .Q(\top_ihp.oisc.regs[60][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1366),
    .D(_02172_),
    .Q_N(_11308_),
    .Q(\top_ihp.oisc.regs[60][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1340),
    .D(_02173_),
    .Q_N(_11307_),
    .Q(\top_ihp.oisc.regs[60][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1298),
    .D(_02174_),
    .Q_N(_11306_),
    .Q(\top_ihp.oisc.regs[60][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1323),
    .D(_02175_),
    .Q_N(_11305_),
    .Q(\top_ihp.oisc.regs[60][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1319),
    .D(_02176_),
    .Q_N(_11304_),
    .Q(\top_ihp.oisc.regs[60][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1321),
    .D(_02177_),
    .Q_N(_11303_),
    .Q(\top_ihp.oisc.regs[60][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1302),
    .D(_02178_),
    .Q_N(_11302_),
    .Q(\top_ihp.oisc.regs[60][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1304),
    .D(_02179_),
    .Q_N(_11301_),
    .Q(\top_ihp.oisc.regs[60][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1306),
    .D(_02180_),
    .Q_N(_11300_),
    .Q(\top_ihp.oisc.regs[60][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1295),
    .D(_02181_),
    .Q_N(_11299_),
    .Q(\top_ihp.oisc.regs[60][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1346),
    .D(_02182_),
    .Q_N(_11298_),
    .Q(\top_ihp.oisc.regs[61][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1286),
    .D(_02183_),
    .Q_N(_11297_),
    .Q(\top_ihp.oisc.regs[61][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1205),
    .D(_02184_),
    .Q_N(_11296_),
    .Q(\top_ihp.oisc.regs[61][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1278),
    .D(_02185_),
    .Q_N(_11295_),
    .Q(\top_ihp.oisc.regs[61][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1252),
    .D(_02186_),
    .Q_N(_11294_),
    .Q(\top_ihp.oisc.regs[61][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1288),
    .D(_02187_),
    .Q_N(_11293_),
    .Q(\top_ihp.oisc.regs[61][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1197),
    .D(_02188_),
    .Q_N(_11292_),
    .Q(\top_ihp.oisc.regs[61][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1252),
    .D(_02189_),
    .Q_N(_11291_),
    .Q(\top_ihp.oisc.regs[61][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1207),
    .D(_02190_),
    .Q_N(_11290_),
    .Q(\top_ihp.oisc.regs[61][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1291),
    .D(_02191_),
    .Q_N(_11289_),
    .Q(\top_ihp.oisc.regs[61][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1212),
    .D(_02192_),
    .Q_N(_11288_),
    .Q(\top_ihp.oisc.regs[61][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1251),
    .D(_02193_),
    .Q_N(_11287_),
    .Q(\top_ihp.oisc.regs[61][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1349),
    .D(_02194_),
    .Q_N(_11286_),
    .Q(\top_ihp.oisc.regs[61][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1253),
    .D(_02195_),
    .Q_N(_11285_),
    .Q(\top_ihp.oisc.regs[61][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1347),
    .D(_02196_),
    .Q_N(_11284_),
    .Q(\top_ihp.oisc.regs[61][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1264),
    .D(_02197_),
    .Q_N(_11283_),
    .Q(\top_ihp.oisc.regs[61][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1345),
    .D(_02198_),
    .Q_N(_11282_),
    .Q(\top_ihp.oisc.regs[61][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1336),
    .D(_02199_),
    .Q_N(_11281_),
    .Q(\top_ihp.oisc.regs[61][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1378),
    .D(_02200_),
    .Q_N(_11280_),
    .Q(\top_ihp.oisc.regs[61][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1379),
    .D(_02201_),
    .Q_N(_11279_),
    .Q(\top_ihp.oisc.regs[61][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1375),
    .D(_02202_),
    .Q_N(_11278_),
    .Q(\top_ihp.oisc.regs[61][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1374),
    .D(_02203_),
    .Q_N(_11277_),
    .Q(\top_ihp.oisc.regs[61][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1366),
    .D(_02204_),
    .Q_N(_11276_),
    .Q(\top_ihp.oisc.regs[61][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1371),
    .D(_02205_),
    .Q_N(_11275_),
    .Q(\top_ihp.oisc.regs[61][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1323),
    .D(_02206_),
    .Q_N(_11274_),
    .Q(\top_ihp.oisc.regs[61][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1331),
    .D(_02207_),
    .Q_N(_11273_),
    .Q(\top_ihp.oisc.regs[61][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1327),
    .D(_02208_),
    .Q_N(_11272_),
    .Q(\top_ihp.oisc.regs[61][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1316),
    .D(_02209_),
    .Q_N(_11271_),
    .Q(\top_ihp.oisc.regs[61][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1316),
    .D(_02210_),
    .Q_N(_11270_),
    .Q(\top_ihp.oisc.regs[61][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1316),
    .D(_02211_),
    .Q_N(_11269_),
    .Q(\top_ihp.oisc.regs[61][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1319),
    .D(_02212_),
    .Q_N(_11268_),
    .Q(\top_ihp.oisc.regs[61][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1293),
    .D(_02213_),
    .Q_N(_11267_),
    .Q(\top_ihp.oisc.regs[61][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1349),
    .D(_02214_),
    .Q_N(_11266_),
    .Q(\top_ihp.oisc.regs[62][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1286),
    .D(_02215_),
    .Q_N(_11265_),
    .Q(\top_ihp.oisc.regs[62][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1273),
    .D(_02216_),
    .Q_N(_11264_),
    .Q(\top_ihp.oisc.regs[62][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1279),
    .D(_02217_),
    .Q_N(_11263_),
    .Q(\top_ihp.oisc.regs[62][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1254),
    .D(_02218_),
    .Q_N(_11262_),
    .Q(\top_ihp.oisc.regs[62][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1289),
    .D(_02219_),
    .Q_N(_11261_),
    .Q(\top_ihp.oisc.regs[62][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1216),
    .D(_02220_),
    .Q_N(_11260_),
    .Q(\top_ihp.oisc.regs[62][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1254),
    .D(_02221_),
    .Q_N(_11259_),
    .Q(\top_ihp.oisc.regs[62][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1216),
    .D(_02222_),
    .Q_N(_11258_),
    .Q(\top_ihp.oisc.regs[62][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1255),
    .D(_02223_),
    .Q_N(_11257_),
    .Q(\top_ihp.oisc.regs[62][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1217),
    .D(_02224_),
    .Q_N(_11256_),
    .Q(\top_ihp.oisc.regs[62][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1296),
    .D(_02225_),
    .Q_N(_11255_),
    .Q(\top_ihp.oisc.regs[62][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1270),
    .D(_02226_),
    .Q_N(_11254_),
    .Q(\top_ihp.oisc.regs[62][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1342),
    .D(_02227_),
    .Q_N(_11253_),
    .Q(\top_ihp.oisc.regs[62][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1348),
    .D(_02228_),
    .Q_N(_11252_),
    .Q(\top_ihp.oisc.regs[62][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1265),
    .D(_02229_),
    .Q_N(_11251_),
    .Q(\top_ihp.oisc.regs[62][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1355),
    .D(_02230_),
    .Q_N(_11250_),
    .Q(\top_ihp.oisc.regs[62][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1380),
    .D(_02231_),
    .Q_N(_11249_),
    .Q(\top_ihp.oisc.regs[62][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1381),
    .D(_02232_),
    .Q_N(_11248_),
    .Q(\top_ihp.oisc.regs[62][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1379),
    .D(_02233_),
    .Q_N(_11247_),
    .Q(\top_ihp.oisc.regs[62][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1375),
    .D(_02234_),
    .Q_N(_11246_),
    .Q(\top_ihp.oisc.regs[62][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1374),
    .D(_02235_),
    .Q_N(_11245_),
    .Q(\top_ihp.oisc.regs[62][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1372),
    .D(_02236_),
    .Q_N(_11244_),
    .Q(\top_ihp.oisc.regs[62][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1372),
    .D(_02237_),
    .Q_N(_11243_),
    .Q(\top_ihp.oisc.regs[62][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1331),
    .D(_02238_),
    .Q_N(_11242_),
    .Q(\top_ihp.oisc.regs[62][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1332),
    .D(_02239_),
    .Q_N(_11241_),
    .Q(\top_ihp.oisc.regs[62][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1328),
    .D(_02240_),
    .Q_N(_11240_),
    .Q(\top_ihp.oisc.regs[62][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1316),
    .D(_02241_),
    .Q_N(_11239_),
    .Q(\top_ihp.oisc.regs[62][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1312),
    .D(_02242_),
    .Q_N(_11238_),
    .Q(\top_ihp.oisc.regs[62][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1315),
    .D(_02243_),
    .Q_N(_11237_),
    .Q(\top_ihp.oisc.regs[62][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1306),
    .D(_02244_),
    .Q_N(_11236_),
    .Q(\top_ihp.oisc.regs[62][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1282),
    .D(_02245_),
    .Q_N(_11235_),
    .Q(\top_ihp.oisc.regs[62][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1258),
    .D(_02246_),
    .Q_N(_11234_),
    .Q(\top_ihp.oisc.regs[63][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1194),
    .D(_02247_),
    .Q_N(_11233_),
    .Q(\top_ihp.oisc.regs[63][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1195),
    .D(_02248_),
    .Q_N(_11232_),
    .Q(\top_ihp.oisc.regs[63][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1209),
    .D(_02249_),
    .Q_N(_11231_),
    .Q(\top_ihp.oisc.regs[63][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1213),
    .D(_02250_),
    .Q_N(_11230_),
    .Q(\top_ihp.oisc.regs[63][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1194),
    .D(_02251_),
    .Q_N(_11229_),
    .Q(\top_ihp.oisc.regs[63][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1198),
    .D(_02252_),
    .Q_N(_11228_),
    .Q(\top_ihp.oisc.regs[63][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1213),
    .D(_02253_),
    .Q_N(_11227_),
    .Q(\top_ihp.oisc.regs[63][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1195),
    .D(_02254_),
    .Q_N(_11226_),
    .Q(\top_ihp.oisc.regs[63][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1213),
    .D(_02255_),
    .Q_N(_11225_),
    .Q(\top_ihp.oisc.regs[63][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1210),
    .D(_02256_),
    .Q_N(_11224_),
    .Q(\top_ihp.oisc.regs[63][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1246),
    .D(_02257_),
    .Q_N(_11223_),
    .Q(\top_ihp.oisc.regs[63][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1257),
    .D(_02258_),
    .Q_N(_11222_),
    .Q(\top_ihp.oisc.regs[63][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1248),
    .D(_02259_),
    .Q_N(_11221_),
    .Q(\top_ihp.oisc.regs[63][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1357),
    .D(_02260_),
    .Q_N(_11220_),
    .Q(\top_ihp.oisc.regs[63][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1257),
    .D(_02261_),
    .Q_N(_11219_),
    .Q(\top_ihp.oisc.regs[63][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1387),
    .D(_02262_),
    .Q_N(_11218_),
    .Q(\top_ihp.oisc.regs[63][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1248),
    .D(_02263_),
    .Q_N(_11217_),
    .Q(\top_ihp.oisc.regs[63][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1248),
    .D(_02264_),
    .Q_N(_11216_),
    .Q(\top_ihp.oisc.regs[63][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1388),
    .D(_02265_),
    .Q_N(_11215_),
    .Q(\top_ihp.oisc.regs[63][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1391),
    .D(_02266_),
    .Q_N(_11214_),
    .Q(\top_ihp.oisc.regs[63][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1253),
    .D(_02267_),
    .Q_N(_11213_),
    .Q(\top_ihp.oisc.regs[63][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1365),
    .D(_02268_),
    .Q_N(_11212_),
    .Q(\top_ihp.oisc.regs[63][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1246),
    .D(_02269_),
    .Q_N(_11211_),
    .Q(\top_ihp.oisc.regs[63][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1330),
    .D(_02270_),
    .Q_N(_11210_),
    .Q(\top_ihp.oisc.regs[63][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1330),
    .D(_02271_),
    .Q_N(_11209_),
    .Q(\top_ihp.oisc.regs[63][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1328),
    .D(_02272_),
    .Q_N(_11208_),
    .Q(\top_ihp.oisc.regs[63][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1308),
    .D(_02273_),
    .Q_N(_11207_),
    .Q(\top_ihp.oisc.regs[63][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1195),
    .D(_02274_),
    .Q_N(_11206_),
    .Q(\top_ihp.oisc.regs[63][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1307),
    .D(_02275_),
    .Q_N(_11205_),
    .Q(\top_ihp.oisc.regs[63][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1191),
    .D(_02276_),
    .Q_N(_11204_),
    .Q(\top_ihp.oisc.regs[63][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1194),
    .D(_02277_),
    .Q_N(_11203_),
    .Q(\top_ihp.oisc.regs[63][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1165),
    .D(_02278_),
    .Q_N(_11202_),
    .Q(\top_ihp.oisc.regs[6][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1171),
    .D(_02279_),
    .Q_N(_11201_),
    .Q(\top_ihp.oisc.regs[6][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1171),
    .D(_02280_),
    .Q_N(_11200_),
    .Q(\top_ihp.oisc.regs[6][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1181),
    .D(_02281_),
    .Q_N(_11199_),
    .Q(\top_ihp.oisc.regs[6][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1223),
    .D(_02282_),
    .Q_N(_11198_),
    .Q(\top_ihp.oisc.regs[6][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1180),
    .D(_02283_),
    .Q_N(_11197_),
    .Q(\top_ihp.oisc.regs[6][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1172),
    .D(_02284_),
    .Q_N(_11196_),
    .Q(\top_ihp.oisc.regs[6][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1224),
    .D(_02285_),
    .Q_N(_11195_),
    .Q(\top_ihp.oisc.regs[6][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1180),
    .D(_02286_),
    .Q_N(_11194_),
    .Q(\top_ihp.oisc.regs[6][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1182),
    .D(_02287_),
    .Q_N(_11193_),
    .Q(\top_ihp.oisc.regs[6][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1183),
    .D(_02288_),
    .Q_N(_11192_),
    .Q(\top_ihp.oisc.regs[6][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1153),
    .D(_02289_),
    .Q_N(_11191_),
    .Q(\top_ihp.oisc.regs[6][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1241),
    .D(_02290_),
    .Q_N(_11190_),
    .Q(\top_ihp.oisc.regs[6][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1226),
    .D(_02291_),
    .Q_N(_11189_),
    .Q(\top_ihp.oisc.regs[6][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1163),
    .D(_02292_),
    .Q_N(_11188_),
    .Q(\top_ihp.oisc.regs[6][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1165),
    .D(_02293_),
    .Q_N(_11187_),
    .Q(\top_ihp.oisc.regs[6][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1155),
    .D(_02294_),
    .Q_N(_11186_),
    .Q(\top_ihp.oisc.regs[6][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1162),
    .D(_02295_),
    .Q_N(_11185_),
    .Q(\top_ihp.oisc.regs[6][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1156),
    .D(_02296_),
    .Q_N(_11184_),
    .Q(\top_ihp.oisc.regs[6][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1234),
    .D(_02297_),
    .Q_N(_11183_),
    .Q(\top_ihp.oisc.regs[6][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1234),
    .D(_02298_),
    .Q_N(_11182_),
    .Q(\top_ihp.oisc.regs[6][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1226),
    .D(_02299_),
    .Q_N(_11181_),
    .Q(\top_ihp.oisc.regs[6][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1224),
    .D(_02300_),
    .Q_N(_11180_),
    .Q(\top_ihp.oisc.regs[6][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1223),
    .D(_02301_),
    .Q_N(_11179_),
    .Q(\top_ihp.oisc.regs[6][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1182),
    .D(_02302_),
    .Q_N(_11178_),
    .Q(\top_ihp.oisc.regs[6][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1183),
    .D(_02303_),
    .Q_N(_11177_),
    .Q(\top_ihp.oisc.regs[6][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1181),
    .D(_02304_),
    .Q_N(_11176_),
    .Q(\top_ihp.oisc.regs[6][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1181),
    .D(_02305_),
    .Q_N(_11175_),
    .Q(\top_ihp.oisc.regs[6][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1170),
    .D(_02306_),
    .Q_N(_11174_),
    .Q(\top_ihp.oisc.regs[6][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1170),
    .D(_02307_),
    .Q_N(_11173_),
    .Q(\top_ihp.oisc.regs[6][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1170),
    .D(_02308_),
    .Q_N(_11172_),
    .Q(\top_ihp.oisc.regs[6][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1173),
    .D(_02309_),
    .Q_N(_11171_),
    .Q(\top_ihp.oisc.regs[6][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1236),
    .D(_02310_),
    .Q_N(_11170_),
    .Q(\top_ihp.oisc.regs[7][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1120),
    .D(_02311_),
    .Q_N(_11169_),
    .Q(\top_ihp.oisc.regs[7][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1120),
    .D(_02312_),
    .Q_N(_11168_),
    .Q(\top_ihp.oisc.regs[7][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1120),
    .D(_02313_),
    .Q_N(_11167_),
    .Q(\top_ihp.oisc.regs[7][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1235),
    .D(_02314_),
    .Q_N(_11166_),
    .Q(\top_ihp.oisc.regs[7][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1124),
    .D(_02315_),
    .Q_N(_11165_),
    .Q(\top_ihp.oisc.regs[7][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1170),
    .D(_02316_),
    .Q_N(_11164_),
    .Q(\top_ihp.oisc.regs[7][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1236),
    .D(_02317_),
    .Q_N(_11163_),
    .Q(\top_ihp.oisc.regs[7][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1127),
    .D(_02318_),
    .Q_N(_11162_),
    .Q(\top_ihp.oisc.regs[7][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1180),
    .D(_02319_),
    .Q_N(_11161_),
    .Q(\top_ihp.oisc.regs[7][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1131),
    .D(_02320_),
    .Q_N(_11160_),
    .Q(\top_ihp.oisc.regs[7][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1131),
    .D(_02321_),
    .Q_N(_11159_),
    .Q(\top_ihp.oisc.regs[7][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1150),
    .D(_02322_),
    .Q_N(_11158_),
    .Q(\top_ihp.oisc.regs[7][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1156),
    .D(_02323_),
    .Q_N(_11157_),
    .Q(\top_ihp.oisc.regs[7][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1165),
    .D(_02324_),
    .Q_N(_11156_),
    .Q(\top_ihp.oisc.regs[7][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1160),
    .D(_02325_),
    .Q_N(_11155_),
    .Q(\top_ihp.oisc.regs[7][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1151),
    .D(_02326_),
    .Q_N(_11154_),
    .Q(\top_ihp.oisc.regs[7][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1151),
    .D(_02327_),
    .Q_N(_11153_),
    .Q(\top_ihp.oisc.regs[7][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1156),
    .D(_02328_),
    .Q_N(_11152_),
    .Q(\top_ihp.oisc.regs[7][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1233),
    .D(_02329_),
    .Q_N(_11151_),
    .Q(\top_ihp.oisc.regs[7][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1233),
    .D(_02330_),
    .Q_N(_11150_),
    .Q(\top_ihp.oisc.regs[7][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1226),
    .D(_02331_),
    .Q_N(_11149_),
    .Q(\top_ihp.oisc.regs[7][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1152),
    .D(_02332_),
    .Q_N(_11148_),
    .Q(\top_ihp.oisc.regs[7][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1154),
    .D(_02333_),
    .Q_N(_11147_),
    .Q(\top_ihp.oisc.regs[7][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1223),
    .D(_02334_),
    .Q_N(_11146_),
    .Q(\top_ihp.oisc.regs[7][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1115),
    .D(_02335_),
    .Q_N(_11145_),
    .Q(\top_ihp.oisc.regs[7][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1117),
    .D(_02336_),
    .Q_N(_11144_),
    .Q(\top_ihp.oisc.regs[7][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1132),
    .D(_02337_),
    .Q_N(_11143_),
    .Q(\top_ihp.oisc.regs[7][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1111),
    .D(_02338_),
    .Q_N(_11142_),
    .Q(\top_ihp.oisc.regs[7][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1111),
    .D(_02339_),
    .Q_N(_11141_),
    .Q(\top_ihp.oisc.regs[7][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1111),
    .D(_02340_),
    .Q_N(_11140_),
    .Q(\top_ihp.oisc.regs[7][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1120),
    .D(_02341_),
    .Q_N(_11139_),
    .Q(\top_ihp.oisc.regs[7][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1159),
    .D(_02342_),
    .Q_N(_11138_),
    .Q(\top_ihp.oisc.regs[8][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1127),
    .D(_02343_),
    .Q_N(_11137_),
    .Q(\top_ihp.oisc.regs[8][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1126),
    .D(_02344_),
    .Q_N(_11136_),
    .Q(\top_ihp.oisc.regs[8][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1171),
    .D(_02345_),
    .Q_N(_11135_),
    .Q(\top_ihp.oisc.regs[8][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1154),
    .D(_02346_),
    .Q_N(_11134_),
    .Q(\top_ihp.oisc.regs[8][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1134),
    .D(_02347_),
    .Q_N(_11133_),
    .Q(\top_ihp.oisc.regs[8][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1171),
    .D(_02348_),
    .Q_N(_11132_),
    .Q(\top_ihp.oisc.regs[8][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1154),
    .D(_02349_),
    .Q_N(_11131_),
    .Q(\top_ihp.oisc.regs[8][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1180),
    .D(_02350_),
    .Q_N(_11130_),
    .Q(\top_ihp.oisc.regs[8][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1182),
    .D(_02351_),
    .Q_N(_11129_),
    .Q(\top_ihp.oisc.regs[8][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1134),
    .D(_02352_),
    .Q_N(_11128_),
    .Q(\top_ihp.oisc.regs[8][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1149),
    .D(_02353_),
    .Q_N(_11127_),
    .Q(\top_ihp.oisc.regs[8][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1159),
    .D(_02354_),
    .Q_N(_11126_),
    .Q(\top_ihp.oisc.regs[8][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1150),
    .D(_02355_),
    .Q_N(_11125_),
    .Q(\top_ihp.oisc.regs[8][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1158),
    .D(_02356_),
    .Q_N(_11124_),
    .Q(\top_ihp.oisc.regs[8][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1159),
    .D(_02357_),
    .Q_N(_11123_),
    .Q(\top_ihp.oisc.regs[8][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1150),
    .D(_02358_),
    .Q_N(_11122_),
    .Q(\top_ihp.oisc.regs[8][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1158),
    .D(_02359_),
    .Q_N(_11121_),
    .Q(\top_ihp.oisc.regs[8][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1150),
    .D(_02360_),
    .Q_N(_11120_),
    .Q(\top_ihp.oisc.regs[8][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1148),
    .D(_02361_),
    .Q_N(_11119_),
    .Q(\top_ihp.oisc.regs[8][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1158),
    .D(_02362_),
    .Q_N(_11118_),
    .Q(\top_ihp.oisc.regs[8][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1140),
    .D(_02363_),
    .Q_N(_11117_),
    .Q(\top_ihp.oisc.regs[8][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1150),
    .D(_02364_),
    .Q_N(_11116_),
    .Q(\top_ihp.oisc.regs[8][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1149),
    .D(_02365_),
    .Q_N(_11115_),
    .Q(\top_ihp.oisc.regs[8][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1136),
    .D(_02366_),
    .Q_N(_11114_),
    .Q(\top_ihp.oisc.regs[8][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1135),
    .D(_02367_),
    .Q_N(_11113_),
    .Q(\top_ihp.oisc.regs[8][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1134),
    .D(_02368_),
    .Q_N(_11112_),
    .Q(\top_ihp.oisc.regs[8][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1129),
    .D(_02369_),
    .Q_N(_11111_),
    .Q(\top_ihp.oisc.regs[8][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1119),
    .D(_02370_),
    .Q_N(_11110_),
    .Q(\top_ihp.oisc.regs[8][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1119),
    .D(_02371_),
    .Q_N(_11109_),
    .Q(\top_ihp.oisc.regs[8][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1110),
    .D(_02372_),
    .Q_N(_11108_),
    .Q(\top_ihp.oisc.regs[8][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1122),
    .D(_02373_),
    .Q_N(_11107_),
    .Q(\top_ihp.oisc.regs[8][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1151),
    .D(_02374_),
    .Q_N(_11106_),
    .Q(\top_ihp.oisc.regs[9][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1125),
    .D(_02375_),
    .Q_N(_11105_),
    .Q(\top_ihp.oisc.regs[9][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1126),
    .D(_02376_),
    .Q_N(_11104_),
    .Q(\top_ihp.oisc.regs[9][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1125),
    .D(_02377_),
    .Q_N(_11103_),
    .Q(\top_ihp.oisc.regs[9][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1166),
    .D(_02378_),
    .Q_N(_11102_),
    .Q(\top_ihp.oisc.regs[9][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1133),
    .D(_02379_),
    .Q_N(_11101_),
    .Q(\top_ihp.oisc.regs[9][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1125),
    .D(_02380_),
    .Q_N(_11100_),
    .Q(\top_ihp.oisc.regs[9][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1235),
    .D(_02381_),
    .Q_N(_11099_),
    .Q(\top_ihp.oisc.regs[9][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1134),
    .D(_02382_),
    .Q_N(_11098_),
    .Q(\top_ihp.oisc.regs[9][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1136),
    .D(_02383_),
    .Q_N(_11097_),
    .Q(\top_ihp.oisc.regs[9][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1116),
    .D(_02384_),
    .Q_N(_11096_),
    .Q(\top_ihp.oisc.regs[9][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1116),
    .D(_02385_),
    .Q_N(_11095_),
    .Q(\top_ihp.oisc.regs[9][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1141),
    .D(_02386_),
    .Q_N(_11094_),
    .Q(\top_ihp.oisc.regs[9][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1141),
    .D(_02387_),
    .Q_N(_11093_),
    .Q(\top_ihp.oisc.regs[9][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1235),
    .D(_02388_),
    .Q_N(_11092_),
    .Q(\top_ihp.oisc.regs[9][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1160),
    .D(_02389_),
    .Q_N(_11091_),
    .Q(\top_ihp.oisc.regs[9][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1141),
    .D(_02390_),
    .Q_N(_11090_),
    .Q(\top_ihp.oisc.regs[9][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1141),
    .D(_02391_),
    .Q_N(_11089_),
    .Q(\top_ihp.oisc.regs[9][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1141),
    .D(_02392_),
    .Q_N(_11088_),
    .Q(\top_ihp.oisc.regs[9][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1146),
    .D(_02393_),
    .Q_N(_11087_),
    .Q(\top_ihp.oisc.regs[9][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1146),
    .D(_02394_),
    .Q_N(_11086_),
    .Q(\top_ihp.oisc.regs[9][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1141),
    .D(_02395_),
    .Q_N(_11085_),
    .Q(\top_ihp.oisc.regs[9][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1142),
    .D(_02396_),
    .Q_N(_11084_),
    .Q(\top_ihp.oisc.regs[9][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1142),
    .D(_02397_),
    .Q_N(_11083_),
    .Q(\top_ihp.oisc.regs[9][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1116),
    .D(_02398_),
    .Q_N(_11082_),
    .Q(\top_ihp.oisc.regs[9][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1116),
    .D(_02399_),
    .Q_N(_11081_),
    .Q(\top_ihp.oisc.regs[9][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1114),
    .D(_02400_),
    .Q_N(_11080_),
    .Q(\top_ihp.oisc.regs[9][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1117),
    .D(_02401_),
    .Q_N(_11079_),
    .Q(\top_ihp.oisc.regs[9][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1110),
    .D(_02402_),
    .Q_N(_11078_),
    .Q(\top_ihp.oisc.regs[9][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1110),
    .D(_02403_),
    .Q_N(_11077_),
    .Q(\top_ihp.oisc.regs[9][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1110),
    .D(_02404_),
    .Q_N(_11076_),
    .Q(\top_ihp.oisc.regs[9][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1110),
    .D(_02405_),
    .Q_N(_11075_),
    .Q(\top_ihp.oisc.regs[9][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1105),
    .D(_02406_),
    .Q_N(\top_ihp.oisc.state[0] ),
    .Q(_13205_));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1103),
    .D(_02407_),
    .Q_N(_11074_),
    .Q(\top_ihp.oisc.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1103),
    .D(_02408_),
    .Q_N(_00075_),
    .Q(\top_ihp.oisc.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1103),
    .D(_02409_),
    .Q_N(_00074_),
    .Q(\top_ihp.oisc.state[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1103),
    .D(_02410_),
    .Q_N(_00076_),
    .Q(\top_ihp.oisc.state[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1104),
    .D(_00002_),
    .Q_N(_00069_),
    .Q(\top_ihp.oisc.state[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1103),
    .D(_02411_),
    .Q_N(_11073_),
    .Q(\top_ihp.oisc.state[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1080),
    .D(_02412_),
    .Q_N(_00091_),
    .Q(\top_ihp.oisc.wb_dat_o[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1071),
    .D(_02413_),
    .Q_N(_11072_),
    .Q(\top_ihp.oisc.wb_dat_o[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1071),
    .D(_02414_),
    .Q_N(_11071_),
    .Q(\top_ihp.oisc.wb_dat_o[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1071),
    .D(_02415_),
    .Q_N(_11070_),
    .Q(\top_ihp.oisc.wb_dat_o[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1071),
    .D(_02416_),
    .Q_N(_11069_),
    .Q(\top_ihp.oisc.wb_dat_o[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1070),
    .D(_02417_),
    .Q_N(_11068_),
    .Q(\top_ihp.oisc.wb_dat_o[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1071),
    .D(_02418_),
    .Q_N(_11067_),
    .Q(\top_ihp.oisc.wb_dat_o[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1073),
    .D(_02419_),
    .Q_N(_11066_),
    .Q(\top_ihp.oisc.wb_dat_o[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1074),
    .D(_02420_),
    .Q_N(_11065_),
    .Q(\top_ihp.oisc.wb_dat_o[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1081),
    .D(_02421_),
    .Q_N(_11064_),
    .Q(\top_ihp.oisc.wb_dat_o[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1081),
    .D(_02422_),
    .Q_N(_11063_),
    .Q(\top_ihp.oisc.wb_dat_o[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1072),
    .D(_02423_),
    .Q_N(_00092_),
    .Q(\top_ihp.oisc.wb_dat_o[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1080),
    .D(_02424_),
    .Q_N(_11062_),
    .Q(\top_ihp.oisc.wb_dat_o[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1080),
    .D(_02425_),
    .Q_N(_11061_),
    .Q(\top_ihp.oisc.wb_dat_o[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1080),
    .D(_02426_),
    .Q_N(_11060_),
    .Q(\top_ihp.oisc.wb_dat_o[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1080),
    .D(_02427_),
    .Q_N(_11059_),
    .Q(\top_ihp.oisc.wb_dat_o[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1074),
    .D(_02428_),
    .Q_N(_11058_),
    .Q(\top_ihp.oisc.wb_dat_o[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1073),
    .D(_02429_),
    .Q_N(_11057_),
    .Q(\top_ihp.oisc.wb_dat_o[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1073),
    .D(_02430_),
    .Q_N(_11056_),
    .Q(\top_ihp.oisc.wb_dat_o[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1072),
    .D(_02431_),
    .Q_N(_11055_),
    .Q(\top_ihp.oisc.wb_dat_o[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1073),
    .D(_02432_),
    .Q_N(_11054_),
    .Q(\top_ihp.oisc.wb_dat_o[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1073),
    .D(_02433_),
    .Q_N(_11053_),
    .Q(\top_ihp.oisc.wb_dat_o[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1072),
    .D(_02434_),
    .Q_N(_00093_),
    .Q(\top_ihp.oisc.wb_dat_o[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1073),
    .D(_02435_),
    .Q_N(_11052_),
    .Q(\top_ihp.oisc.wb_dat_o[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1073),
    .D(_02436_),
    .Q_N(_11051_),
    .Q(\top_ihp.oisc.wb_dat_o[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1072),
    .D(_02437_),
    .Q_N(_00094_),
    .Q(\top_ihp.oisc.wb_dat_o[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1072),
    .D(_02438_),
    .Q_N(_00095_),
    .Q(\top_ihp.oisc.wb_dat_o[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1074),
    .D(_02439_),
    .Q_N(_00096_),
    .Q(\top_ihp.oisc.wb_dat_o[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1070),
    .D(_02440_),
    .Q_N(_00097_),
    .Q(\top_ihp.oisc.wb_dat_o[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1072),
    .D(_02441_),
    .Q_N(_00098_),
    .Q(\top_ihp.oisc.wb_dat_o[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1070),
    .D(_02442_),
    .Q_N(_11050_),
    .Q(\top_ihp.oisc.wb_dat_o[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1071),
    .D(_02443_),
    .Q_N(_11049_),
    .Q(\top_ihp.oisc.wb_dat_o[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1957),
    .D(_02444_),
    .Q_N(_00138_),
    .Q(\top_ihp.wb_emem.bit_counter[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1958),
    .D(_02445_),
    .Q_N(_11048_),
    .Q(\top_ihp.wb_emem.bit_counter[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1959),
    .D(_02446_),
    .Q_N(_11047_),
    .Q(\top_ihp.wb_emem.bit_counter[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1960),
    .D(_02447_),
    .Q_N(_11046_),
    .Q(\top_ihp.wb_emem.bit_counter[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1961),
    .D(_02448_),
    .Q_N(_11045_),
    .Q(\top_ihp.wb_emem.bit_counter[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1962),
    .D(_02449_),
    .Q_N(_11044_),
    .Q(\top_ihp.wb_emem.bit_counter[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1963),
    .D(_02450_),
    .Q_N(_11043_),
    .Q(\top_ihp.wb_emem.bit_counter[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1964),
    .D(_02451_),
    .Q_N(_11042_),
    .Q(\top_ihp.wb_emem.bit_counter[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[0]$_DFFE_NN0P_  (.CLK(net2095),
    .RESET_B(net1076),
    .D(_02452_),
    .Q_N(_11041_),
    .Q(\top_ihp.wb_dati_ram[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[10]$_DFFE_NN0P_  (.CLK(net2094),
    .RESET_B(net1061),
    .D(_02453_),
    .Q_N(_11040_),
    .Q(\top_ihp.wb_dati_ram[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[11]$_DFFE_NN0P_  (.CLK(net2093),
    .RESET_B(net1076),
    .D(_02454_),
    .Q_N(_11039_),
    .Q(\top_ihp.wb_dati_ram[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[12]$_DFFE_NN0P_  (.CLK(net2092),
    .RESET_B(net1076),
    .D(_02455_),
    .Q_N(_11038_),
    .Q(\top_ihp.wb_dati_ram[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[13]$_DFFE_NN0P_  (.CLK(net2091),
    .RESET_B(net1076),
    .D(_02456_),
    .Q_N(_11037_),
    .Q(\top_ihp.wb_dati_ram[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[14]$_DFFE_NN0P_  (.CLK(net2090),
    .RESET_B(net1076),
    .D(_02457_),
    .Q_N(_11036_),
    .Q(\top_ihp.wb_dati_ram[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[15]$_DFFE_NN0P_  (.CLK(net2089),
    .RESET_B(net1076),
    .D(_02458_),
    .Q_N(_11035_),
    .Q(\top_ihp.wb_dati_ram[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[16]$_DFFE_NN0P_  (.CLK(net2088),
    .RESET_B(net1068),
    .D(_02459_),
    .Q_N(_11034_),
    .Q(\top_ihp.wb_dati_ram[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[17]$_DFFE_NN0P_  (.CLK(net2087),
    .RESET_B(net1067),
    .D(_02460_),
    .Q_N(_11033_),
    .Q(\top_ihp.wb_dati_ram[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[18]$_DFFE_NN0P_  (.CLK(net2086),
    .RESET_B(net1067),
    .D(_02461_),
    .Q_N(_11032_),
    .Q(\top_ihp.wb_dati_ram[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[19]$_DFFE_NN0P_  (.CLK(net2085),
    .RESET_B(net1067),
    .D(_02462_),
    .Q_N(_11031_),
    .Q(\top_ihp.wb_dati_ram[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[1]$_DFFE_NN0P_  (.CLK(net2084),
    .RESET_B(net1053),
    .D(_02463_),
    .Q_N(_11030_),
    .Q(\top_ihp.wb_dati_ram[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[20]$_DFFE_NN0P_  (.CLK(net2083),
    .RESET_B(net1050),
    .D(_02464_),
    .Q_N(_11029_),
    .Q(\top_ihp.wb_dati_ram[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[21]$_DFFE_NN0P_  (.CLK(net2082),
    .RESET_B(net1050),
    .D(_02465_),
    .Q_N(_11028_),
    .Q(\top_ihp.wb_dati_ram[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[22]$_DFFE_NN0P_  (.CLK(net2081),
    .RESET_B(net1051),
    .D(_02466_),
    .Q_N(_11027_),
    .Q(\top_ihp.wb_dati_ram[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[23]$_DFFE_NN0P_  (.CLK(net2080),
    .RESET_B(net1061),
    .D(_02467_),
    .Q_N(_11026_),
    .Q(\top_ihp.wb_dati_ram[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[24]$_DFFE_NN0P_  (.CLK(net2079),
    .RESET_B(net1061),
    .D(_02468_),
    .Q_N(_11025_),
    .Q(\top_ihp.wb_dati_ram[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[25]$_DFFE_NN0P_  (.CLK(net2078),
    .RESET_B(net1061),
    .D(_02469_),
    .Q_N(_11024_),
    .Q(\top_ihp.wb_dati_ram[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[26]$_DFFE_NN0P_  (.CLK(net2077),
    .RESET_B(net1053),
    .D(_02470_),
    .Q_N(_11023_),
    .Q(\top_ihp.wb_dati_ram[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[27]$_DFFE_NN0P_  (.CLK(net2076),
    .RESET_B(net1053),
    .D(_02471_),
    .Q_N(_11022_),
    .Q(\top_ihp.wb_dati_ram[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[28]$_DFFE_NN0P_  (.CLK(net2075),
    .RESET_B(net1053),
    .D(_02472_),
    .Q_N(_11021_),
    .Q(\top_ihp.wb_dati_ram[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[29]$_DFFE_NN0P_  (.CLK(net2074),
    .RESET_B(net1051),
    .D(_02473_),
    .Q_N(_11020_),
    .Q(\top_ihp.wb_dati_ram[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[2]$_DFFE_NN0P_  (.CLK(net2073),
    .RESET_B(net1068),
    .D(_02474_),
    .Q_N(_11019_),
    .Q(\top_ihp.wb_dati_ram[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[30]$_DFFE_NN0P_  (.CLK(net2072),
    .RESET_B(net1053),
    .D(_02475_),
    .Q_N(_11018_),
    .Q(\top_ihp.wb_dati_ram[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[31]$_DFFE_NN0P_  (.CLK(net2071),
    .RESET_B(net1061),
    .D(_02476_),
    .Q_N(_11017_),
    .Q(\top_ihp.wb_dati_ram[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[32]$_DFFE_NN0P_  (.CLK(net2070),
    .RESET_B(net1064),
    .D(_02477_),
    .Q_N(_11016_),
    .Q(\top_ihp.wb_emem.cmd[32] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[33]$_DFFE_NN0P_  (.CLK(net2069),
    .RESET_B(net1064),
    .D(_02478_),
    .Q_N(_11015_),
    .Q(\top_ihp.wb_emem.cmd[33] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[34]$_DFFE_NN0P_  (.CLK(net2068),
    .RESET_B(net1061),
    .D(_02479_),
    .Q_N(_11014_),
    .Q(\top_ihp.wb_emem.cmd[34] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[35]$_DFFE_NN0P_  (.CLK(net2067),
    .RESET_B(net1062),
    .D(_02480_),
    .Q_N(_11013_),
    .Q(\top_ihp.wb_emem.cmd[35] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[36]$_DFFE_NN0P_  (.CLK(net2066),
    .RESET_B(net1063),
    .D(_02481_),
    .Q_N(_11012_),
    .Q(\top_ihp.wb_emem.cmd[36] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[37]$_DFFE_NN0P_  (.CLK(net2065),
    .RESET_B(net1063),
    .D(_02482_),
    .Q_N(_11011_),
    .Q(\top_ihp.wb_emem.cmd[37] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[38]$_DFFE_NN0P_  (.CLK(net2064),
    .RESET_B(net1057),
    .D(_02483_),
    .Q_N(_11010_),
    .Q(\top_ihp.wb_emem.cmd[38] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[39]$_DFFE_NN0P_  (.CLK(net2063),
    .RESET_B(net1057),
    .D(_02484_),
    .Q_N(_11009_),
    .Q(\top_ihp.wb_emem.cmd[39] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[3]$_DFFE_NN0P_  (.CLK(net2062),
    .RESET_B(net1068),
    .D(_02485_),
    .Q_N(_11008_),
    .Q(\top_ihp.wb_dati_ram[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[40]$_DFFE_NN0P_  (.CLK(net2061),
    .RESET_B(net1063),
    .D(_02486_),
    .Q_N(_11007_),
    .Q(\top_ihp.wb_emem.cmd[40] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[41]$_DFFE_NN0P_  (.CLK(net2060),
    .RESET_B(net1063),
    .D(_02487_),
    .Q_N(_11006_),
    .Q(\top_ihp.wb_emem.cmd[41] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[42]$_DFFE_NN0P_  (.CLK(net2059),
    .RESET_B(net1063),
    .D(_02488_),
    .Q_N(_11005_),
    .Q(\top_ihp.wb_emem.cmd[42] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[43]$_DFFE_NN0P_  (.CLK(net2058),
    .RESET_B(net1063),
    .D(_02489_),
    .Q_N(_11004_),
    .Q(\top_ihp.wb_emem.cmd[43] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[44]$_DFFE_NN0P_  (.CLK(net2057),
    .RESET_B(net1063),
    .D(_02490_),
    .Q_N(_11003_),
    .Q(\top_ihp.wb_emem.cmd[44] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[45]$_DFFE_NN0P_  (.CLK(net2056),
    .RESET_B(net1063),
    .D(_02491_),
    .Q_N(_11002_),
    .Q(\top_ihp.wb_emem.cmd[45] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[46]$_DFFE_NN0P_  (.CLK(net2055),
    .RESET_B(net1064),
    .D(_02492_),
    .Q_N(_11001_),
    .Q(\top_ihp.wb_emem.cmd[46] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[47]$_DFFE_NN0P_  (.CLK(net2054),
    .RESET_B(net1064),
    .D(_02493_),
    .Q_N(_11000_),
    .Q(\top_ihp.wb_emem.cmd[47] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[48]$_DFFE_NN1P_  (.CLK(net2053),
    .RESET_B(net1064),
    .D(_02494_),
    .Q_N(\top_ihp.wb_emem.cmd[48] ),
    .Q(_00214_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[49]$_DFFE_NN0P_  (.CLK(net2052),
    .RESET_B(net1065),
    .D(_02495_),
    .Q_N(_10999_),
    .Q(\top_ihp.wb_emem.cmd[49] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[4]$_DFFE_NN0P_  (.CLK(net2051),
    .RESET_B(net1054),
    .D(_02496_),
    .Q_N(_10998_),
    .Q(\top_ihp.wb_dati_ram[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[50]$_DFFE_NN0P_  (.CLK(net2050),
    .RESET_B(net1064),
    .D(_02497_),
    .Q_N(_10997_),
    .Q(\top_ihp.wb_emem.cmd[50] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[51]$_DFFE_NN1P_  (.CLK(net2049),
    .RESET_B(net1064),
    .D(_02498_),
    .Q_N(\top_ihp.wb_emem.cmd[51] ),
    .Q(_00215_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[52]$_DFFE_NN1P_  (.CLK(net2048),
    .RESET_B(net1087),
    .D(_02499_),
    .Q_N(\top_ihp.wb_emem.cmd[52] ),
    .Q(_00216_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[53]$_DFFE_NN0P_  (.CLK(net2047),
    .RESET_B(net1087),
    .D(_02500_),
    .Q_N(_10996_),
    .Q(\top_ihp.wb_emem.cmd[53] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[54]$_DFFE_NN0P_  (.CLK(net2046),
    .RESET_B(net1087),
    .D(_02501_),
    .Q_N(_10995_),
    .Q(\top_ihp.wb_emem.cmd[54] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[55]$_DFFE_NN1P_  (.CLK(net2045),
    .RESET_B(net1087),
    .D(_02502_),
    .Q_N(\top_ihp.wb_emem.cmd[55] ),
    .Q(_00217_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[56]$_DFFE_NN0P_  (.CLK(net2044),
    .RESET_B(net1062),
    .D(_02503_),
    .Q_N(_10994_),
    .Q(\top_ihp.wb_emem.cmd[56] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[57]$_DFFE_NN1P_  (.CLK(net2043),
    .RESET_B(net1057),
    .D(_02504_),
    .Q_N(\top_ihp.wb_emem.cmd[57] ),
    .Q(_00218_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[58]$_DFFE_NN1P_  (.CLK(net2042),
    .RESET_B(net1057),
    .D(_02505_),
    .Q_N(\top_ihp.wb_emem.cmd[58] ),
    .Q(_00219_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[59]$_DFFE_NN0P_  (.CLK(net2041),
    .RESET_B(net1057),
    .D(_02506_),
    .Q_N(_10993_),
    .Q(\top_ihp.wb_emem.cmd[59] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[5]$_DFFE_NN0P_  (.CLK(net2040),
    .RESET_B(net1054),
    .D(_02507_),
    .Q_N(_10992_),
    .Q(\top_ihp.wb_dati_ram[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[60]$_DFFE_NN0P_  (.CLK(net2039),
    .RESET_B(net1058),
    .D(_02508_),
    .Q_N(_10991_),
    .Q(\top_ihp.wb_emem.cmd[60] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[61]$_DFFE_NN1P_  (.CLK(net2038),
    .RESET_B(net1058),
    .D(_02509_),
    .Q_N(\top_ihp.wb_emem.cmd[61] ),
    .Q(_00220_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[62]$_DFFE_NN1P_  (.CLK(net2037),
    .RESET_B(net1058),
    .D(_02510_),
    .Q_N(\top_ihp.wb_emem.cmd[62] ),
    .Q(_00221_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[63]$_DFFE_NN0P_  (.CLK(net2036),
    .RESET_B(net1087),
    .D(_02511_),
    .Q_N(_10990_),
    .Q(\top_ihp.wb_emem.cmd[63] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[6]$_DFFE_NN0P_  (.CLK(net2035),
    .RESET_B(net1054),
    .D(_02512_),
    .Q_N(_10989_),
    .Q(\top_ihp.wb_dati_ram[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[7]$_DFFE_NN0P_  (.CLK(net2034),
    .RESET_B(net1061),
    .D(_02513_),
    .Q_N(_10988_),
    .Q(\top_ihp.wb_dati_ram[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[8]$_DFFE_NN0P_  (.CLK(net2033),
    .RESET_B(net1061),
    .D(_02514_),
    .Q_N(_10987_),
    .Q(\top_ihp.wb_dati_ram[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[9]$_DFFE_NN0P_  (.CLK(net2032),
    .RESET_B(net1062),
    .D(_02515_),
    .Q_N(_10986_),
    .Q(\top_ihp.wb_dati_ram[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.last_bit$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1965),
    .D(_02516_),
    .Q_N(_10985_),
    .Q(\top_ihp.wb_emem.last_bit ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.last_wait$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1966),
    .D(_02517_),
    .Q_N(_10984_),
    .Q(\top_ihp.wb_emem.last_wait ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[3]$_SDFFCE_NP1P_  (.CLK(net2031),
    .RESET_B(net1967),
    .D(_02518_),
    .Q_N(_10983_),
    .Q(\top_ihp.wb_emem.nbits[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[4]$_SDFFCE_NP0P_  (.CLK(net2030),
    .RESET_B(net1968),
    .D(_02519_),
    .Q_N(_10982_),
    .Q(\top_ihp.wb_emem.nbits[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[5]$_SDFFCE_NP0P_  (.CLK(net2029),
    .RESET_B(net1969),
    .D(_02520_),
    .Q_N(_10981_),
    .Q(\top_ihp.wb_emem.nbits[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[6]$_SDFFCE_NP0P_  (.CLK(net2028),
    .RESET_B(net1970),
    .D(_02521_),
    .Q_N(_10980_),
    .Q(\top_ihp.wb_emem.nbits[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[0]$_DFFE_NN0P_  (.CLK(net2027),
    .RESET_B(net1055),
    .D(_02522_),
    .Q_N(_10979_),
    .Q(\top_ihp.wb_emem.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[1]$_DFFE_NN0P_  (.CLK(net2026),
    .RESET_B(net1060),
    .D(_02523_),
    .Q_N(_10978_),
    .Q(\top_ihp.wb_emem.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[2]$_DFFE_NN0P_  (.CLK(net2025),
    .RESET_B(net1062),
    .D(_02524_),
    .Q_N(_10977_),
    .Q(\top_ihp.wb_emem.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[3]$_DFFE_NN0P_  (.CLK(net2024),
    .RESET_B(net1062),
    .D(_02525_),
    .Q_N(\top_ihp.ram_cs_o ),
    .Q(\top_ihp.wb_emem.state[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1971),
    .D(_02526_),
    .Q_N(_00139_),
    .Q(\top_ihp.wb_emem.wait_counter[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1972),
    .D(_02527_),
    .Q_N(_10976_),
    .Q(\top_ihp.wb_emem.wait_counter[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1973),
    .D(_02528_),
    .Q_N(_10975_),
    .Q(\top_ihp.wb_emem.wait_counter[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1974),
    .D(_02529_),
    .Q_N(_10974_),
    .Q(\top_ihp.wb_emem.wait_counter[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1975),
    .D(_02530_),
    .Q_N(_10973_),
    .Q(\top_ihp.wb_emem.wait_counter[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1976),
    .D(_02531_),
    .Q_N(_10972_),
    .Q(\top_ihp.wb_emem.wait_counter[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1977),
    .D(_02532_),
    .Q_N(_10971_),
    .Q(\top_ihp.wb_emem.wait_counter[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1978),
    .D(_02533_),
    .Q_N(_13134_),
    .Q(\top_ihp.wb_emem.wait_counter[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1096),
    .D(_00003_),
    .Q_N(_00072_),
    .Q(\top_ihp.wb_ack_gpio ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1102),
    .D(_02534_),
    .Q_N(_10970_),
    .Q(\top_ihp.wb_dati_gpio[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1099),
    .D(_02535_),
    .Q_N(_10969_),
    .Q(\top_ihp.gpio_o_1 ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1099),
    .D(_02536_),
    .Q_N(\top_ihp.gpio_o_2 ),
    .Q(_00222_));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1101),
    .D(_02537_),
    .Q_N(_10968_),
    .Q(\top_ihp.gpio_o_3 ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1093),
    .D(_02538_),
    .Q_N(\top_ihp.gpio_o_4 ),
    .Q(_00223_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[0]$_DFFE_NN0P_  (.CLK(net2023),
    .RESET_B(net1089),
    .D(_02539_),
    .Q_N(_10967_),
    .Q(\top_ihp.wb_imem.bits_left[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[1]$_DFFE_NN0P_  (.CLK(net2022),
    .RESET_B(net1089),
    .D(_02540_),
    .Q_N(_10966_),
    .Q(\top_ihp.wb_imem.bits_left[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[2]$_DFFE_NN0P_  (.CLK(net2021),
    .RESET_B(net1087),
    .D(_02541_),
    .Q_N(_10965_),
    .Q(\top_ihp.wb_imem.bits_left[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[3]$_DFFE_NN0P_  (.CLK(net2020),
    .RESET_B(net1087),
    .D(_02542_),
    .Q_N(_10964_),
    .Q(\top_ihp.wb_imem.bits_left[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[4]$_DFFE_NN0P_  (.CLK(net2019),
    .RESET_B(net1087),
    .D(_02543_),
    .Q_N(_10963_),
    .Q(\top_ihp.wb_imem.bits_left[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[5]$_DFFE_NN0P_  (.CLK(net2018),
    .RESET_B(net1088),
    .D(_02544_),
    .Q_N(_10962_),
    .Q(\top_ihp.wb_imem.bits_left[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[0]$_DFFE_NN0P_  (.CLK(net2017),
    .RESET_B(net1096),
    .D(_02545_),
    .Q_N(_10961_),
    .Q(\top_ihp.wb_dati_rom[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[10]$_DFFE_NN0P_  (.CLK(net2016),
    .RESET_B(net1088),
    .D(_02546_),
    .Q_N(_10960_),
    .Q(\top_ihp.wb_dati_rom[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[11]$_DFFE_NN0P_  (.CLK(net2015),
    .RESET_B(net1094),
    .D(_02547_),
    .Q_N(_10959_),
    .Q(\top_ihp.wb_dati_rom[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[12]$_DFFE_NN0P_  (.CLK(net2014),
    .RESET_B(net1077),
    .D(_02548_),
    .Q_N(_10958_),
    .Q(\top_ihp.wb_dati_rom[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[13]$_DFFE_NN0P_  (.CLK(net2013),
    .RESET_B(net1077),
    .D(_02549_),
    .Q_N(_10957_),
    .Q(\top_ihp.wb_dati_rom[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[14]$_DFFE_NN0P_  (.CLK(net2012),
    .RESET_B(net1077),
    .D(_02550_),
    .Q_N(_10956_),
    .Q(\top_ihp.wb_dati_rom[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[15]$_DFFE_NN0P_  (.CLK(net2011),
    .RESET_B(net1077),
    .D(_02551_),
    .Q_N(_10955_),
    .Q(\top_ihp.wb_dati_rom[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[16]$_DFFE_NN0P_  (.CLK(net2010),
    .RESET_B(net1077),
    .D(_02552_),
    .Q_N(_10954_),
    .Q(\top_ihp.wb_dati_rom[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[17]$_DFFE_NN0P_  (.CLK(net2009),
    .RESET_B(net1077),
    .D(_02553_),
    .Q_N(_10953_),
    .Q(\top_ihp.wb_dati_rom[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[18]$_DFFE_NN0P_  (.CLK(net2008),
    .RESET_B(net1065),
    .D(_02554_),
    .Q_N(_10952_),
    .Q(\top_ihp.wb_dati_rom[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[19]$_DFFE_NN0P_  (.CLK(net2007),
    .RESET_B(net1088),
    .D(_02555_),
    .Q_N(_10951_),
    .Q(\top_ihp.wb_dati_rom[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[1]$_DFFE_NN0P_  (.CLK(net2006),
    .RESET_B(net1094),
    .D(_02556_),
    .Q_N(_10950_),
    .Q(\top_ihp.wb_dati_rom[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[20]$_DFFE_NN0P_  (.CLK(net2005),
    .RESET_B(net1094),
    .D(_02557_),
    .Q_N(_10949_),
    .Q(\top_ihp.wb_dati_rom[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[21]$_DFFE_NN0P_  (.CLK(net2004),
    .RESET_B(net1094),
    .D(_02558_),
    .Q_N(_10948_),
    .Q(\top_ihp.wb_dati_rom[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[22]$_DFFE_NN0P_  (.CLK(net2003),
    .RESET_B(net1094),
    .D(_02559_),
    .Q_N(_10947_),
    .Q(\top_ihp.wb_dati_rom[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[23]$_DFFE_NN0P_  (.CLK(net2002),
    .RESET_B(net1094),
    .D(_02560_),
    .Q_N(_10946_),
    .Q(\top_ihp.wb_dati_rom[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[24]$_DFFE_NN0P_  (.CLK(net2001),
    .RESET_B(net1094),
    .D(_02561_),
    .Q_N(_10945_),
    .Q(\top_ihp.wb_dati_rom[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[25]$_DFFE_NN0P_  (.CLK(net2000),
    .RESET_B(net1094),
    .D(_02562_),
    .Q_N(_10944_),
    .Q(\top_ihp.wb_dati_rom[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[26]$_DFFE_NN0P_  (.CLK(net1999),
    .RESET_B(net1096),
    .D(_02563_),
    .Q_N(_10943_),
    .Q(\top_ihp.wb_dati_rom[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[27]$_DFFE_NN0P_  (.CLK(net1998),
    .RESET_B(net1096),
    .D(_02564_),
    .Q_N(_10942_),
    .Q(\top_ihp.wb_dati_rom[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[28]$_DFFE_NN0P_  (.CLK(net1997),
    .RESET_B(net1096),
    .D(_02565_),
    .Q_N(_10941_),
    .Q(\top_ihp.wb_dati_rom[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[29]$_DFFE_NN0P_  (.CLK(net1996),
    .RESET_B(net1089),
    .D(_02566_),
    .Q_N(_10940_),
    .Q(\top_ihp.wb_dati_rom[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[2]$_DFFE_NN0P_  (.CLK(net1995),
    .RESET_B(net1077),
    .D(_02567_),
    .Q_N(_10939_),
    .Q(\top_ihp.wb_dati_rom[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[30]$_DFFE_NN0P_  (.CLK(net1994),
    .RESET_B(net1090),
    .D(_02568_),
    .Q_N(_10938_),
    .Q(\top_ihp.wb_dati_rom[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[31]$_DFFE_NN0P_  (.CLK(net1993),
    .RESET_B(net1090),
    .D(_02569_),
    .Q_N(_10937_),
    .Q(\top_ihp.wb_dati_rom[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[3]$_DFFE_NN0P_  (.CLK(net1992),
    .RESET_B(net1077),
    .D(_02570_),
    .Q_N(_10936_),
    .Q(\top_ihp.wb_dati_rom[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[4]$_DFFE_NN0P_  (.CLK(net1991),
    .RESET_B(net1078),
    .D(_02571_),
    .Q_N(_10935_),
    .Q(\top_ihp.wb_dati_rom[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[5]$_DFFE_NN0P_  (.CLK(net1990),
    .RESET_B(net1078),
    .D(_02572_),
    .Q_N(_10934_),
    .Q(\top_ihp.wb_dati_rom[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[6]$_DFFE_NN0P_  (.CLK(net1989),
    .RESET_B(net1065),
    .D(_02573_),
    .Q_N(_10933_),
    .Q(\top_ihp.wb_dati_rom[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[7]$_DFFE_NN0P_  (.CLK(net1988),
    .RESET_B(net1088),
    .D(_02574_),
    .Q_N(_10932_),
    .Q(\top_ihp.wb_dati_rom[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[8]$_DFFE_NN0P_  (.CLK(net1987),
    .RESET_B(net1088),
    .D(_02575_),
    .Q_N(_10931_),
    .Q(\top_ihp.wb_dati_rom[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[9]$_DFFE_NN0P_  (.CLK(net1986),
    .RESET_B(net1088),
    .D(_02576_),
    .Q_N(_10930_),
    .Q(\top_ihp.wb_dati_rom[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.spi_cs_o$_DFFE_NN1P_  (.CLK(net1985),
    .RESET_B(net1090),
    .D(_02577_),
    .Q_N(\top_ihp.rom_cs_o ),
    .Q(_00224_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[0]$_DFF_NN1_  (.CLK(net1984),
    .RESET_B(net1090),
    .D(_00229_),
    .Q_N(\top_ihp.wb_imem.state[0] ),
    .Q(_13206_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[1]$_DFF_NN0_  (.CLK(net1983),
    .RESET_B(net1088),
    .D(_00000_),
    .Q_N(_00077_),
    .Q(\top_ihp.wb_imem.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[2]$_DFF_NN0_  (.CLK(net1982),
    .RESET_B(net1090),
    .D(_00001_),
    .Q_N(_13135_),
    .Q(\top_ihp.wb_imem.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1078),
    .D(_13209_),
    .Q_N(_10929_),
    .Q(\top_ihp.wb_ack_spi ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1066),
    .D(_02578_),
    .Q_N(_10928_),
    .Q(\top_ihp.wb_spi.bits_left[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1070),
    .D(_02579_),
    .Q_N(_10927_),
    .Q(\top_ihp.wb_spi.bits_left[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1070),
    .D(_02580_),
    .Q_N(_10926_),
    .Q(\top_ihp.wb_spi.bits_left[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1070),
    .D(_02581_),
    .Q_N(_10925_),
    .Q(\top_ihp.wb_spi.bits_left[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1070),
    .D(_02582_),
    .Q_N(_10924_),
    .Q(\top_ihp.wb_spi.bits_left[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1070),
    .D(_02583_),
    .Q_N(_10923_),
    .Q(\top_ihp.wb_spi.bits_left[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1076),
    .D(_02584_),
    .Q_N(_10922_),
    .Q(\top_ihp.wb_dati_spi[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1068),
    .D(_02585_),
    .Q_N(_10921_),
    .Q(\top_ihp.wb_dati_spi[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1066),
    .D(_02586_),
    .Q_N(_10920_),
    .Q(\top_ihp.wb_dati_spi[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1069),
    .D(_02587_),
    .Q_N(_10919_),
    .Q(\top_ihp.wb_dati_spi[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1066),
    .D(_02588_),
    .Q_N(_10918_),
    .Q(\top_ihp.wb_dati_spi[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1069),
    .D(_02589_),
    .Q_N(_10917_),
    .Q(\top_ihp.wb_dati_spi[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1066),
    .D(_02590_),
    .Q_N(_10916_),
    .Q(\top_ihp.wb_dati_spi[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1066),
    .D(_02591_),
    .Q_N(_10915_),
    .Q(\top_ihp.wb_dati_spi[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1076),
    .D(_02592_),
    .Q_N(_10914_),
    .Q(\top_ihp.wb_dati_spi[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1079),
    .D(_02593_),
    .Q_N(_10913_),
    .Q(\top_ihp.wb_dati_spi[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1079),
    .D(_02594_),
    .Q_N(_10912_),
    .Q(\top_ihp.wb_dati_spi[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1068),
    .D(_02595_),
    .Q_N(_10911_),
    .Q(\top_ihp.wb_dati_spi[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1079),
    .D(_02596_),
    .Q_N(_10910_),
    .Q(\top_ihp.wb_dati_spi[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1080),
    .D(_02597_),
    .Q_N(_10909_),
    .Q(\top_ihp.wb_dati_spi[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1080),
    .D(_02598_),
    .Q_N(_10908_),
    .Q(\top_ihp.wb_dati_spi[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1080),
    .D(_02599_),
    .Q_N(_10907_),
    .Q(\top_ihp.wb_dati_spi[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1066),
    .D(_02600_),
    .Q_N(_10906_),
    .Q(\top_ihp.wb_dati_spi[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1066),
    .D(_02601_),
    .Q_N(_10905_),
    .Q(\top_ihp.wb_dati_spi[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1067),
    .D(_02602_),
    .Q_N(_10904_),
    .Q(\top_ihp.wb_dati_spi[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1067),
    .D(_02603_),
    .Q_N(_10903_),
    .Q(\top_ihp.wb_dati_spi[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1067),
    .D(_02604_),
    .Q_N(_10902_),
    .Q(\top_ihp.wb_dati_spi[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1067),
    .D(_02605_),
    .Q_N(_10901_),
    .Q(\top_ihp.wb_dati_spi[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1068),
    .D(_02606_),
    .Q_N(_10900_),
    .Q(\top_ihp.wb_dati_spi[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1067),
    .D(_02607_),
    .Q_N(_10899_),
    .Q(\top_ihp.wb_dati_spi[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1066),
    .D(_02608_),
    .Q_N(_10898_),
    .Q(\top_ihp.wb_dati_spi[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1068),
    .D(_02609_),
    .Q_N(_10897_),
    .Q(\top_ihp.wb_dati_spi[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1074),
    .D(_02610_),
    .Q_N(_10896_),
    .Q(\top_ihp.wb_dati_spi[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1074),
    .D(_02611_),
    .Q_N(_10895_),
    .Q(\top_ihp.wb_dati_spi[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1072),
    .D(_02612_),
    .Q_N(_10894_),
    .Q(\top_ihp.wb_dati_spi[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1072),
    .D(_02613_),
    .Q_N(_10893_),
    .Q(\top_ihp.wb_dati_spi[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1068),
    .D(_02614_),
    .Q_N(_10892_),
    .Q(\top_ihp.wb_dati_spi[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1069),
    .D(_02615_),
    .Q_N(_10891_),
    .Q(\top_ihp.wb_dati_spi[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_clk_cnt[0]$_DFF_NN0_  (.CLK(net1981),
    .RESET_B(net1099),
    .D(_10864_),
    .Q_N(_10864_),
    .Q(\top_ihp.wb_spi.spi_clk_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_clk_cnt[1]$_DFF_NN0_  (.CLK(net1980),
    .RESET_B(net1101),
    .D(_00140_),
    .Q_N(_10890_),
    .Q(\top_ihp.spi_clk_o ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_1$_DFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1083),
    .D(_02616_),
    .Q_N(\top_ihp.spi_cs_o_1 ),
    .Q(_00225_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_2$_DFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1083),
    .D(_02617_),
    .Q_N(\top_ihp.spi_cs_o_2 ),
    .Q(_00226_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_3$_DFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1083),
    .D(_02618_),
    .Q_N(\top_ihp.spi_cs_o_3 ),
    .Q(_00227_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.state$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1079),
    .D(_13210_),
    .Q_N(_00078_),
    .Q(\top_ihp.wb_spi.state ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.ack_o$_SDFFCE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1979),
    .D(_02619_),
    .Q_N(_00071_),
    .Q(\top_ihp.wb_ack_uart ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.state[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1089),
    .D(_02620_),
    .Q_N(_10889_),
    .Q(\top_ihp.wb_uart.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1089),
    .D(_02621_),
    .Q_N(_10888_),
    .Q(\top_ihp.wb_uart.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1083),
    .D(_02622_),
    .Q_N(_00089_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1083),
    .D(_02623_),
    .Q_N(_10887_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1083),
    .D(_02624_),
    .Q_N(_10886_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(_02625_),
    .Q_N(_13136_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_00004_),
    .Q_N(_13137_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1056),
    .D(_00005_),
    .Q_N(_13138_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1058),
    .D(_00006_),
    .Q_N(_13139_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1058),
    .D(_00007_),
    .Q_N(_13140_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1057),
    .D(_00008_),
    .Q_N(_13141_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1057),
    .D(_00009_),
    .Q_N(_13142_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1057),
    .D(_00010_),
    .Q_N(_13143_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[16]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1060),
    .D(_00011_),
    .Q_N(_13144_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[17]$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1055),
    .D(_00012_),
    .Q_N(_13145_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[18]$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1055),
    .D(_00013_),
    .Q_N(_13146_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[19]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1056),
    .D(_00014_),
    .Q_N(_13147_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1084),
    .D(_00015_),
    .Q_N(_13148_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[20]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1056),
    .D(_00016_),
    .Q_N(_13149_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[21]$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1055),
    .D(_00017_),
    .Q_N(_13150_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[22]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1055),
    .D(_00018_),
    .Q_N(_13151_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[23]$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1055),
    .D(_00019_),
    .Q_N(_13152_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[24]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1055),
    .D(_00020_),
    .Q_N(_13153_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[25]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1056),
    .D(_00021_),
    .Q_N(_13154_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[26]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1055),
    .D(_00022_),
    .Q_N(_13155_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[27]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1056),
    .D(_00023_),
    .Q_N(_13156_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[28]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1056),
    .D(_00024_),
    .Q_N(_13157_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[29]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1056),
    .D(_00025_),
    .Q_N(_13158_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1083),
    .D(_00026_),
    .Q_N(_13159_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[30]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1056),
    .D(_00027_),
    .Q_N(_13160_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[31]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1059),
    .D(_00028_),
    .Q_N(_13161_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1083),
    .D(_00029_),
    .Q_N(_13162_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1084),
    .D(_00030_),
    .Q_N(_13163_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_00031_),
    .Q_N(_00079_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_00032_),
    .Q_N(_13164_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_00033_),
    .Q_N(_13165_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1084),
    .D(_00034_),
    .Q_N(_13166_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1084),
    .D(_00035_),
    .Q_N(_10885_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(_02626_),
    .Q_N(_10884_),
    .Q(\top_ihp.wb_dati_uart[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1086),
    .D(_02627_),
    .Q_N(_10883_),
    .Q(\top_ihp.wb_dati_uart[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1089),
    .D(_02628_),
    .Q_N(_10882_),
    .Q(\top_ihp.wb_dati_uart[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1089),
    .D(_02629_),
    .Q_N(_10881_),
    .Q(\top_ihp.wb_dati_uart[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(_02630_),
    .Q_N(_10880_),
    .Q(\top_ihp.wb_dati_uart[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1085),
    .D(_02631_),
    .Q_N(_10879_),
    .Q(\top_ihp.wb_dati_uart[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1086),
    .D(_02632_),
    .Q_N(_10878_),
    .Q(\top_ihp.wb_dati_uart[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1086),
    .D(_02633_),
    .Q_N(_10877_),
    .Q(\top_ihp.wb_dati_uart[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data_ready$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(_02634_),
    .Q_N(_13167_),
    .Q(\top_ihp.wb_uart.rx_ready ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[0]$_DFF_PN0_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(\top_ihp.wb_uart.uart_rx.next_state[0] ),
    .Q_N(_13168_),
    .Q(\top_ihp.wb_uart.uart_rx.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(\top_ihp.wb_uart.uart_rx.next_state[1] ),
    .Q_N(_13169_),
    .Q(\top_ihp.wb_uart.uart_rx.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1085),
    .D(\top_ihp.wb_uart.uart_rx.next_state[2] ),
    .Q_N(_00080_),
    .Q(\top_ihp.wb_uart.uart_rx.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1052),
    .D(_02635_),
    .Q_N(_10876_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1052),
    .D(_02636_),
    .Q_N(_10875_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1052),
    .D(_02637_),
    .Q_N(_00090_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1052),
    .D(_02638_),
    .Q_N(_13170_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1045),
    .D(_00036_),
    .Q_N(_13171_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1048),
    .D(_00037_),
    .Q_N(_13172_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1048),
    .D(_00038_),
    .Q_N(_13173_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1048),
    .D(_00039_),
    .Q_N(_13174_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1048),
    .D(_00040_),
    .Q_N(_13175_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1048),
    .D(_00041_),
    .Q_N(_13176_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1048),
    .D(_00042_),
    .Q_N(_13177_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[16]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1048),
    .D(_00043_),
    .Q_N(_13178_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[17]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1048),
    .D(_00044_),
    .Q_N(_13179_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[18]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1049),
    .D(_00045_),
    .Q_N(_13180_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[19]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1049),
    .D(_00046_),
    .Q_N(_13181_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1045),
    .D(_00047_),
    .Q_N(_13182_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[20]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1049),
    .D(_00048_),
    .Q_N(_13183_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[21]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1049),
    .D(_00049_),
    .Q_N(_13184_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[22]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1046),
    .D(_00050_),
    .Q_N(_13185_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[23]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1046),
    .D(_00051_),
    .Q_N(_13186_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[24]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1047),
    .D(_00052_),
    .Q_N(_13187_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[25]$_DFF_PN0_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1047),
    .D(_00053_),
    .Q_N(_13188_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[26]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1046),
    .D(_00054_),
    .Q_N(_13189_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[27]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1046),
    .D(_00055_),
    .Q_N(_13190_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[28]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1046),
    .D(_00056_),
    .Q_N(_13191_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[29]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1046),
    .D(_00057_),
    .Q_N(_13192_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1045),
    .D(_00058_),
    .Q_N(_13193_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[30]$_DFF_PN0_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1046),
    .D(_00059_),
    .Q_N(_13194_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[31]$_DFF_PN0_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1046),
    .D(_00060_),
    .Q_N(_13195_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1045),
    .D(_00061_),
    .Q_N(_13196_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1045),
    .D(_00062_),
    .Q_N(_13197_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1045),
    .D(_00063_),
    .Q_N(_13198_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1045),
    .D(_00064_),
    .Q_N(_13199_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1045),
    .D(_00065_),
    .Q_N(_13200_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1047),
    .D(_00066_),
    .Q_N(_13201_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1047),
    .D(_00067_),
    .Q_N(_13202_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.state[0]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1052),
    .D(\top_ihp.wb_uart.uart_tx.next_state[0] ),
    .Q_N(_13203_),
    .Q(\top_ihp.wb_uart.uart_tx.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1052),
    .D(\top_ihp.wb_uart.uart_tx.next_state[1] ),
    .Q_N(_10874_),
    .Q(\top_ihp.wb_uart.uart_tx.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1050),
    .D(_02639_),
    .Q_N(_10873_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1051),
    .D(_02640_),
    .Q_N(_10872_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1050),
    .D(_02641_),
    .Q_N(_10871_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1051),
    .D(_02642_),
    .Q_N(_10870_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1050),
    .D(_02643_),
    .Q_N(_10869_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1050),
    .D(_02644_),
    .Q_N(_10868_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1050),
    .D(_02645_),
    .Q_N(_10867_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1050),
    .D(_02646_),
    .Q_N(_10866_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_ready$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1052),
    .D(_02647_),
    .Q_N(_10865_),
    .Q(\top_ihp.wb_uart.tx_ready ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_reg$_DFF_PN1_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1052),
    .D(_00230_),
    .Q_N(\top_ihp.tx ),
    .Q(_13207_));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[6]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[7]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout25 (.A(_03108_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_03053_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_02709_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_02693_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_02670_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_02668_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_02652_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_10855_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_10831_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_10495_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_10457_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_10455_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_10441_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_10429_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_10404_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_09981_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_03145_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_03106_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_03094_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_03092_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_03090_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_03078_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_02718_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_02655_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_02650_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_02648_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_10848_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_10846_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_10443_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_10439_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_10437_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_10422_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_10420_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_10203_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_10117_),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(_10088_));
 sg13g2_buf_2 fanout61 (.A(_10087_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_10084_),
    .X(net62));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(_10081_));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(_10074_));
 sg13g2_buf_4 fanout65 (.X(net65),
    .A(_10063_));
 sg13g2_buf_2 fanout66 (.A(_09944_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_09930_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_09914_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_09762_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_09714_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_09703_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_09599_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_09375_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_09270_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_06169_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_05538_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_05354_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_05210_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_05101_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_04811_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_03658_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_03639_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_03611_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03598_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_03216_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_03203_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_03190_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_03150_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_03118_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_03088_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_03083_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_03073_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_03071_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_03069_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03065_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_02753_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_02714_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_02712_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_02707_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_02697_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_02685_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_02680_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_02664_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_02662_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_10862_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_10859_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_10850_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_10841_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_10838_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_10811_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_10799_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_10767_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_10753_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_10686_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_10673_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_10540_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_10500_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_10498_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_10493_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_10473_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_10468_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_10452_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_10450_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_10435_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_10433_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_10424_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_10416_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_10413_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_10214_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_10163_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_10130_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_10122_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_10083_),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_10079_));
 sg13g2_buf_2 fanout135 (.A(_10071_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_10070_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_10032_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_09986_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_09782_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_09724_),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(_09702_));
 sg13g2_buf_2 fanout142 (.A(_09679_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_09623_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_09483_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_09462_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_09437_),
    .X(net146));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(_09374_));
 sg13g2_buf_2 fanout148 (.A(_09304_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_08140_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_08115_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_08093_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_06065_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_05211_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_05105_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_03614_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_03601_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_03599_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_03597_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_03530_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_03517_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_03374_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03361_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03304_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03301_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03292_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03289_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_03280_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_03279_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_03218_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03206_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_03204_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03202_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_03168_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03148_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_03143_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_03123_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_03103_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_03101_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_03086_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_03061_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_02987_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_02974_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_02864_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02851_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_02740_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_02727_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_02666_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_10807_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_10793_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_10769_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_10762_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_10756_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_10754_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_10752_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_10718_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_10711_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_10688_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_10676_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_10674_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_10672_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_10639_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_10568_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_10555_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_10549_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_10525_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_10512_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_10427_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_10408_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_10189_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_10107_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_10086_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_10085_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_10078_),
    .X(net213));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_10077_));
 sg13g2_buf_2 fanout215 (.A(_10072_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_10068_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_10066_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_10064_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_10061_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_10048_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_10047_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_10044_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_10038_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_10036_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_10027_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_10020_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_10015_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_10014_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_09995_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_09994_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_09978_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_09977_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_09966_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_09965_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_09895_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_09872_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_09841_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_09808_),
    .X(net238));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(_09781_));
 sg13g2_buf_2 fanout240 (.A(_09754_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_09669_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_09654_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_09643_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_09622_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_09573_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_09512_),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_09436_));
 sg13g2_buf_2 fanout248 (.A(_09419_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_09404_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_09348_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_09303_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_08008_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_07983_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_07963_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_05758_),
    .X(net255));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(_05334_));
 sg13g2_buf_2 fanout257 (.A(_05321_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_05320_),
    .X(net258));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_05307_));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_05300_));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_05294_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_05224_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_05219_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_05193_));
 sg13g2_buf_2 fanout265 (.A(_05191_),
    .X(net265));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_05189_));
 sg13g2_buf_2 fanout267 (.A(_05170_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_05114_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_05110_),
    .X(net269));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_05107_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_05090_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_05073_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_05037_));
 sg13g2_buf_2 fanout274 (.A(_03665_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_03651_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_03636_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_03578_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_03572_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_03563_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_03558_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_03557_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_03533_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_03520_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_03518_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_03516_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_03492_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_03479_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_03462_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_03457_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_03446_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_03440_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_03439_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_03422_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_03417_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_03406_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_03400_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_03399_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_03376_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_03364_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_03362_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_03360_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_03341_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_03335_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_03326_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_03321_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_03320_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_03254_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_03241_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_03182_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_03165_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_03163_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_03159_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_03084_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_03079_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_03062_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_03057_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_03037_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_03032_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_03021_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_03015_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_03014_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_02989_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_02977_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_02975_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_02973_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_02946_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_02933_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_02905_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_02892_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_02867_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_02854_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_02852_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_02850_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_02845_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_02824_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_02811_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_02742_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_02730_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_02728_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_02726_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_02704_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_02699_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_02686_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_02678_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_02677_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_02674_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_02653_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_10860_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_10843_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_10835_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_10834_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_10809_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_10796_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_10794_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_10792_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_10733_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_10715_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_10714_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_10709_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_10653_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_10636_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_10634_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_10630_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_10607_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_10594_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_10570_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_10558_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_10556_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_10554_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_10528_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_10515_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_10513_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_10511_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_10490_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_10485_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_10474_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_10466_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_10465_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_10430_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_10426_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_10411_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_10409_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_10407_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_10381_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_10377_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_10369_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_10364_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_10363_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_10342_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_10337_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_10328_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_10324_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_10323_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_10250_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_10237_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_10181_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_10180_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_10169_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_10168_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_10156_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_10155_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_10097_),
    .X(net402));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(_10082_));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_10067_));
 sg13g2_buf_2 fanout405 (.A(_10060_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_10035_),
    .X(net406));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_09946_));
 sg13g2_buf_2 fanout408 (.A(_09910_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_09554_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_09514_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_09204_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_09199_),
    .X(net412));
 sg13g2_buf_4 fanout413 (.X(net413),
    .A(_05760_));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(_05707_));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(_05597_));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(_05591_));
 sg13g2_buf_2 fanout417 (.A(_05590_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_05547_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_05485_),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(_05481_));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_05467_));
 sg13g2_buf_2 fanout422 (.A(_05462_),
    .X(net422));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(_05401_));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(_05383_));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(_05380_));
 sg13g2_buf_2 fanout426 (.A(_05377_),
    .X(net426));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(_05367_));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(_05345_));
 sg13g2_buf_2 fanout429 (.A(_05342_),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(_05310_));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(_05302_));
 sg13g2_buf_2 fanout432 (.A(_05290_),
    .X(net432));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_05255_));
 sg13g2_buf_4 fanout434 (.X(net434),
    .A(_05226_));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(_05221_));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(_05217_));
 sg13g2_buf_2 fanout437 (.A(_05215_),
    .X(net437));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(_05192_));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(_05188_));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_05180_));
 sg13g2_buf_2 fanout441 (.A(_05179_),
    .X(net441));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(_05177_));
 sg13g2_buf_2 fanout443 (.A(_05173_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_05171_),
    .X(net444));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(_05164_));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(_05116_));
 sg13g2_buf_2 fanout447 (.A(_05112_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_05109_),
    .X(net448));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(_05094_));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(_05089_));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(_05086_));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(_05080_));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(_05077_));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(_05072_));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(_05068_));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(_05059_));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(_05055_));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(_05044_));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(_05036_));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(_05028_));
 sg13g2_buf_2 fanout461 (.A(_04995_),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(_04989_));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(_04966_));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_04949_));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_04941_));
 sg13g2_buf_2 fanout466 (.A(_04937_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_04927_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_04921_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_04909_),
    .X(net469));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(_04903_));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(_04899_));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_04894_));
 sg13g2_buf_2 fanout473 (.A(_04890_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_04876_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_04871_),
    .X(net475));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(_04844_));
 sg13g2_buf_2 fanout477 (.A(_04827_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_03556_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_03554_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_03494_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_03482_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_03480_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_03478_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_03396_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_03319_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_03257_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_03244_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_03242_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_03240_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_03158_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_03140_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_03135_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_03124_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_03116_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_03115_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_03075_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_03058_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_03056_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_03011_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_02948_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_02936_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_02934_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_02932_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_02908_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_02895_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_02893_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_02891_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_02826_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_02814_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_02812_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_02810_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_02793_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_02788_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_02777_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_02771_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_02770_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_10852_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_10830_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_10629_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_10609_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_10597_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_10595_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_10593_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_10462_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_10362_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_10322_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_10278_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_10253_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_10240_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_10238_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_10236_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_10215_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_10211_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_10201_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_10197_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_10138_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_10133_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_10120_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_10113_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_10112_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_10109_),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_10103_));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_10100_));
 sg13g2_buf_2 fanout544 (.A(_10096_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_10029_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_09600_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_09553_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_09305_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_09271_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_09203_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_08090_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_05705_),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(_05620_));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_05520_));
 sg13g2_buf_2 fanout555 (.A(_05514_),
    .X(net555));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_05474_));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(_05472_));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_05460_));
 sg13g2_buf_2 fanout559 (.A(_05424_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_05398_),
    .X(net560));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_05393_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_05361_));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(_05359_));
 sg13g2_buf_2 fanout564 (.A(_05344_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_05329_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_05309_),
    .X(net566));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(_05299_));
 sg13g2_buf_2 fanout568 (.A(_05297_),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_05276_));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_05268_));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(_05266_));
 sg13g2_buf_2 fanout572 (.A(_05264_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_05250_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_05238_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_05214_),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_05201_));
 sg13g2_buf_2 fanout577 (.A(_05196_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_05185_),
    .X(net578));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(_05183_));
 sg13g2_buf_2 fanout580 (.A(_05182_),
    .X(net580));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(_05174_));
 sg13g2_buf_2 fanout582 (.A(_05166_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_05158_),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(_05154_));
 sg13g2_buf_2 fanout585 (.A(_05150_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_05144_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_05142_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_05131_),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_05115_));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(_05097_));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(_05067_));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(_05062_));
 sg13g2_buf_2 fanout593 (.A(_05052_),
    .X(net593));
 sg13g2_buf_4 fanout594 (.X(net594),
    .A(_05047_));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(_05040_));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_05031_));
 sg13g2_buf_2 fanout597 (.A(_05022_),
    .X(net597));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(_05016_));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_05012_));
 sg13g2_buf_2 fanout600 (.A(_05009_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_05004_),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_04999_));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(_04984_));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(_04979_));
 sg13g2_buf_4 fanout605 (.X(net605),
    .A(_04975_));
 sg13g2_buf_2 fanout606 (.A(_04970_),
    .X(net606));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(_04940_));
 sg13g2_buf_2 fanout608 (.A(_04936_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_04926_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_04920_),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(_04908_));
 sg13g2_buf_2 fanout612 (.A(_04902_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_04893_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_04889_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_04870_),
    .X(net615));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(_04866_));
 sg13g2_buf_2 fanout617 (.A(_04847_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_04821_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_04817_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_04562_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_04366_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_04356_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_04336_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_04319_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_04299_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_04297_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_04221_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_04172_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_03436_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_03316_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_03112_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_02767_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_10304_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_10299_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_10288_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_10282_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_10281_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_10198_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_10196_),
    .X(net639));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_05655_));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(_05464_));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(_05412_));
 sg13g2_buf_2 fanout643 (.A(_05409_),
    .X(net643));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(_05282_));
 sg13g2_buf_2 fanout645 (.A(_05204_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_05200_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_05146_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_05141_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_05139_),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(_05135_));
 sg13g2_buf_2 fanout651 (.A(_05019_),
    .X(net651));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(_04931_));
 sg13g2_buf_2 fanout653 (.A(_04925_),
    .X(net653));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(_04911_));
 sg13g2_buf_2 fanout655 (.A(_04888_),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(_04877_));
 sg13g2_buf_2 fanout657 (.A(_04846_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_04834_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_04227_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_04182_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_04171_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_04169_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_10398_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_10318_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_10151_),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(_05326_));
 sg13g2_buf_2 fanout667 (.A(_05281_),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_05280_));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_05134_));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(_05132_));
 sg13g2_buf_2 fanout671 (.A(_05127_),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(_05122_));
 sg13g2_buf_2 fanout673 (.A(_05083_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_04992_),
    .X(net674));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_04959_));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_04953_));
 sg13g2_buf_2 fanout677 (.A(_04944_),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_04910_));
 sg13g2_buf_2 fanout679 (.A(_04896_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_04873_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_04777_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_10460_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_07024_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_06853_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_06228_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_05653_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_05418_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_05272_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_05130_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_05126_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_05017_),
    .X(net691));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(_04958_));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(_04952_));
 sg13g2_buf_2 fanout694 (.A(_04943_),
    .X(net694));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(_04917_));
 sg13g2_buf_2 fanout696 (.A(_04878_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_04837_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_04829_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_04828_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_04818_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_04814_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_04813_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_04812_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_04792_));
 sg13g2_buf_2 fanout705 (.A(_04789_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_04776_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_04580_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_04552_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_03692_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_10092_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_09960_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_07027_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_07011_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_07005_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_06960_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_06938_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_06927_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_05609_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_05119_),
    .X(net719));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(_04930_));
 sg13g2_buf_2 fanout721 (.A(_04916_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_04853_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_04767_),
    .X(net723));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(_04759_));
 sg13g2_buf_2 fanout725 (.A(_04754_),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(_04744_));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_04720_));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_04710_));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(_04678_));
 sg13g2_buf_2 fanout730 (.A(_04570_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_04567_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_04534_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_04533_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_03925_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_03691_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_09855_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_09104_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_08224_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_07047_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_07016_),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(_06988_));
 sg13g2_buf_2 fanout742 (.A(_06987_),
    .X(net742));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_06985_));
 sg13g2_buf_2 fanout744 (.A(_06984_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_06978_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_06976_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_06975_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_06967_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_06966_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_06951_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_06950_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_06945_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_06944_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_06942_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_06939_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_06932_),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(_06929_));
 sg13g2_buf_2 fanout758 (.A(_06928_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_06891_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_06886_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_06883_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_06875_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_05410_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_05202_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_04772_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_04571_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_04532_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_04332_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_03900_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_03892_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_03697_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_03690_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_03680_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_08246_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_08225_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_08223_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_07441_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_07152_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_07050_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_07046_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_07042_),
    .X(net781));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(_06998_));
 sg13g2_buf_2 fanout783 (.A(_06995_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_06993_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_06962_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_06957_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_06948_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_06947_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_06941_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_06936_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_06931_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_06902_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_06894_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_06878_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_06866_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_06857_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_04851_));
 sg13g2_buf_2 fanout798 (.A(_04547_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_04359_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_04327_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_04084_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_03843_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_03689_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_09332_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_08222_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_07658_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_07440_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_07031_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_06968_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_06935_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_06898_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_06856_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_04311_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_04206_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_04161_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_04083_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_03841_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_03816_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_03810_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_03807_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_09166_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_08942_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_08244_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_07657_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_07168_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_07038_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_06956_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_06855_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_04199_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_04160_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_03929_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_03921_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_03862_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_03857_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_03834_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_03814_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_03809_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_03802_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_09174_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_09165_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_09146_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_08974_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_08384_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_08254_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_08220_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_07758_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_06924_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_06906_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_04194_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_03885_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_03884_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_03852_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_03827_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_03821_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_03818_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_03815_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_03812_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_03805_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_09351_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_09307_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_09145_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_08206_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_07757_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_06923_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_06905_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_03804_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_09350_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_09337_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_09250_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_09210_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_09205_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_09141_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_09123_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_08522_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_08436_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_08426_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_07799_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_07756_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_07436_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_03737_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_03717_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_09321_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_09310_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_09274_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_09221_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_09188_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_09181_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_08605_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_08551_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_08506_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_08449_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_08442_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_08429_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_08391_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_08386_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_08364_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_08334_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_08332_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_08320_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_08314_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_08273_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_08268_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_08200_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_07620_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_03946_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_03933_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_03918_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_03733_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_03719_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_03716_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_03715_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_03683_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_09290_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_09248_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_09180_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_09169_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_09157_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_09144_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_08653_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_08622_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_08569_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_08510_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_08427_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_08423_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_08390_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_08369_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_08348_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_08344_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_08322_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_08321_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_08318_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_08313_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_08310_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_08304_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_08300_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_08283_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_08272_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_08267_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_08230_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_08169_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_04394_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_04344_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_04323_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_04320_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_04073_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_04012_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_03917_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_09294_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_09245_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_09168_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_09164_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_09156_),
    .X(net952));
 sg13g2_buf_1 fanout953 (.A(_09143_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_09138_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_09122_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_09110_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_08466_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_08465_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_08422_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_08394_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_08377_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_08372_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_08350_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_08343_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_08327_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_08317_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_08309_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_08306_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_08299_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_08295_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_08291_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_08290_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_08286_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_08277_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_08271_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_08266_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_08260_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_08257_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_08247_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_08218_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_08194_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_07678_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_07675_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_07648_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_07634_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_04333_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_04315_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_09240_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_09189_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_09163_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_09161_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_09152_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_09135_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_09118_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_09111_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_09109_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_09090_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_09071_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_08944_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_08538_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_08464_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_08435_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_08366_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_08324_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_08316_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_08305_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_08302_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_08281_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_08270_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_08265_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_08262_),
    .X(net1011));
 sg13g2_buf_1 fanout1012 (.A(_08211_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_08186_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_07674_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_07580_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_07423_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_07418_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_09136_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_09054_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_08274_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_08269_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_08261_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_08258_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_08042_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_07762_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_07715_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_07680_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_07679_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_07626_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_07614_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_07550_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_07547_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_07539_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_07525_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_07517_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_07510_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_07496_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_07490_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_07487_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_07482_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_07478_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_07459_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_07455_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_07445_),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(net1047));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1047));
 sg13g2_buf_2 fanout1047 (.A(net1054),
    .X(net1047));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(net1054));
 sg13g2_buf_2 fanout1049 (.A(net1054),
    .X(net1049));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(net1053));
 sg13g2_buf_2 fanout1051 (.A(net1053),
    .X(net1051));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(net1053));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1054));
 sg13g2_buf_2 fanout1054 (.A(net1082),
    .X(net1054));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(net1060));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(net1059));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(net1059));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_1 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_1 fanout1060 (.A(net1082),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(net1062));
 sg13g2_buf_2 fanout1062 (.A(net1065),
    .X(net1062));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1064));
 sg13g2_buf_4 fanout1064 (.X(net1064),
    .A(net1065));
 sg13g2_buf_2 fanout1065 (.A(net1082),
    .X(net1065));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net1069));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(net1069));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(net1069));
 sg13g2_buf_2 fanout1069 (.A(net1075),
    .X(net1069));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(net1075));
 sg13g2_buf_2 fanout1071 (.A(net1075),
    .X(net1071));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1074));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(net1074));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(net1075));
 sg13g2_buf_1 fanout1075 (.A(net1082),
    .X(net1075));
 sg13g2_buf_4 fanout1076 (.X(net1076),
    .A(net1079));
 sg13g2_buf_4 fanout1077 (.X(net1077),
    .A(net1078));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1079));
 sg13g2_buf_2 fanout1079 (.A(net1082),
    .X(net1079));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1081));
 sg13g2_buf_2 fanout1081 (.A(net1082),
    .X(net1081));
 sg13g2_buf_1 fanout1082 (.A(net1169),
    .X(net1082));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(net1086));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(net1086));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(net1086));
 sg13g2_buf_2 fanout1086 (.A(net1091),
    .X(net1086));
 sg13g2_buf_4 fanout1087 (.X(net1087),
    .A(net1088));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(net1091));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1091));
 sg13g2_buf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_1 fanout1091 (.A(net1093),
    .X(net1091));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(net1093));
 sg13g2_buf_1 fanout1093 (.A(net1106),
    .X(net1093));
 sg13g2_buf_4 fanout1094 (.X(net1094),
    .A(net1096));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_4 fanout1096 (.X(net1096),
    .A(net1097));
 sg13g2_buf_2 fanout1097 (.A(net1106),
    .X(net1097));
 sg13g2_buf_4 fanout1098 (.X(net1098),
    .A(net1101));
 sg13g2_buf_2 fanout1099 (.A(net1101),
    .X(net1099));
 sg13g2_buf_4 fanout1100 (.X(net1100),
    .A(net1101));
 sg13g2_buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_4 fanout1102 (.X(net1102),
    .A(net1106));
 sg13g2_buf_4 fanout1103 (.X(net1103),
    .A(net1104));
 sg13g2_buf_2 fanout1104 (.A(net1105),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_1 fanout1106 (.A(net1169),
    .X(net1106));
 sg13g2_buf_4 fanout1107 (.X(net1107),
    .A(net1108));
 sg13g2_buf_2 fanout1108 (.A(net1118),
    .X(net1108));
 sg13g2_buf_4 fanout1109 (.X(net1109),
    .A(net1111));
 sg13g2_buf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(net1118),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(net1113));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(net1118));
 sg13g2_buf_4 fanout1114 (.X(net1114),
    .A(net1117));
 sg13g2_buf_4 fanout1115 (.X(net1115),
    .A(net1117));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(net1138),
    .X(net1118));
 sg13g2_buf_4 fanout1119 (.X(net1119),
    .A(net1123));
 sg13g2_buf_2 fanout1120 (.A(net1123),
    .X(net1120));
 sg13g2_buf_4 fanout1121 (.X(net1121),
    .A(net1123));
 sg13g2_buf_4 fanout1122 (.X(net1122),
    .A(net1123));
 sg13g2_buf_1 fanout1123 (.A(net1128),
    .X(net1123));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(net1125));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(net1128));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(net1128));
 sg13g2_buf_2 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_1 fanout1128 (.A(net1138),
    .X(net1128));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(net1132));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(net1132));
 sg13g2_buf_2 fanout1131 (.A(net1132),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(net1138),
    .X(net1132));
 sg13g2_buf_4 fanout1133 (.X(net1133),
    .A(net1137));
 sg13g2_buf_2 fanout1134 (.A(net1137),
    .X(net1134));
 sg13g2_buf_4 fanout1135 (.X(net1135),
    .A(net1137));
 sg13g2_buf_2 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_1 fanout1138 (.A(net1169),
    .X(net1138));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(net1143));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(net1143));
 sg13g2_buf_2 fanout1141 (.A(net1143),
    .X(net1141));
 sg13g2_buf_4 fanout1142 (.X(net1142),
    .A(net1143));
 sg13g2_buf_2 fanout1143 (.A(net1168),
    .X(net1143));
 sg13g2_buf_4 fanout1144 (.X(net1144),
    .A(net1145));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(net1168));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1148));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(net1148));
 sg13g2_buf_2 fanout1148 (.A(net1168),
    .X(net1148));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(net1152));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(net1152));
 sg13g2_buf_2 fanout1151 (.A(net1152),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(net1167),
    .X(net1152));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(net1157));
 sg13g2_buf_2 fanout1154 (.A(net1157),
    .X(net1154));
 sg13g2_buf_4 fanout1155 (.X(net1155),
    .A(net1157));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(net1157));
 sg13g2_buf_1 fanout1157 (.A(net1167),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1161));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(net1161));
 sg13g2_buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(net1167),
    .X(net1161));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(net1166));
 sg13g2_buf_2 fanout1163 (.A(net1166),
    .X(net1163));
 sg13g2_buf_4 fanout1164 (.X(net1164),
    .A(net1165));
 sg13g2_buf_4 fanout1165 (.X(net1165),
    .A(net1166));
 sg13g2_buf_1 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_1 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_1 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_buf_1 fanout1169 (.A(net1),
    .X(net1169));
 sg13g2_buf_4 fanout1170 (.X(net1170),
    .A(net1173));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(net1173));
 sg13g2_buf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_1 fanout1173 (.A(net1190),
    .X(net1173));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(net1179));
 sg13g2_buf_2 fanout1175 (.A(net1179),
    .X(net1175));
 sg13g2_buf_4 fanout1176 (.X(net1176),
    .A(net1179));
 sg13g2_buf_2 fanout1177 (.A(net1178),
    .X(net1177));
 sg13g2_buf_4 fanout1178 (.X(net1178),
    .A(net1179));
 sg13g2_buf_1 fanout1179 (.A(net1190),
    .X(net1179));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(net1184));
 sg13g2_buf_4 fanout1181 (.X(net1181),
    .A(net1184));
 sg13g2_buf_4 fanout1182 (.X(net1182),
    .A(net1184));
 sg13g2_buf_2 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_1 fanout1184 (.A(net1190),
    .X(net1184));
 sg13g2_buf_4 fanout1185 (.X(net1185),
    .A(net1186));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(net1189));
 sg13g2_buf_4 fanout1187 (.X(net1187),
    .A(net1188));
 sg13g2_buf_4 fanout1188 (.X(net1188),
    .A(net1189));
 sg13g2_buf_2 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_1 fanout1190 (.A(net1394),
    .X(net1190));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(net1194));
 sg13g2_buf_4 fanout1192 (.X(net1192),
    .A(net1194));
 sg13g2_buf_2 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(net1208),
    .X(net1194));
 sg13g2_buf_4 fanout1195 (.X(net1195),
    .A(net1198));
 sg13g2_buf_4 fanout1196 (.X(net1196),
    .A(net1198));
 sg13g2_buf_2 fanout1197 (.A(net1198),
    .X(net1197));
 sg13g2_buf_1 fanout1198 (.A(net1208),
    .X(net1198));
 sg13g2_buf_4 fanout1199 (.X(net1199),
    .A(net1203));
 sg13g2_buf_2 fanout1200 (.A(net1203),
    .X(net1200));
 sg13g2_buf_4 fanout1201 (.X(net1201),
    .A(net1203));
 sg13g2_buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_1 fanout1203 (.A(net1208),
    .X(net1203));
 sg13g2_buf_4 fanout1204 (.X(net1204),
    .A(net1207));
 sg13g2_buf_4 fanout1205 (.X(net1205),
    .A(net1207));
 sg13g2_buf_2 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_2 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_1 fanout1208 (.A(net1222),
    .X(net1208));
 sg13g2_buf_4 fanout1209 (.X(net1209),
    .A(net1210));
 sg13g2_buf_4 fanout1210 (.X(net1210),
    .A(net1214));
 sg13g2_buf_2 fanout1211 (.A(net1214),
    .X(net1211));
 sg13g2_buf_4 fanout1212 (.X(net1212),
    .A(net1213));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net1214));
 sg13g2_buf_2 fanout1214 (.A(net1222),
    .X(net1214));
 sg13g2_buf_4 fanout1215 (.X(net1215),
    .A(net1218));
 sg13g2_buf_4 fanout1216 (.X(net1216),
    .A(net1218));
 sg13g2_buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(net1222),
    .X(net1218));
 sg13g2_buf_4 fanout1219 (.X(net1219),
    .A(net1221));
 sg13g2_buf_4 fanout1220 (.X(net1220),
    .A(net1221));
 sg13g2_buf_2 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_1 fanout1222 (.A(net1394),
    .X(net1222));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(net1227));
 sg13g2_buf_2 fanout1224 (.A(net1227),
    .X(net1224));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(net1227));
 sg13g2_buf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_1 fanout1227 (.A(net1271),
    .X(net1227));
 sg13g2_buf_4 fanout1228 (.X(net1228),
    .A(net1232));
 sg13g2_buf_2 fanout1229 (.A(net1232),
    .X(net1229));
 sg13g2_buf_4 fanout1230 (.X(net1230),
    .A(net1231));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1232));
 sg13g2_buf_1 fanout1232 (.A(net1271),
    .X(net1232));
 sg13g2_buf_4 fanout1233 (.X(net1233),
    .A(net1234));
 sg13g2_buf_4 fanout1234 (.X(net1234),
    .A(net1243));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(net1243));
 sg13g2_buf_2 fanout1236 (.A(net1243),
    .X(net1236));
 sg13g2_buf_4 fanout1237 (.X(net1237),
    .A(net1238));
 sg13g2_buf_4 fanout1238 (.X(net1238),
    .A(net1242));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1241));
 sg13g2_buf_2 fanout1240 (.A(net1241),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_1 fanout1242 (.A(net1243),
    .X(net1242));
 sg13g2_buf_1 fanout1243 (.A(net1271),
    .X(net1243));
 sg13g2_buf_4 fanout1244 (.X(net1244),
    .A(net1246));
 sg13g2_buf_2 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(net1255),
    .X(net1246));
 sg13g2_buf_4 fanout1247 (.X(net1247),
    .A(net1248));
 sg13g2_buf_2 fanout1248 (.A(net1255),
    .X(net1248));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(net1251));
 sg13g2_buf_2 fanout1250 (.A(net1251),
    .X(net1250));
 sg13g2_buf_4 fanout1251 (.X(net1251),
    .A(net1255));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(net1254));
 sg13g2_buf_4 fanout1253 (.X(net1253),
    .A(net1254));
 sg13g2_buf_2 fanout1254 (.A(net1255),
    .X(net1254));
 sg13g2_buf_2 fanout1255 (.A(net1271),
    .X(net1255));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(net1257));
 sg13g2_buf_4 fanout1257 (.X(net1257),
    .A(net1263));
 sg13g2_buf_4 fanout1258 (.X(net1258),
    .A(net1262));
 sg13g2_buf_2 fanout1259 (.A(net1262),
    .X(net1259));
 sg13g2_buf_4 fanout1260 (.X(net1260),
    .A(net1262));
 sg13g2_buf_2 fanout1261 (.A(net1262),
    .X(net1261));
 sg13g2_buf_1 fanout1262 (.A(net1263),
    .X(net1262));
 sg13g2_buf_1 fanout1263 (.A(net1271),
    .X(net1263));
 sg13g2_buf_4 fanout1264 (.X(net1264),
    .A(net1265));
 sg13g2_buf_4 fanout1265 (.X(net1265),
    .A(net1270));
 sg13g2_buf_4 fanout1266 (.X(net1266),
    .A(net1269));
 sg13g2_buf_4 fanout1267 (.X(net1267),
    .A(net1269));
 sg13g2_buf_2 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_2 fanout1269 (.A(net1270),
    .X(net1269));
 sg13g2_buf_2 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_1 fanout1271 (.A(net1394),
    .X(net1271));
 sg13g2_buf_4 fanout1272 (.X(net1272),
    .A(net1276));
 sg13g2_buf_2 fanout1273 (.A(net1276),
    .X(net1273));
 sg13g2_buf_4 fanout1274 (.X(net1274),
    .A(net1276));
 sg13g2_buf_2 fanout1275 (.A(net1276),
    .X(net1275));
 sg13g2_buf_1 fanout1276 (.A(net1279),
    .X(net1276));
 sg13g2_buf_4 fanout1277 (.X(net1277),
    .A(net1279));
 sg13g2_buf_4 fanout1278 (.X(net1278),
    .A(net1279));
 sg13g2_buf_2 fanout1279 (.A(net1300),
    .X(net1279));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(net1283));
 sg13g2_buf_4 fanout1281 (.X(net1281),
    .A(net1283));
 sg13g2_buf_2 fanout1282 (.A(net1283),
    .X(net1282));
 sg13g2_buf_2 fanout1283 (.A(net1300),
    .X(net1283));
 sg13g2_buf_4 fanout1284 (.X(net1284),
    .A(net1286));
 sg13g2_buf_4 fanout1285 (.X(net1285),
    .A(net1286));
 sg13g2_buf_2 fanout1286 (.A(net1300),
    .X(net1286));
 sg13g2_buf_4 fanout1287 (.X(net1287),
    .A(net1289));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(net1289));
 sg13g2_buf_2 fanout1289 (.A(net1299),
    .X(net1289));
 sg13g2_buf_4 fanout1290 (.X(net1290),
    .A(net1291));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(net1299));
 sg13g2_buf_2 fanout1292 (.A(net1299),
    .X(net1292));
 sg13g2_buf_4 fanout1293 (.X(net1293),
    .A(net1295));
 sg13g2_buf_4 fanout1294 (.X(net1294),
    .A(net1295));
 sg13g2_buf_2 fanout1295 (.A(net1299),
    .X(net1295));
 sg13g2_buf_4 fanout1296 (.X(net1296),
    .A(net1298));
 sg13g2_buf_4 fanout1297 (.X(net1297),
    .A(net1298));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_1 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_1 fanout1300 (.A(net1393),
    .X(net1300));
 sg13g2_buf_4 fanout1301 (.X(net1301),
    .A(net1305));
 sg13g2_buf_2 fanout1302 (.A(net1305),
    .X(net1302));
 sg13g2_buf_4 fanout1303 (.X(net1303),
    .A(net1305));
 sg13g2_buf_2 fanout1304 (.A(net1305),
    .X(net1304));
 sg13g2_buf_1 fanout1305 (.A(net1318),
    .X(net1305));
 sg13g2_buf_4 fanout1306 (.X(net1306),
    .A(net1308));
 sg13g2_buf_4 fanout1307 (.X(net1307),
    .A(net1308));
 sg13g2_buf_2 fanout1308 (.A(net1318),
    .X(net1308));
 sg13g2_buf_4 fanout1309 (.X(net1309),
    .A(net1313));
 sg13g2_buf_2 fanout1310 (.A(net1313),
    .X(net1310));
 sg13g2_buf_4 fanout1311 (.X(net1311),
    .A(net1313));
 sg13g2_buf_2 fanout1312 (.A(net1313),
    .X(net1312));
 sg13g2_buf_1 fanout1313 (.A(net1318),
    .X(net1313));
 sg13g2_buf_4 fanout1314 (.X(net1314),
    .A(net1317));
 sg13g2_buf_4 fanout1315 (.X(net1315),
    .A(net1317));
 sg13g2_buf_4 fanout1316 (.X(net1316),
    .A(net1317));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_1 fanout1318 (.A(net1393),
    .X(net1318));
 sg13g2_buf_4 fanout1319 (.X(net1319),
    .A(net1322));
 sg13g2_buf_2 fanout1320 (.A(net1322),
    .X(net1320));
 sg13g2_buf_4 fanout1321 (.X(net1321),
    .A(net1322));
 sg13g2_buf_1 fanout1322 (.A(net1333),
    .X(net1322));
 sg13g2_buf_4 fanout1323 (.X(net1323),
    .A(net1325));
 sg13g2_buf_4 fanout1324 (.X(net1324),
    .A(net1325));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1333));
 sg13g2_buf_4 fanout1326 (.X(net1326),
    .A(net1328));
 sg13g2_buf_4 fanout1327 (.X(net1327),
    .A(net1328));
 sg13g2_buf_2 fanout1328 (.A(net1333),
    .X(net1328));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(net1332));
 sg13g2_buf_4 fanout1330 (.X(net1330),
    .A(net1331));
 sg13g2_buf_4 fanout1331 (.X(net1331),
    .A(net1332));
 sg13g2_buf_2 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_buf_1 fanout1333 (.A(net1393),
    .X(net1333));
 sg13g2_buf_4 fanout1334 (.X(net1334),
    .A(net1335));
 sg13g2_buf_4 fanout1335 (.X(net1335),
    .A(net1344));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(net1338));
 sg13g2_buf_4 fanout1337 (.X(net1337),
    .A(net1338));
 sg13g2_buf_2 fanout1338 (.A(net1344),
    .X(net1338));
 sg13g2_buf_4 fanout1339 (.X(net1339),
    .A(net1344));
 sg13g2_buf_2 fanout1340 (.A(net1344),
    .X(net1340));
 sg13g2_buf_4 fanout1341 (.X(net1341),
    .A(net1343));
 sg13g2_buf_4 fanout1342 (.X(net1342),
    .A(net1343));
 sg13g2_buf_4 fanout1343 (.X(net1343),
    .A(net1344));
 sg13g2_buf_1 fanout1344 (.A(net1392),
    .X(net1344));
 sg13g2_buf_4 fanout1345 (.X(net1345),
    .A(net1348));
 sg13g2_buf_2 fanout1346 (.A(net1348),
    .X(net1346));
 sg13g2_buf_4 fanout1347 (.X(net1347),
    .A(net1348));
 sg13g2_buf_1 fanout1348 (.A(net1362),
    .X(net1348));
 sg13g2_buf_4 fanout1349 (.X(net1349),
    .A(net1352));
 sg13g2_buf_2 fanout1350 (.A(net1352),
    .X(net1350));
 sg13g2_buf_4 fanout1351 (.X(net1351),
    .A(net1352));
 sg13g2_buf_2 fanout1352 (.A(net1362),
    .X(net1352));
 sg13g2_buf_4 fanout1353 (.X(net1353),
    .A(net1356));
 sg13g2_buf_4 fanout1354 (.X(net1354),
    .A(net1356));
 sg13g2_buf_2 fanout1355 (.A(net1356),
    .X(net1355));
 sg13g2_buf_1 fanout1356 (.A(net1362),
    .X(net1356));
 sg13g2_buf_4 fanout1357 (.X(net1357),
    .A(net1361));
 sg13g2_buf_2 fanout1358 (.A(net1361),
    .X(net1358));
 sg13g2_buf_4 fanout1359 (.X(net1359),
    .A(net1361));
 sg13g2_buf_2 fanout1360 (.A(net1361),
    .X(net1360));
 sg13g2_buf_1 fanout1361 (.A(net1362),
    .X(net1361));
 sg13g2_buf_1 fanout1362 (.A(net1392),
    .X(net1362));
 sg13g2_buf_4 fanout1363 (.X(net1363),
    .A(net1365));
 sg13g2_buf_4 fanout1364 (.X(net1364),
    .A(net1365));
 sg13g2_buf_4 fanout1365 (.X(net1365),
    .A(net1377));
 sg13g2_buf_4 fanout1366 (.X(net1366),
    .A(net1369));
 sg13g2_buf_4 fanout1367 (.X(net1367),
    .A(net1369));
 sg13g2_buf_2 fanout1368 (.A(net1369),
    .X(net1368));
 sg13g2_buf_2 fanout1369 (.A(net1377),
    .X(net1369));
 sg13g2_buf_4 fanout1370 (.X(net1370),
    .A(net1372));
 sg13g2_buf_4 fanout1371 (.X(net1371),
    .A(net1372));
 sg13g2_buf_2 fanout1372 (.A(net1377),
    .X(net1372));
 sg13g2_buf_4 fanout1373 (.X(net1373),
    .A(net1376));
 sg13g2_buf_4 fanout1374 (.X(net1374),
    .A(net1376));
 sg13g2_buf_2 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_2 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_1 fanout1377 (.A(net1392),
    .X(net1377));
 sg13g2_buf_4 fanout1378 (.X(net1378),
    .A(net1380));
 sg13g2_buf_4 fanout1379 (.X(net1379),
    .A(net1380));
 sg13g2_buf_2 fanout1380 (.A(net1391),
    .X(net1380));
 sg13g2_buf_4 fanout1381 (.X(net1381),
    .A(net1385));
 sg13g2_buf_2 fanout1382 (.A(net1385),
    .X(net1382));
 sg13g2_buf_4 fanout1383 (.X(net1383),
    .A(net1385));
 sg13g2_buf_2 fanout1384 (.A(net1385),
    .X(net1384));
 sg13g2_buf_1 fanout1385 (.A(net1391),
    .X(net1385));
 sg13g2_buf_4 fanout1386 (.X(net1386),
    .A(net1388));
 sg13g2_buf_4 fanout1387 (.X(net1387),
    .A(net1388));
 sg13g2_buf_4 fanout1388 (.X(net1388),
    .A(net1391));
 sg13g2_buf_4 fanout1389 (.X(net1389),
    .A(net1390));
 sg13g2_buf_4 fanout1390 (.X(net1390),
    .A(net1391));
 sg13g2_buf_2 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_1 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_1 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_1 fanout1394 (.A(net1),
    .X(net1394));
 sg13g2_tiehi _23936__1395 (.L_HI(net1395));
 sg13g2_tiehi _23937__1396 (.L_HI(net1396));
 sg13g2_tiehi _23938__1397 (.L_HI(net1397));
 sg13g2_tiehi _23939__1398 (.L_HI(net1398));
 sg13g2_tiehi _23940__1399 (.L_HI(net1399));
 sg13g2_tiehi _23941__1400 (.L_HI(net1400));
 sg13g2_tiehi _23942__1401 (.L_HI(net1401));
 sg13g2_tiehi _23943__1402 (.L_HI(net1402));
 sg13g2_tiehi \top_ihp.oisc.mem_addr_lowbits[0]$_DFF_P__1403  (.L_HI(net1403));
 sg13g2_tiehi \top_ihp.oisc.mem_addr_lowbits[1]$_DFF_P__1404  (.L_HI(net1404));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[0]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[1]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[2]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[3]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[4]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[5]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[6]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[7]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \top_ihp.oisc.regs[16][0]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \top_ihp.oisc.regs[16][10]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \top_ihp.oisc.regs[16][11]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \top_ihp.oisc.regs[16][12]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \top_ihp.oisc.regs[16][13]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \top_ihp.oisc.regs[16][14]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \top_ihp.oisc.regs[16][15]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \top_ihp.oisc.regs[16][16]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \top_ihp.oisc.regs[16][17]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \top_ihp.oisc.regs[16][18]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \top_ihp.oisc.regs[16][19]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \top_ihp.oisc.regs[16][1]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \top_ihp.oisc.regs[16][20]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \top_ihp.oisc.regs[16][21]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \top_ihp.oisc.regs[16][22]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \top_ihp.oisc.regs[16][23]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \top_ihp.oisc.regs[16][24]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \top_ihp.oisc.regs[16][25]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \top_ihp.oisc.regs[16][26]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \top_ihp.oisc.regs[16][27]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \top_ihp.oisc.regs[16][28]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \top_ihp.oisc.regs[16][29]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \top_ihp.oisc.regs[16][2]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \top_ihp.oisc.regs[16][30]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \top_ihp.oisc.regs[16][31]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \top_ihp.oisc.regs[16][3]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \top_ihp.oisc.regs[16][4]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \top_ihp.oisc.regs[16][5]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \top_ihp.oisc.regs[16][6]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \top_ihp.oisc.regs[16][7]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \top_ihp.oisc.regs[16][8]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \top_ihp.oisc.regs[16][9]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \top_ihp.oisc.regs[17][0]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \top_ihp.oisc.regs[17][10]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \top_ihp.oisc.regs[17][11]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \top_ihp.oisc.regs[17][12]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \top_ihp.oisc.regs[17][13]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \top_ihp.oisc.regs[17][14]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \top_ihp.oisc.regs[17][15]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \top_ihp.oisc.regs[17][16]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \top_ihp.oisc.regs[17][17]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \top_ihp.oisc.regs[17][18]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \top_ihp.oisc.regs[17][19]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \top_ihp.oisc.regs[17][1]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \top_ihp.oisc.regs[17][20]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \top_ihp.oisc.regs[17][21]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \top_ihp.oisc.regs[17][22]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \top_ihp.oisc.regs[17][23]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \top_ihp.oisc.regs[17][24]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \top_ihp.oisc.regs[17][25]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \top_ihp.oisc.regs[17][26]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \top_ihp.oisc.regs[17][27]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \top_ihp.oisc.regs[17][28]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \top_ihp.oisc.regs[17][29]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \top_ihp.oisc.regs[17][2]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \top_ihp.oisc.regs[17][30]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \top_ihp.oisc.regs[17][31]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \top_ihp.oisc.regs[17][3]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \top_ihp.oisc.regs[17][4]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \top_ihp.oisc.regs[17][5]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \top_ihp.oisc.regs[17][6]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \top_ihp.oisc.regs[17][7]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \top_ihp.oisc.regs[17][8]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \top_ihp.oisc.regs[17][9]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \top_ihp.oisc.regs[18][0]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \top_ihp.oisc.regs[18][10]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \top_ihp.oisc.regs[18][11]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \top_ihp.oisc.regs[18][12]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \top_ihp.oisc.regs[18][13]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \top_ihp.oisc.regs[18][14]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \top_ihp.oisc.regs[18][15]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \top_ihp.oisc.regs[18][16]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \top_ihp.oisc.regs[18][17]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \top_ihp.oisc.regs[18][18]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \top_ihp.oisc.regs[18][19]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \top_ihp.oisc.regs[18][1]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \top_ihp.oisc.regs[18][20]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \top_ihp.oisc.regs[18][21]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \top_ihp.oisc.regs[18][22]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \top_ihp.oisc.regs[18][23]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \top_ihp.oisc.regs[18][24]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \top_ihp.oisc.regs[18][25]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \top_ihp.oisc.regs[18][26]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \top_ihp.oisc.regs[18][27]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \top_ihp.oisc.regs[18][28]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \top_ihp.oisc.regs[18][29]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \top_ihp.oisc.regs[18][2]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \top_ihp.oisc.regs[18][30]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \top_ihp.oisc.regs[18][31]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \top_ihp.oisc.regs[18][3]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \top_ihp.oisc.regs[18][4]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \top_ihp.oisc.regs[18][5]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \top_ihp.oisc.regs[18][6]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \top_ihp.oisc.regs[18][7]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \top_ihp.oisc.regs[18][8]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \top_ihp.oisc.regs[18][9]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \top_ihp.oisc.regs[19][0]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \top_ihp.oisc.regs[19][10]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \top_ihp.oisc.regs[19][11]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \top_ihp.oisc.regs[19][12]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \top_ihp.oisc.regs[19][13]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \top_ihp.oisc.regs[19][14]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \top_ihp.oisc.regs[19][15]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \top_ihp.oisc.regs[19][16]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \top_ihp.oisc.regs[19][17]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \top_ihp.oisc.regs[19][18]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \top_ihp.oisc.regs[19][19]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \top_ihp.oisc.regs[19][1]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \top_ihp.oisc.regs[19][20]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \top_ihp.oisc.regs[19][21]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \top_ihp.oisc.regs[19][22]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \top_ihp.oisc.regs[19][23]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \top_ihp.oisc.regs[19][24]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \top_ihp.oisc.regs[19][25]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \top_ihp.oisc.regs[19][26]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \top_ihp.oisc.regs[19][27]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \top_ihp.oisc.regs[19][28]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \top_ihp.oisc.regs[19][29]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \top_ihp.oisc.regs[19][2]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \top_ihp.oisc.regs[19][30]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \top_ihp.oisc.regs[19][31]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \top_ihp.oisc.regs[19][3]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \top_ihp.oisc.regs[19][4]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \top_ihp.oisc.regs[19][5]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \top_ihp.oisc.regs[19][6]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \top_ihp.oisc.regs[19][7]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \top_ihp.oisc.regs[19][8]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \top_ihp.oisc.regs[19][9]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \top_ihp.oisc.regs[20][0]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \top_ihp.oisc.regs[20][10]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \top_ihp.oisc.regs[20][11]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \top_ihp.oisc.regs[20][12]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \top_ihp.oisc.regs[20][13]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \top_ihp.oisc.regs[20][14]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \top_ihp.oisc.regs[20][15]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \top_ihp.oisc.regs[20][16]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \top_ihp.oisc.regs[20][17]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \top_ihp.oisc.regs[20][18]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \top_ihp.oisc.regs[20][19]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \top_ihp.oisc.regs[20][1]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \top_ihp.oisc.regs[20][20]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \top_ihp.oisc.regs[20][21]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \top_ihp.oisc.regs[20][22]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \top_ihp.oisc.regs[20][23]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \top_ihp.oisc.regs[20][24]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \top_ihp.oisc.regs[20][25]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \top_ihp.oisc.regs[20][26]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \top_ihp.oisc.regs[20][27]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \top_ihp.oisc.regs[20][28]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \top_ihp.oisc.regs[20][29]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \top_ihp.oisc.regs[20][2]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \top_ihp.oisc.regs[20][30]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \top_ihp.oisc.regs[20][31]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \top_ihp.oisc.regs[20][3]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \top_ihp.oisc.regs[20][4]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \top_ihp.oisc.regs[20][5]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \top_ihp.oisc.regs[20][6]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \top_ihp.oisc.regs[20][7]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \top_ihp.oisc.regs[20][8]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \top_ihp.oisc.regs[20][9]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \top_ihp.oisc.regs[21][0]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \top_ihp.oisc.regs[21][10]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \top_ihp.oisc.regs[21][11]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \top_ihp.oisc.regs[21][12]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \top_ihp.oisc.regs[21][13]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \top_ihp.oisc.regs[21][14]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \top_ihp.oisc.regs[21][15]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \top_ihp.oisc.regs[21][16]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \top_ihp.oisc.regs[21][17]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \top_ihp.oisc.regs[21][18]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \top_ihp.oisc.regs[21][19]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \top_ihp.oisc.regs[21][1]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \top_ihp.oisc.regs[21][20]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \top_ihp.oisc.regs[21][21]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \top_ihp.oisc.regs[21][22]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \top_ihp.oisc.regs[21][23]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \top_ihp.oisc.regs[21][24]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \top_ihp.oisc.regs[21][25]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \top_ihp.oisc.regs[21][26]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \top_ihp.oisc.regs[21][27]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \top_ihp.oisc.regs[21][28]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \top_ihp.oisc.regs[21][29]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \top_ihp.oisc.regs[21][2]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \top_ihp.oisc.regs[21][30]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \top_ihp.oisc.regs[21][31]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \top_ihp.oisc.regs[21][3]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \top_ihp.oisc.regs[21][4]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \top_ihp.oisc.regs[21][5]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \top_ihp.oisc.regs[21][6]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \top_ihp.oisc.regs[21][7]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \top_ihp.oisc.regs[21][8]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \top_ihp.oisc.regs[21][9]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \top_ihp.oisc.regs[22][0]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \top_ihp.oisc.regs[22][10]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \top_ihp.oisc.regs[22][11]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \top_ihp.oisc.regs[22][12]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \top_ihp.oisc.regs[22][13]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \top_ihp.oisc.regs[22][14]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \top_ihp.oisc.regs[22][15]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \top_ihp.oisc.regs[22][16]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \top_ihp.oisc.regs[22][17]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \top_ihp.oisc.regs[22][18]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \top_ihp.oisc.regs[22][19]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \top_ihp.oisc.regs[22][1]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \top_ihp.oisc.regs[22][20]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \top_ihp.oisc.regs[22][21]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \top_ihp.oisc.regs[22][22]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \top_ihp.oisc.regs[22][23]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \top_ihp.oisc.regs[22][24]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \top_ihp.oisc.regs[22][25]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \top_ihp.oisc.regs[22][26]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \top_ihp.oisc.regs[22][27]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \top_ihp.oisc.regs[22][28]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \top_ihp.oisc.regs[22][29]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \top_ihp.oisc.regs[22][2]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \top_ihp.oisc.regs[22][30]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \top_ihp.oisc.regs[22][31]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \top_ihp.oisc.regs[22][3]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \top_ihp.oisc.regs[22][4]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \top_ihp.oisc.regs[22][5]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \top_ihp.oisc.regs[22][6]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \top_ihp.oisc.regs[22][7]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \top_ihp.oisc.regs[22][8]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \top_ihp.oisc.regs[22][9]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \top_ihp.oisc.regs[23][0]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \top_ihp.oisc.regs[23][10]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \top_ihp.oisc.regs[23][11]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \top_ihp.oisc.regs[23][12]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \top_ihp.oisc.regs[23][13]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \top_ihp.oisc.regs[23][14]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \top_ihp.oisc.regs[23][15]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \top_ihp.oisc.regs[23][16]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \top_ihp.oisc.regs[23][17]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \top_ihp.oisc.regs[23][18]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \top_ihp.oisc.regs[23][19]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \top_ihp.oisc.regs[23][1]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \top_ihp.oisc.regs[23][20]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \top_ihp.oisc.regs[23][21]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \top_ihp.oisc.regs[23][22]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \top_ihp.oisc.regs[23][23]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \top_ihp.oisc.regs[23][24]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \top_ihp.oisc.regs[23][25]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \top_ihp.oisc.regs[23][26]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \top_ihp.oisc.regs[23][27]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \top_ihp.oisc.regs[23][28]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \top_ihp.oisc.regs[23][29]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \top_ihp.oisc.regs[23][2]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \top_ihp.oisc.regs[23][30]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \top_ihp.oisc.regs[23][31]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \top_ihp.oisc.regs[23][3]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \top_ihp.oisc.regs[23][4]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \top_ihp.oisc.regs[23][5]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \top_ihp.oisc.regs[23][6]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \top_ihp.oisc.regs[23][7]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \top_ihp.oisc.regs[23][8]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \top_ihp.oisc.regs[23][9]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \top_ihp.oisc.regs[24][0]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \top_ihp.oisc.regs[24][10]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \top_ihp.oisc.regs[24][11]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \top_ihp.oisc.regs[24][12]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \top_ihp.oisc.regs[24][13]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \top_ihp.oisc.regs[24][14]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \top_ihp.oisc.regs[24][15]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \top_ihp.oisc.regs[24][16]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \top_ihp.oisc.regs[24][17]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \top_ihp.oisc.regs[24][18]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \top_ihp.oisc.regs[24][19]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \top_ihp.oisc.regs[24][1]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \top_ihp.oisc.regs[24][20]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \top_ihp.oisc.regs[24][21]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \top_ihp.oisc.regs[24][22]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \top_ihp.oisc.regs[24][23]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \top_ihp.oisc.regs[24][24]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \top_ihp.oisc.regs[24][25]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \top_ihp.oisc.regs[24][26]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \top_ihp.oisc.regs[24][27]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \top_ihp.oisc.regs[24][28]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \top_ihp.oisc.regs[24][29]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \top_ihp.oisc.regs[24][2]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \top_ihp.oisc.regs[24][30]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \top_ihp.oisc.regs[24][31]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \top_ihp.oisc.regs[24][3]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \top_ihp.oisc.regs[24][4]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \top_ihp.oisc.regs[24][5]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \top_ihp.oisc.regs[24][6]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \top_ihp.oisc.regs[24][7]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \top_ihp.oisc.regs[24][8]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \top_ihp.oisc.regs[24][9]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \top_ihp.oisc.regs[25][0]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \top_ihp.oisc.regs[25][10]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \top_ihp.oisc.regs[25][11]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \top_ihp.oisc.regs[25][12]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \top_ihp.oisc.regs[25][13]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \top_ihp.oisc.regs[25][14]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \top_ihp.oisc.regs[25][15]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \top_ihp.oisc.regs[25][16]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \top_ihp.oisc.regs[25][17]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \top_ihp.oisc.regs[25][18]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \top_ihp.oisc.regs[25][19]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \top_ihp.oisc.regs[25][1]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \top_ihp.oisc.regs[25][20]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \top_ihp.oisc.regs[25][21]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \top_ihp.oisc.regs[25][22]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \top_ihp.oisc.regs[25][23]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \top_ihp.oisc.regs[25][24]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \top_ihp.oisc.regs[25][25]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \top_ihp.oisc.regs[25][26]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \top_ihp.oisc.regs[25][27]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \top_ihp.oisc.regs[25][28]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \top_ihp.oisc.regs[25][29]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \top_ihp.oisc.regs[25][2]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \top_ihp.oisc.regs[25][30]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \top_ihp.oisc.regs[25][31]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \top_ihp.oisc.regs[25][3]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \top_ihp.oisc.regs[25][4]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \top_ihp.oisc.regs[25][5]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \top_ihp.oisc.regs[25][6]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \top_ihp.oisc.regs[25][7]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \top_ihp.oisc.regs[25][8]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \top_ihp.oisc.regs[25][9]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \top_ihp.oisc.regs[26][0]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \top_ihp.oisc.regs[26][10]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \top_ihp.oisc.regs[26][11]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \top_ihp.oisc.regs[26][12]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \top_ihp.oisc.regs[26][13]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \top_ihp.oisc.regs[26][14]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \top_ihp.oisc.regs[26][15]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \top_ihp.oisc.regs[26][16]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \top_ihp.oisc.regs[26][17]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \top_ihp.oisc.regs[26][18]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \top_ihp.oisc.regs[26][19]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \top_ihp.oisc.regs[26][1]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \top_ihp.oisc.regs[26][20]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \top_ihp.oisc.regs[26][21]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \top_ihp.oisc.regs[26][22]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \top_ihp.oisc.regs[26][23]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \top_ihp.oisc.regs[26][24]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \top_ihp.oisc.regs[26][25]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \top_ihp.oisc.regs[26][26]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \top_ihp.oisc.regs[26][27]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \top_ihp.oisc.regs[26][28]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \top_ihp.oisc.regs[26][29]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \top_ihp.oisc.regs[26][2]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \top_ihp.oisc.regs[26][30]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \top_ihp.oisc.regs[26][31]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \top_ihp.oisc.regs[26][3]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \top_ihp.oisc.regs[26][4]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \top_ihp.oisc.regs[26][5]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \top_ihp.oisc.regs[26][6]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \top_ihp.oisc.regs[26][7]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \top_ihp.oisc.regs[26][8]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \top_ihp.oisc.regs[26][9]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \top_ihp.oisc.regs[27][0]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \top_ihp.oisc.regs[27][10]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \top_ihp.oisc.regs[27][11]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \top_ihp.oisc.regs[27][12]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \top_ihp.oisc.regs[27][13]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \top_ihp.oisc.regs[27][14]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \top_ihp.oisc.regs[27][15]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \top_ihp.oisc.regs[27][16]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \top_ihp.oisc.regs[27][17]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \top_ihp.oisc.regs[27][18]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \top_ihp.oisc.regs[27][19]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \top_ihp.oisc.regs[27][1]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \top_ihp.oisc.regs[27][20]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \top_ihp.oisc.regs[27][21]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \top_ihp.oisc.regs[27][22]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \top_ihp.oisc.regs[27][23]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \top_ihp.oisc.regs[27][24]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \top_ihp.oisc.regs[27][25]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \top_ihp.oisc.regs[27][26]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \top_ihp.oisc.regs[27][27]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \top_ihp.oisc.regs[27][28]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \top_ihp.oisc.regs[27][29]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \top_ihp.oisc.regs[27][2]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \top_ihp.oisc.regs[27][30]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \top_ihp.oisc.regs[27][31]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \top_ihp.oisc.regs[27][3]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \top_ihp.oisc.regs[27][4]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \top_ihp.oisc.regs[27][5]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \top_ihp.oisc.regs[27][6]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \top_ihp.oisc.regs[27][7]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \top_ihp.oisc.regs[27][8]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \top_ihp.oisc.regs[27][9]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \top_ihp.oisc.regs[28][0]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \top_ihp.oisc.regs[28][10]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \top_ihp.oisc.regs[28][11]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \top_ihp.oisc.regs[28][12]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \top_ihp.oisc.regs[28][13]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \top_ihp.oisc.regs[28][14]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \top_ihp.oisc.regs[28][15]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \top_ihp.oisc.regs[28][16]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \top_ihp.oisc.regs[28][17]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \top_ihp.oisc.regs[28][18]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \top_ihp.oisc.regs[28][19]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \top_ihp.oisc.regs[28][1]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \top_ihp.oisc.regs[28][20]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \top_ihp.oisc.regs[28][21]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \top_ihp.oisc.regs[28][22]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \top_ihp.oisc.regs[28][23]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \top_ihp.oisc.regs[28][24]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \top_ihp.oisc.regs[28][25]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \top_ihp.oisc.regs[28][26]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \top_ihp.oisc.regs[28][27]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \top_ihp.oisc.regs[28][28]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \top_ihp.oisc.regs[28][29]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \top_ihp.oisc.regs[28][2]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \top_ihp.oisc.regs[28][30]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \top_ihp.oisc.regs[28][31]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \top_ihp.oisc.regs[28][3]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \top_ihp.oisc.regs[28][4]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \top_ihp.oisc.regs[28][5]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \top_ihp.oisc.regs[28][6]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \top_ihp.oisc.regs[28][7]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \top_ihp.oisc.regs[28][8]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \top_ihp.oisc.regs[28][9]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \top_ihp.oisc.regs[29][0]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \top_ihp.oisc.regs[29][10]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \top_ihp.oisc.regs[29][11]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \top_ihp.oisc.regs[29][12]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \top_ihp.oisc.regs[29][13]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \top_ihp.oisc.regs[29][14]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \top_ihp.oisc.regs[29][15]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \top_ihp.oisc.regs[29][16]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \top_ihp.oisc.regs[29][17]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \top_ihp.oisc.regs[29][18]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \top_ihp.oisc.regs[29][19]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \top_ihp.oisc.regs[29][1]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \top_ihp.oisc.regs[29][20]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \top_ihp.oisc.regs[29][21]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \top_ihp.oisc.regs[29][22]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \top_ihp.oisc.regs[29][23]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \top_ihp.oisc.regs[29][24]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \top_ihp.oisc.regs[29][25]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \top_ihp.oisc.regs[29][26]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \top_ihp.oisc.regs[29][27]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \top_ihp.oisc.regs[29][28]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \top_ihp.oisc.regs[29][29]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \top_ihp.oisc.regs[29][2]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \top_ihp.oisc.regs[29][30]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \top_ihp.oisc.regs[29][31]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \top_ihp.oisc.regs[29][3]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \top_ihp.oisc.regs[29][4]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \top_ihp.oisc.regs[29][5]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \top_ihp.oisc.regs[29][6]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \top_ihp.oisc.regs[29][7]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \top_ihp.oisc.regs[29][8]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \top_ihp.oisc.regs[29][9]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \top_ihp.oisc.regs[30][0]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \top_ihp.oisc.regs[30][10]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \top_ihp.oisc.regs[30][11]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \top_ihp.oisc.regs[30][12]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \top_ihp.oisc.regs[30][13]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \top_ihp.oisc.regs[30][14]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \top_ihp.oisc.regs[30][15]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \top_ihp.oisc.regs[30][16]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \top_ihp.oisc.regs[30][17]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \top_ihp.oisc.regs[30][18]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \top_ihp.oisc.regs[30][19]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \top_ihp.oisc.regs[30][1]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \top_ihp.oisc.regs[30][20]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \top_ihp.oisc.regs[30][21]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \top_ihp.oisc.regs[30][22]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \top_ihp.oisc.regs[30][23]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \top_ihp.oisc.regs[30][24]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \top_ihp.oisc.regs[30][25]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \top_ihp.oisc.regs[30][26]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \top_ihp.oisc.regs[30][27]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \top_ihp.oisc.regs[30][28]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \top_ihp.oisc.regs[30][29]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \top_ihp.oisc.regs[30][2]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \top_ihp.oisc.regs[30][30]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \top_ihp.oisc.regs[30][31]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \top_ihp.oisc.regs[30][3]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \top_ihp.oisc.regs[30][4]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \top_ihp.oisc.regs[30][5]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \top_ihp.oisc.regs[30][6]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \top_ihp.oisc.regs[30][7]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \top_ihp.oisc.regs[30][8]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \top_ihp.oisc.regs[30][9]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \top_ihp.oisc.regs[31][0]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \top_ihp.oisc.regs[31][10]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \top_ihp.oisc.regs[31][11]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \top_ihp.oisc.regs[31][12]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \top_ihp.oisc.regs[31][13]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \top_ihp.oisc.regs[31][14]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \top_ihp.oisc.regs[31][15]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \top_ihp.oisc.regs[31][16]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \top_ihp.oisc.regs[31][17]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \top_ihp.oisc.regs[31][18]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \top_ihp.oisc.regs[31][19]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \top_ihp.oisc.regs[31][1]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \top_ihp.oisc.regs[31][20]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \top_ihp.oisc.regs[31][21]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \top_ihp.oisc.regs[31][22]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \top_ihp.oisc.regs[31][23]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \top_ihp.oisc.regs[31][24]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \top_ihp.oisc.regs[31][25]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \top_ihp.oisc.regs[31][26]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \top_ihp.oisc.regs[31][27]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \top_ihp.oisc.regs[31][28]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \top_ihp.oisc.regs[31][29]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \top_ihp.oisc.regs[31][2]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \top_ihp.oisc.regs[31][30]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \top_ihp.oisc.regs[31][31]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \top_ihp.oisc.regs[31][3]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \top_ihp.oisc.regs[31][4]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \top_ihp.oisc.regs[31][5]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \top_ihp.oisc.regs[31][6]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \top_ihp.oisc.regs[31][7]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \top_ihp.oisc.regs[31][8]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \top_ihp.oisc.regs[31][9]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \top_ihp.oisc.regs[32][0]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \top_ihp.oisc.regs[32][10]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \top_ihp.oisc.regs[32][11]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \top_ihp.oisc.regs[32][12]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \top_ihp.oisc.regs[32][13]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \top_ihp.oisc.regs[32][14]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \top_ihp.oisc.regs[32][15]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \top_ihp.oisc.regs[32][16]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \top_ihp.oisc.regs[32][17]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \top_ihp.oisc.regs[32][18]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \top_ihp.oisc.regs[32][19]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \top_ihp.oisc.regs[32][1]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \top_ihp.oisc.regs[32][20]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \top_ihp.oisc.regs[32][21]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \top_ihp.oisc.regs[32][22]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \top_ihp.oisc.regs[32][23]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \top_ihp.oisc.regs[32][24]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \top_ihp.oisc.regs[32][25]$_DFFE_PP__1942  (.L_HI(net1942));
 sg13g2_tiehi \top_ihp.oisc.regs[32][26]$_DFFE_PP__1943  (.L_HI(net1943));
 sg13g2_tiehi \top_ihp.oisc.regs[32][27]$_DFFE_PP__1944  (.L_HI(net1944));
 sg13g2_tiehi \top_ihp.oisc.regs[32][28]$_DFFE_PP__1945  (.L_HI(net1945));
 sg13g2_tiehi \top_ihp.oisc.regs[32][29]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \top_ihp.oisc.regs[32][2]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \top_ihp.oisc.regs[32][30]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \top_ihp.oisc.regs[32][31]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \top_ihp.oisc.regs[32][3]$_DFFE_PP__1950  (.L_HI(net1950));
 sg13g2_tiehi \top_ihp.oisc.regs[32][4]$_DFFE_PP__1951  (.L_HI(net1951));
 sg13g2_tiehi \top_ihp.oisc.regs[32][5]$_DFFE_PP__1952  (.L_HI(net1952));
 sg13g2_tiehi \top_ihp.oisc.regs[32][6]$_DFFE_PP__1953  (.L_HI(net1953));
 sg13g2_tiehi \top_ihp.oisc.regs[32][7]$_DFFE_PP__1954  (.L_HI(net1954));
 sg13g2_tiehi \top_ihp.oisc.regs[32][8]$_DFFE_PP__1955  (.L_HI(net1955));
 sg13g2_tiehi \top_ihp.oisc.regs[32][9]$_DFFE_PP__1956  (.L_HI(net1956));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[0]$_SDFFCE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[1]$_SDFFCE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[2]$_SDFFCE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[3]$_SDFFCE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[4]$_SDFFCE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[5]$_SDFFCE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[6]$_SDFFCE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[7]$_SDFFCE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \top_ihp.wb_emem.last_bit$_DFFE_PP__1965  (.L_HI(net1965));
 sg13g2_tiehi \top_ihp.wb_emem.last_wait$_DFFE_PP__1966  (.L_HI(net1966));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[3]$_SDFFCE_NP1P__1967  (.L_HI(net1967));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[4]$_SDFFCE_NP0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[5]$_SDFFCE_NP0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[6]$_SDFFCE_NP0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[0]$_SDFFCE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[1]$_SDFFCE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[2]$_SDFFCE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[3]$_SDFFCE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[4]$_SDFFCE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[5]$_SDFFCE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[6]$_SDFFCE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[7]$_SDFFCE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \top_ihp.wb_uart.ack_o$_SDFFCE_PP0P__1979  (.L_HI(net1979));
 sg13g2_inv_1 net1791_2 (.Y(net1981),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 net1791_3 (.Y(net1982),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net1791_4 (.Y(net1983),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_5 (.Y(net1984),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 net1791_6 (.Y(net1985),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net1791_7 (.Y(net1986),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_8 (.Y(net1987),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_9 (.Y(net1988),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_10 (.Y(net1989),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_11 (.Y(net1990),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 net1791_12 (.Y(net1991),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 net1791_13 (.Y(net1992),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 net1791_14 (.Y(net1993),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net1791_15 (.Y(net1994),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net1791_16 (.Y(net1995),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 net1791_17 (.Y(net1996),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net1791_18 (.Y(net1997),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net1791_19 (.Y(net1998),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net1791_20 (.Y(net1999),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net1791_21 (.Y(net2000),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_22 (.Y(net2001),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_23 (.Y(net2002),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_24 (.Y(net2003),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_25 (.Y(net2004),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net1791_26 (.Y(net2005),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_27 (.Y(net2006),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net1791_28 (.Y(net2007),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 net1791_29 (.Y(net2008),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 net1791_30 (.Y(net2009),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 net1791_31 (.Y(net2010),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 net1791_32 (.Y(net2011),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 net1791_33 (.Y(net2012),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 net1791_34 (.Y(net2013),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _35 (.Y(net2014),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _35_36 (.Y(net2015),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _35_37 (.Y(net2016),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _35_38 (.Y(net2017),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _35_39 (.Y(net2018),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _35_40 (.Y(net2019),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _35_41 (.Y(net2020),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _35_42 (.Y(net2021),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _35_43 (.Y(net2022),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _35_44 (.Y(net2023),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _35_45 (.Y(net2024),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _35_46 (.Y(net2025),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_47 (.Y(net2026),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _35_48 (.Y(net2027),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _35_49 (.Y(net2028),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_50 (.Y(net2029),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_51 (.Y(net2030),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _35_52 (.Y(net2031),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_53 (.Y(net2032),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_54 (.Y(net2033),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_55 (.Y(net2034),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_56 (.Y(net2035),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_57 (.Y(net2036),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _35_58 (.Y(net2037),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _35_59 (.Y(net2038),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _35_60 (.Y(net2039),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _35_61 (.Y(net2040),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_62 (.Y(net2041),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _35_63 (.Y(net2042),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _35_64 (.Y(net2043),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _35_65 (.Y(net2044),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_66 (.Y(net2045),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _35_67 (.Y(net2046),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _35_68 (.Y(net2047),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _35_69 (.Y(net2048),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _35_70 (.Y(net2049),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _35_71 (.Y(net2050),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _35_72 (.Y(net2051),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_73 (.Y(net2052),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _35_74 (.Y(net2053),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _35_75 (.Y(net2054),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _35_76 (.Y(net2055),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _35_77 (.Y(net2056),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _35_78 (.Y(net2057),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _35_79 (.Y(net2058),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _35_80 (.Y(net2059),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _35_81 (.Y(net2060),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _35_82 (.Y(net2061),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_83 (.Y(net2062),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _35_84 (.Y(net2063),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _35_85 (.Y(net2064),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _35_86 (.Y(net2065),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_87 (.Y(net2066),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_88 (.Y(net2067),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _35_89 (.Y(net2068),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_90 (.Y(net2069),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_91 (.Y(net2070),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_92 (.Y(net2071),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_93 (.Y(net2072),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_94 (.Y(net2073),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _35_95 (.Y(net2074),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _35_96 (.Y(net2075),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _35_97 (.Y(net2076),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _35_98 (.Y(net2077),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_99 (.Y(net2078),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_100 (.Y(net2079),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_101 (.Y(net2080),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_102 (.Y(net2081),
    .A(clknet_leaf_310_clk));
 sg13g2_inv_1 _35_103 (.Y(net2082),
    .A(clknet_leaf_310_clk));
 sg13g2_inv_1 _35_104 (.Y(net2083),
    .A(clknet_leaf_310_clk));
 sg13g2_inv_1 _35_105 (.Y(net2084),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _35_106 (.Y(net2085),
    .A(clknet_leaf_309_clk));
 sg13g2_inv_1 _35_107 (.Y(net2086),
    .A(clknet_leaf_309_clk));
 sg13g2_inv_1 _35_108 (.Y(net2087),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _35_109 (.Y(net2088),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _35_110 (.Y(net2089),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_111 (.Y(net2090),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_112 (.Y(net2091),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_113 (.Y(net2092),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _35_114 (.Y(net2093),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_115 (.Y(net2094),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _35_116 (.Y(net2095),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _35_117 (.Y(net2096),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _35_118 (.Y(net2097),
    .A(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_313_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_41_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00294_));
 sg13g2_antennanp ANTENNA_2 (.A(_00294_));
 sg13g2_antennanp ANTENNA_3 (.A(_00296_));
 sg13g2_antennanp ANTENNA_4 (.A(_00296_));
 sg13g2_antennanp ANTENNA_5 (.A(_00296_));
 sg13g2_antennanp ANTENNA_6 (.A(_00299_));
 sg13g2_antennanp ANTENNA_7 (.A(_00300_));
 sg13g2_antennanp ANTENNA_8 (.A(_00300_));
 sg13g2_antennanp ANTENNA_9 (.A(_00300_));
 sg13g2_antennanp ANTENNA_10 (.A(_00305_));
 sg13g2_antennanp ANTENNA_11 (.A(_00307_));
 sg13g2_antennanp ANTENNA_12 (.A(_00307_));
 sg13g2_antennanp ANTENNA_13 (.A(_00311_));
 sg13g2_antennanp ANTENNA_14 (.A(_00311_));
 sg13g2_antennanp ANTENNA_15 (.A(_00316_));
 sg13g2_antennanp ANTENNA_16 (.A(_00316_));
 sg13g2_antennanp ANTENNA_17 (.A(_00316_));
 sg13g2_antennanp ANTENNA_18 (.A(_00319_));
 sg13g2_antennanp ANTENNA_19 (.A(_00320_));
 sg13g2_antennanp ANTENNA_20 (.A(_00322_));
 sg13g2_antennanp ANTENNA_21 (.A(_00322_));
 sg13g2_antennanp ANTENNA_22 (.A(_00323_));
 sg13g2_antennanp ANTENNA_23 (.A(_00324_));
 sg13g2_antennanp ANTENNA_24 (.A(_02668_));
 sg13g2_antennanp ANTENNA_25 (.A(_02668_));
 sg13g2_antennanp ANTENNA_26 (.A(_02668_));
 sg13g2_antennanp ANTENNA_27 (.A(_02668_));
 sg13g2_antennanp ANTENNA_28 (.A(_02670_));
 sg13g2_antennanp ANTENNA_29 (.A(_02670_));
 sg13g2_antennanp ANTENNA_30 (.A(_02670_));
 sg13g2_antennanp ANTENNA_31 (.A(_02670_));
 sg13g2_antennanp ANTENNA_32 (.A(_02718_));
 sg13g2_antennanp ANTENNA_33 (.A(_02718_));
 sg13g2_antennanp ANTENNA_34 (.A(_02718_));
 sg13g2_antennanp ANTENNA_35 (.A(_02777_));
 sg13g2_antennanp ANTENNA_36 (.A(_02777_));
 sg13g2_antennanp ANTENNA_37 (.A(_02777_));
 sg13g2_antennanp ANTENNA_38 (.A(_02845_));
 sg13g2_antennanp ANTENNA_39 (.A(_02845_));
 sg13g2_antennanp ANTENNA_40 (.A(_02845_));
 sg13g2_antennanp ANTENNA_41 (.A(_02845_));
 sg13g2_antennanp ANTENNA_42 (.A(_02845_));
 sg13g2_antennanp ANTENNA_43 (.A(_02845_));
 sg13g2_antennanp ANTENNA_44 (.A(_02845_));
 sg13g2_antennanp ANTENNA_45 (.A(_03021_));
 sg13g2_antennanp ANTENNA_46 (.A(_03021_));
 sg13g2_antennanp ANTENNA_47 (.A(_03021_));
 sg13g2_antennanp ANTENNA_48 (.A(_03090_));
 sg13g2_antennanp ANTENNA_49 (.A(_03090_));
 sg13g2_antennanp ANTENNA_50 (.A(_03090_));
 sg13g2_antennanp ANTENNA_51 (.A(_03090_));
 sg13g2_antennanp ANTENNA_52 (.A(_03090_));
 sg13g2_antennanp ANTENNA_53 (.A(_03101_));
 sg13g2_antennanp ANTENNA_54 (.A(_03101_));
 sg13g2_antennanp ANTENNA_55 (.A(_03101_));
 sg13g2_antennanp ANTENNA_56 (.A(_03101_));
 sg13g2_antennanp ANTENNA_57 (.A(_03148_));
 sg13g2_antennanp ANTENNA_58 (.A(_03148_));
 sg13g2_antennanp ANTENNA_59 (.A(_03148_));
 sg13g2_antennanp ANTENNA_60 (.A(_03148_));
 sg13g2_antennanp ANTENNA_61 (.A(_03148_));
 sg13g2_antennanp ANTENNA_62 (.A(_03148_));
 sg13g2_antennanp ANTENNA_63 (.A(_03148_));
 sg13g2_antennanp ANTENNA_64 (.A(_03148_));
 sg13g2_antennanp ANTENNA_65 (.A(_03713_));
 sg13g2_antennanp ANTENNA_66 (.A(_04741_));
 sg13g2_antennanp ANTENNA_67 (.A(_04741_));
 sg13g2_antennanp ANTENNA_68 (.A(_04741_));
 sg13g2_antennanp ANTENNA_69 (.A(_04741_));
 sg13g2_antennanp ANTENNA_70 (.A(_04741_));
 sg13g2_antennanp ANTENNA_71 (.A(_04741_));
 sg13g2_antennanp ANTENNA_72 (.A(_04741_));
 sg13g2_antennanp ANTENNA_73 (.A(_04741_));
 sg13g2_antennanp ANTENNA_74 (.A(_04799_));
 sg13g2_antennanp ANTENNA_75 (.A(_04799_));
 sg13g2_antennanp ANTENNA_76 (.A(_04799_));
 sg13g2_antennanp ANTENNA_77 (.A(_04799_));
 sg13g2_antennanp ANTENNA_78 (.A(_04799_));
 sg13g2_antennanp ANTENNA_79 (.A(_04799_));
 sg13g2_antennanp ANTENNA_80 (.A(_04847_));
 sg13g2_antennanp ANTENNA_81 (.A(_04847_));
 sg13g2_antennanp ANTENNA_82 (.A(_04847_));
 sg13g2_antennanp ANTENNA_83 (.A(_04847_));
 sg13g2_antennanp ANTENNA_84 (.A(_04851_));
 sg13g2_antennanp ANTENNA_85 (.A(_04851_));
 sg13g2_antennanp ANTENNA_86 (.A(_04851_));
 sg13g2_antennanp ANTENNA_87 (.A(_04851_));
 sg13g2_antennanp ANTENNA_88 (.A(_04857_));
 sg13g2_antennanp ANTENNA_89 (.A(_04871_));
 sg13g2_antennanp ANTENNA_90 (.A(_04871_));
 sg13g2_antennanp ANTENNA_91 (.A(_04871_));
 sg13g2_antennanp ANTENNA_92 (.A(_04873_));
 sg13g2_antennanp ANTENNA_93 (.A(_04873_));
 sg13g2_antennanp ANTENNA_94 (.A(_04873_));
 sg13g2_antennanp ANTENNA_95 (.A(_04883_));
 sg13g2_antennanp ANTENNA_96 (.A(_04912_));
 sg13g2_antennanp ANTENNA_97 (.A(_04917_));
 sg13g2_antennanp ANTENNA_98 (.A(_04917_));
 sg13g2_antennanp ANTENNA_99 (.A(_04917_));
 sg13g2_antennanp ANTENNA_100 (.A(_04917_));
 sg13g2_antennanp ANTENNA_101 (.A(_04917_));
 sg13g2_antennanp ANTENNA_102 (.A(_04917_));
 sg13g2_antennanp ANTENNA_103 (.A(_04920_));
 sg13g2_antennanp ANTENNA_104 (.A(_04920_));
 sg13g2_antennanp ANTENNA_105 (.A(_04920_));
 sg13g2_antennanp ANTENNA_106 (.A(_04921_));
 sg13g2_antennanp ANTENNA_107 (.A(_04921_));
 sg13g2_antennanp ANTENNA_108 (.A(_04921_));
 sg13g2_antennanp ANTENNA_109 (.A(_04925_));
 sg13g2_antennanp ANTENNA_110 (.A(_04925_));
 sg13g2_antennanp ANTENNA_111 (.A(_04932_));
 sg13g2_antennanp ANTENNA_112 (.A(_05012_));
 sg13g2_antennanp ANTENNA_113 (.A(_05012_));
 sg13g2_antennanp ANTENNA_114 (.A(_05012_));
 sg13g2_antennanp ANTENNA_115 (.A(_05012_));
 sg13g2_antennanp ANTENNA_116 (.A(_05012_));
 sg13g2_antennanp ANTENNA_117 (.A(_05012_));
 sg13g2_antennanp ANTENNA_118 (.A(_05024_));
 sg13g2_antennanp ANTENNA_119 (.A(_05024_));
 sg13g2_antennanp ANTENNA_120 (.A(_05047_));
 sg13g2_antennanp ANTENNA_121 (.A(_05047_));
 sg13g2_antennanp ANTENNA_122 (.A(_05047_));
 sg13g2_antennanp ANTENNA_123 (.A(_05047_));
 sg13g2_antennanp ANTENNA_124 (.A(_05100_));
 sg13g2_antennanp ANTENNA_125 (.A(_05101_));
 sg13g2_antennanp ANTENNA_126 (.A(_05101_));
 sg13g2_antennanp ANTENNA_127 (.A(_05101_));
 sg13g2_antennanp ANTENNA_128 (.A(_05101_));
 sg13g2_antennanp ANTENNA_129 (.A(_05101_));
 sg13g2_antennanp ANTENNA_130 (.A(_05101_));
 sg13g2_antennanp ANTENNA_131 (.A(_05102_));
 sg13g2_antennanp ANTENNA_132 (.A(_05118_));
 sg13g2_antennanp ANTENNA_133 (.A(_05124_));
 sg13g2_antennanp ANTENNA_134 (.A(_05128_));
 sg13g2_antennanp ANTENNA_135 (.A(_05130_));
 sg13g2_antennanp ANTENNA_136 (.A(_05130_));
 sg13g2_antennanp ANTENNA_137 (.A(_05130_));
 sg13g2_antennanp ANTENNA_138 (.A(_05130_));
 sg13g2_antennanp ANTENNA_139 (.A(_05130_));
 sg13g2_antennanp ANTENNA_140 (.A(_05130_));
 sg13g2_antennanp ANTENNA_141 (.A(_05130_));
 sg13g2_antennanp ANTENNA_142 (.A(_05130_));
 sg13g2_antennanp ANTENNA_143 (.A(_05130_));
 sg13g2_antennanp ANTENNA_144 (.A(_05130_));
 sg13g2_antennanp ANTENNA_145 (.A(_05134_));
 sg13g2_antennanp ANTENNA_146 (.A(_05134_));
 sg13g2_antennanp ANTENNA_147 (.A(_05134_));
 sg13g2_antennanp ANTENNA_148 (.A(_05134_));
 sg13g2_antennanp ANTENNA_149 (.A(_05134_));
 sg13g2_antennanp ANTENNA_150 (.A(_05134_));
 sg13g2_antennanp ANTENNA_151 (.A(_05134_));
 sg13g2_antennanp ANTENNA_152 (.A(_05134_));
 sg13g2_antennanp ANTENNA_153 (.A(_05134_));
 sg13g2_antennanp ANTENNA_154 (.A(_05136_));
 sg13g2_antennanp ANTENNA_155 (.A(_05164_));
 sg13g2_antennanp ANTENNA_156 (.A(_05164_));
 sg13g2_antennanp ANTENNA_157 (.A(_05164_));
 sg13g2_antennanp ANTENNA_158 (.A(_05171_));
 sg13g2_antennanp ANTENNA_159 (.A(_05171_));
 sg13g2_antennanp ANTENNA_160 (.A(_05171_));
 sg13g2_antennanp ANTENNA_161 (.A(_05198_));
 sg13g2_antennanp ANTENNA_162 (.A(_05201_));
 sg13g2_antennanp ANTENNA_163 (.A(_05201_));
 sg13g2_antennanp ANTENNA_164 (.A(_05201_));
 sg13g2_antennanp ANTENNA_165 (.A(_05201_));
 sg13g2_antennanp ANTENNA_166 (.A(_05201_));
 sg13g2_antennanp ANTENNA_167 (.A(_05201_));
 sg13g2_antennanp ANTENNA_168 (.A(_05201_));
 sg13g2_antennanp ANTENNA_169 (.A(_05205_));
 sg13g2_antennanp ANTENNA_170 (.A(_05209_));
 sg13g2_antennanp ANTENNA_171 (.A(_05238_));
 sg13g2_antennanp ANTENNA_172 (.A(_05238_));
 sg13g2_antennanp ANTENNA_173 (.A(_05238_));
 sg13g2_antennanp ANTENNA_174 (.A(_05238_));
 sg13g2_antennanp ANTENNA_175 (.A(_05252_));
 sg13g2_antennanp ANTENNA_176 (.A(_05258_));
 sg13g2_antennanp ANTENNA_177 (.A(_05286_));
 sg13g2_antennanp ANTENNA_178 (.A(_05286_));
 sg13g2_antennanp ANTENNA_179 (.A(_05302_));
 sg13g2_antennanp ANTENNA_180 (.A(_05302_));
 sg13g2_antennanp ANTENNA_181 (.A(_05302_));
 sg13g2_antennanp ANTENNA_182 (.A(_05302_));
 sg13g2_antennanp ANTENNA_183 (.A(_05302_));
 sg13g2_antennanp ANTENNA_184 (.A(_05302_));
 sg13g2_antennanp ANTENNA_185 (.A(_05302_));
 sg13g2_antennanp ANTENNA_186 (.A(_05302_));
 sg13g2_antennanp ANTENNA_187 (.A(_05302_));
 sg13g2_antennanp ANTENNA_188 (.A(_05309_));
 sg13g2_antennanp ANTENNA_189 (.A(_05309_));
 sg13g2_antennanp ANTENNA_190 (.A(_05309_));
 sg13g2_antennanp ANTENNA_191 (.A(_05309_));
 sg13g2_antennanp ANTENNA_192 (.A(_05318_));
 sg13g2_antennanp ANTENNA_193 (.A(_05328_));
 sg13g2_antennanp ANTENNA_194 (.A(_05339_));
 sg13g2_antennanp ANTENNA_195 (.A(_05342_));
 sg13g2_antennanp ANTENNA_196 (.A(_05342_));
 sg13g2_antennanp ANTENNA_197 (.A(_05342_));
 sg13g2_antennanp ANTENNA_198 (.A(_05344_));
 sg13g2_antennanp ANTENNA_199 (.A(_05344_));
 sg13g2_antennanp ANTENNA_200 (.A(_05344_));
 sg13g2_antennanp ANTENNA_201 (.A(_05344_));
 sg13g2_antennanp ANTENNA_202 (.A(_05344_));
 sg13g2_antennanp ANTENNA_203 (.A(_05344_));
 sg13g2_antennanp ANTENNA_204 (.A(_05344_));
 sg13g2_antennanp ANTENNA_205 (.A(_05344_));
 sg13g2_antennanp ANTENNA_206 (.A(_05344_));
 sg13g2_antennanp ANTENNA_207 (.A(_05346_));
 sg13g2_antennanp ANTENNA_208 (.A(_05350_));
 sg13g2_antennanp ANTENNA_209 (.A(_05377_));
 sg13g2_antennanp ANTENNA_210 (.A(_05377_));
 sg13g2_antennanp ANTENNA_211 (.A(_05377_));
 sg13g2_antennanp ANTENNA_212 (.A(_05377_));
 sg13g2_antennanp ANTENNA_213 (.A(_05389_));
 sg13g2_antennanp ANTENNA_214 (.A(_05390_));
 sg13g2_antennanp ANTENNA_215 (.A(_05404_));
 sg13g2_antennanp ANTENNA_216 (.A(_05415_));
 sg13g2_antennanp ANTENNA_217 (.A(_05424_));
 sg13g2_antennanp ANTENNA_218 (.A(_05424_));
 sg13g2_antennanp ANTENNA_219 (.A(_05424_));
 sg13g2_antennanp ANTENNA_220 (.A(_05424_));
 sg13g2_antennanp ANTENNA_221 (.A(_05442_));
 sg13g2_antennanp ANTENNA_222 (.A(_05459_));
 sg13g2_antennanp ANTENNA_223 (.A(_05477_));
 sg13g2_antennanp ANTENNA_224 (.A(_05485_));
 sg13g2_antennanp ANTENNA_225 (.A(_05485_));
 sg13g2_antennanp ANTENNA_226 (.A(_05485_));
 sg13g2_antennanp ANTENNA_227 (.A(_05500_));
 sg13g2_antennanp ANTENNA_228 (.A(_05524_));
 sg13g2_antennanp ANTENNA_229 (.A(_05576_));
 sg13g2_antennanp ANTENNA_230 (.A(_05584_));
 sg13g2_antennanp ANTENNA_231 (.A(_05584_));
 sg13g2_antennanp ANTENNA_232 (.A(_05591_));
 sg13g2_antennanp ANTENNA_233 (.A(_05591_));
 sg13g2_antennanp ANTENNA_234 (.A(_05591_));
 sg13g2_antennanp ANTENNA_235 (.A(_05609_));
 sg13g2_antennanp ANTENNA_236 (.A(_05609_));
 sg13g2_antennanp ANTENNA_237 (.A(_05609_));
 sg13g2_antennanp ANTENNA_238 (.A(_05609_));
 sg13g2_antennanp ANTENNA_239 (.A(_05611_));
 sg13g2_antennanp ANTENNA_240 (.A(_05633_));
 sg13g2_antennanp ANTENNA_241 (.A(_05657_));
 sg13g2_antennanp ANTENNA_242 (.A(_05670_));
 sg13g2_antennanp ANTENNA_243 (.A(_05681_));
 sg13g2_antennanp ANTENNA_244 (.A(_05681_));
 sg13g2_antennanp ANTENNA_245 (.A(_05705_));
 sg13g2_antennanp ANTENNA_246 (.A(_05705_));
 sg13g2_antennanp ANTENNA_247 (.A(_05705_));
 sg13g2_antennanp ANTENNA_248 (.A(_05726_));
 sg13g2_antennanp ANTENNA_249 (.A(_05750_));
 sg13g2_antennanp ANTENNA_250 (.A(_05777_));
 sg13g2_antennanp ANTENNA_251 (.A(_05814_));
 sg13g2_antennanp ANTENNA_252 (.A(_05816_));
 sg13g2_antennanp ANTENNA_253 (.A(_05818_));
 sg13g2_antennanp ANTENNA_254 (.A(_05827_));
 sg13g2_antennanp ANTENNA_255 (.A(_05829_));
 sg13g2_antennanp ANTENNA_256 (.A(_05874_));
 sg13g2_antennanp ANTENNA_257 (.A(_05886_));
 sg13g2_antennanp ANTENNA_258 (.A(_05890_));
 sg13g2_antennanp ANTENNA_259 (.A(_05897_));
 sg13g2_antennanp ANTENNA_260 (.A(_05904_));
 sg13g2_antennanp ANTENNA_261 (.A(_05924_));
 sg13g2_antennanp ANTENNA_262 (.A(_05924_));
 sg13g2_antennanp ANTENNA_263 (.A(_05939_));
 sg13g2_antennanp ANTENNA_264 (.A(_05946_));
 sg13g2_antennanp ANTENNA_265 (.A(_05951_));
 sg13g2_antennanp ANTENNA_266 (.A(_05951_));
 sg13g2_antennanp ANTENNA_267 (.A(_05957_));
 sg13g2_antennanp ANTENNA_268 (.A(_05997_));
 sg13g2_antennanp ANTENNA_269 (.A(_05998_));
 sg13g2_antennanp ANTENNA_270 (.A(_06018_));
 sg13g2_antennanp ANTENNA_271 (.A(_06023_));
 sg13g2_antennanp ANTENNA_272 (.A(_06046_));
 sg13g2_antennanp ANTENNA_273 (.A(_06050_));
 sg13g2_antennanp ANTENNA_274 (.A(_06053_));
 sg13g2_antennanp ANTENNA_275 (.A(_06053_));
 sg13g2_antennanp ANTENNA_276 (.A(_06064_));
 sg13g2_antennanp ANTENNA_277 (.A(_06075_));
 sg13g2_antennanp ANTENNA_278 (.A(_06083_));
 sg13g2_antennanp ANTENNA_279 (.A(_06091_));
 sg13g2_antennanp ANTENNA_280 (.A(_06116_));
 sg13g2_antennanp ANTENNA_281 (.A(_06134_));
 sg13g2_antennanp ANTENNA_282 (.A(_06139_));
 sg13g2_antennanp ANTENNA_283 (.A(_06146_));
 sg13g2_antennanp ANTENNA_284 (.A(_06146_));
 sg13g2_antennanp ANTENNA_285 (.A(_06146_));
 sg13g2_antennanp ANTENNA_286 (.A(_06151_));
 sg13g2_antennanp ANTENNA_287 (.A(_06167_));
 sg13g2_antennanp ANTENNA_288 (.A(_06179_));
 sg13g2_antennanp ANTENNA_289 (.A(_06189_));
 sg13g2_antennanp ANTENNA_290 (.A(_06196_));
 sg13g2_antennanp ANTENNA_291 (.A(_06209_));
 sg13g2_antennanp ANTENNA_292 (.A(_06225_));
 sg13g2_antennanp ANTENNA_293 (.A(_06227_));
 sg13g2_antennanp ANTENNA_294 (.A(_06244_));
 sg13g2_antennanp ANTENNA_295 (.A(_06249_));
 sg13g2_antennanp ANTENNA_296 (.A(_06250_));
 sg13g2_antennanp ANTENNA_297 (.A(_06271_));
 sg13g2_antennanp ANTENNA_298 (.A(_06281_));
 sg13g2_antennanp ANTENNA_299 (.A(_06290_));
 sg13g2_antennanp ANTENNA_300 (.A(_06300_));
 sg13g2_antennanp ANTENNA_301 (.A(_06322_));
 sg13g2_antennanp ANTENNA_302 (.A(_06324_));
 sg13g2_antennanp ANTENNA_303 (.A(_06328_));
 sg13g2_antennanp ANTENNA_304 (.A(_06334_));
 sg13g2_antennanp ANTENNA_305 (.A(_06335_));
 sg13g2_antennanp ANTENNA_306 (.A(_06342_));
 sg13g2_antennanp ANTENNA_307 (.A(_06347_));
 sg13g2_antennanp ANTENNA_308 (.A(_06351_));
 sg13g2_antennanp ANTENNA_309 (.A(_06361_));
 sg13g2_antennanp ANTENNA_310 (.A(_06366_));
 sg13g2_antennanp ANTENNA_311 (.A(_06372_));
 sg13g2_antennanp ANTENNA_312 (.A(_06374_));
 sg13g2_antennanp ANTENNA_313 (.A(_06383_));
 sg13g2_antennanp ANTENNA_314 (.A(_06391_));
 sg13g2_antennanp ANTENNA_315 (.A(_06396_));
 sg13g2_antennanp ANTENNA_316 (.A(_06396_));
 sg13g2_antennanp ANTENNA_317 (.A(_06397_));
 sg13g2_antennanp ANTENNA_318 (.A(_06417_));
 sg13g2_antennanp ANTENNA_319 (.A(_06422_));
 sg13g2_antennanp ANTENNA_320 (.A(_06440_));
 sg13g2_antennanp ANTENNA_321 (.A(_06448_));
 sg13g2_antennanp ANTENNA_322 (.A(_06463_));
 sg13g2_antennanp ANTENNA_323 (.A(_06467_));
 sg13g2_antennanp ANTENNA_324 (.A(_06484_));
 sg13g2_antennanp ANTENNA_325 (.A(_06492_));
 sg13g2_antennanp ANTENNA_326 (.A(_06497_));
 sg13g2_antennanp ANTENNA_327 (.A(_06504_));
 sg13g2_antennanp ANTENNA_328 (.A(_06506_));
 sg13g2_antennanp ANTENNA_329 (.A(_06512_));
 sg13g2_antennanp ANTENNA_330 (.A(_06517_));
 sg13g2_antennanp ANTENNA_331 (.A(_06522_));
 sg13g2_antennanp ANTENNA_332 (.A(_06523_));
 sg13g2_antennanp ANTENNA_333 (.A(_06546_));
 sg13g2_antennanp ANTENNA_334 (.A(_06548_));
 sg13g2_antennanp ANTENNA_335 (.A(_06559_));
 sg13g2_antennanp ANTENNA_336 (.A(_06588_));
 sg13g2_antennanp ANTENNA_337 (.A(_06589_));
 sg13g2_antennanp ANTENNA_338 (.A(_06594_));
 sg13g2_antennanp ANTENNA_339 (.A(_06596_));
 sg13g2_antennanp ANTENNA_340 (.A(_06621_));
 sg13g2_antennanp ANTENNA_341 (.A(_06640_));
 sg13g2_antennanp ANTENNA_342 (.A(_06658_));
 sg13g2_antennanp ANTENNA_343 (.A(_06667_));
 sg13g2_antennanp ANTENNA_344 (.A(_06679_));
 sg13g2_antennanp ANTENNA_345 (.A(_06680_));
 sg13g2_antennanp ANTENNA_346 (.A(_06682_));
 sg13g2_antennanp ANTENNA_347 (.A(_06684_));
 sg13g2_antennanp ANTENNA_348 (.A(_06687_));
 sg13g2_antennanp ANTENNA_349 (.A(_06688_));
 sg13g2_antennanp ANTENNA_350 (.A(_06701_));
 sg13g2_antennanp ANTENNA_351 (.A(_06702_));
 sg13g2_antennanp ANTENNA_352 (.A(_06712_));
 sg13g2_antennanp ANTENNA_353 (.A(_06732_));
 sg13g2_antennanp ANTENNA_354 (.A(_06745_));
 sg13g2_antennanp ANTENNA_355 (.A(_06758_));
 sg13g2_antennanp ANTENNA_356 (.A(_06761_));
 sg13g2_antennanp ANTENNA_357 (.A(_06764_));
 sg13g2_antennanp ANTENNA_358 (.A(_06768_));
 sg13g2_antennanp ANTENNA_359 (.A(_06775_));
 sg13g2_antennanp ANTENNA_360 (.A(_06796_));
 sg13g2_antennanp ANTENNA_361 (.A(_06813_));
 sg13g2_antennanp ANTENNA_362 (.A(_06830_));
 sg13g2_antennanp ANTENNA_363 (.A(_06830_));
 sg13g2_antennanp ANTENNA_364 (.A(_06834_));
 sg13g2_antennanp ANTENNA_365 (.A(_06844_));
 sg13g2_antennanp ANTENNA_366 (.A(_06849_));
 sg13g2_antennanp ANTENNA_367 (.A(_06926_));
 sg13g2_antennanp ANTENNA_368 (.A(_06926_));
 sg13g2_antennanp ANTENNA_369 (.A(_06959_));
 sg13g2_antennanp ANTENNA_370 (.A(_07004_));
 sg13g2_antennanp ANTENNA_371 (.A(_07022_));
 sg13g2_antennanp ANTENNA_372 (.A(_07040_));
 sg13g2_antennanp ANTENNA_373 (.A(_07057_));
 sg13g2_antennanp ANTENNA_374 (.A(_07071_));
 sg13g2_antennanp ANTENNA_375 (.A(_07085_));
 sg13g2_antennanp ANTENNA_376 (.A(_07098_));
 sg13g2_antennanp ANTENNA_377 (.A(_07111_));
 sg13g2_antennanp ANTENNA_378 (.A(_07154_));
 sg13g2_antennanp ANTENNA_379 (.A(_07170_));
 sg13g2_antennanp ANTENNA_380 (.A(_07243_));
 sg13g2_antennanp ANTENNA_381 (.A(_07258_));
 sg13g2_antennanp ANTENNA_382 (.A(_07273_));
 sg13g2_antennanp ANTENNA_383 (.A(_07301_));
 sg13g2_antennanp ANTENNA_384 (.A(_07316_));
 sg13g2_antennanp ANTENNA_385 (.A(_07331_));
 sg13g2_antennanp ANTENNA_386 (.A(_07534_));
 sg13g2_antennanp ANTENNA_387 (.A(_07534_));
 sg13g2_antennanp ANTENNA_388 (.A(_07534_));
 sg13g2_antennanp ANTENNA_389 (.A(_07534_));
 sg13g2_antennanp ANTENNA_390 (.A(_07534_));
 sg13g2_antennanp ANTENNA_391 (.A(_07534_));
 sg13g2_antennanp ANTENNA_392 (.A(_07534_));
 sg13g2_antennanp ANTENNA_393 (.A(_07534_));
 sg13g2_antennanp ANTENNA_394 (.A(_07534_));
 sg13g2_antennanp ANTENNA_395 (.A(_07663_));
 sg13g2_antennanp ANTENNA_396 (.A(_09082_));
 sg13g2_antennanp ANTENNA_397 (.A(_09082_));
 sg13g2_antennanp ANTENNA_398 (.A(_09082_));
 sg13g2_antennanp ANTENNA_399 (.A(_09082_));
 sg13g2_antennanp ANTENNA_400 (.A(_09082_));
 sg13g2_antennanp ANTENNA_401 (.A(_09082_));
 sg13g2_antennanp ANTENNA_402 (.A(_09082_));
 sg13g2_antennanp ANTENNA_403 (.A(_09082_));
 sg13g2_antennanp ANTENNA_404 (.A(_09082_));
 sg13g2_antennanp ANTENNA_405 (.A(_09082_));
 sg13g2_antennanp ANTENNA_406 (.A(_09082_));
 sg13g2_antennanp ANTENNA_407 (.A(_09082_));
 sg13g2_antennanp ANTENNA_408 (.A(_09082_));
 sg13g2_antennanp ANTENNA_409 (.A(_09082_));
 sg13g2_antennanp ANTENNA_410 (.A(_09104_));
 sg13g2_antennanp ANTENNA_411 (.A(_09104_));
 sg13g2_antennanp ANTENNA_412 (.A(_09104_));
 sg13g2_antennanp ANTENNA_413 (.A(_09104_));
 sg13g2_antennanp ANTENNA_414 (.A(_09301_));
 sg13g2_antennanp ANTENNA_415 (.A(_09301_));
 sg13g2_antennanp ANTENNA_416 (.A(_09301_));
 sg13g2_antennanp ANTENNA_417 (.A(_09301_));
 sg13g2_antennanp ANTENNA_418 (.A(_09301_));
 sg13g2_antennanp ANTENNA_419 (.A(_09301_));
 sg13g2_antennanp ANTENNA_420 (.A(_09436_));
 sg13g2_antennanp ANTENNA_421 (.A(_09436_));
 sg13g2_antennanp ANTENNA_422 (.A(_09436_));
 sg13g2_antennanp ANTENNA_423 (.A(_09573_));
 sg13g2_antennanp ANTENNA_424 (.A(_09573_));
 sg13g2_antennanp ANTENNA_425 (.A(_09573_));
 sg13g2_antennanp ANTENNA_426 (.A(_09573_));
 sg13g2_antennanp ANTENNA_427 (.A(_09599_));
 sg13g2_antennanp ANTENNA_428 (.A(_09599_));
 sg13g2_antennanp ANTENNA_429 (.A(_09599_));
 sg13g2_antennanp ANTENNA_430 (.A(_09599_));
 sg13g2_antennanp ANTENNA_431 (.A(_09910_));
 sg13g2_antennanp ANTENNA_432 (.A(_09910_));
 sg13g2_antennanp ANTENNA_433 (.A(_09910_));
 sg13g2_antennanp ANTENNA_434 (.A(_09910_));
 sg13g2_antennanp ANTENNA_435 (.A(_09910_));
 sg13g2_antennanp ANTENNA_436 (.A(_09910_));
 sg13g2_antennanp ANTENNA_437 (.A(_09910_));
 sg13g2_antennanp ANTENNA_438 (.A(_09910_));
 sg13g2_antennanp ANTENNA_439 (.A(_09910_));
 sg13g2_antennanp ANTENNA_440 (.A(_09910_));
 sg13g2_antennanp ANTENNA_441 (.A(_09944_));
 sg13g2_antennanp ANTENNA_442 (.A(_09944_));
 sg13g2_antennanp ANTENNA_443 (.A(_09944_));
 sg13g2_antennanp ANTENNA_444 (.A(_09944_));
 sg13g2_antennanp ANTENNA_445 (.A(_09944_));
 sg13g2_antennanp ANTENNA_446 (.A(_09944_));
 sg13g2_antennanp ANTENNA_447 (.A(_09944_));
 sg13g2_antennanp ANTENNA_448 (.A(_09944_));
 sg13g2_antennanp ANTENNA_449 (.A(_09944_));
 sg13g2_antennanp ANTENNA_450 (.A(_09944_));
 sg13g2_antennanp ANTENNA_451 (.A(_09960_));
 sg13g2_antennanp ANTENNA_452 (.A(_09960_));
 sg13g2_antennanp ANTENNA_453 (.A(_09960_));
 sg13g2_antennanp ANTENNA_454 (.A(_09960_));
 sg13g2_antennanp ANTENNA_455 (.A(_10009_));
 sg13g2_antennanp ANTENNA_456 (.A(_10009_));
 sg13g2_antennanp ANTENNA_457 (.A(_10009_));
 sg13g2_antennanp ANTENNA_458 (.A(_10009_));
 sg13g2_antennanp ANTENNA_459 (.A(_10009_));
 sg13g2_antennanp ANTENNA_460 (.A(_10009_));
 sg13g2_antennanp ANTENNA_461 (.A(_10009_));
 sg13g2_antennanp ANTENNA_462 (.A(_10009_));
 sg13g2_antennanp ANTENNA_463 (.A(_10009_));
 sg13g2_antennanp ANTENNA_464 (.A(_10032_));
 sg13g2_antennanp ANTENNA_465 (.A(_10032_));
 sg13g2_antennanp ANTENNA_466 (.A(_10032_));
 sg13g2_antennanp ANTENNA_467 (.A(_10032_));
 sg13g2_antennanp ANTENNA_468 (.A(_10032_));
 sg13g2_antennanp ANTENNA_469 (.A(_10032_));
 sg13g2_antennanp ANTENNA_470 (.A(_10032_));
 sg13g2_antennanp ANTENNA_471 (.A(_10032_));
 sg13g2_antennanp ANTENNA_472 (.A(_10032_));
 sg13g2_antennanp ANTENNA_473 (.A(_10032_));
 sg13g2_antennanp ANTENNA_474 (.A(_10074_));
 sg13g2_antennanp ANTENNA_475 (.A(_10074_));
 sg13g2_antennanp ANTENNA_476 (.A(_10074_));
 sg13g2_antennanp ANTENNA_477 (.A(_10074_));
 sg13g2_antennanp ANTENNA_478 (.A(_10077_));
 sg13g2_antennanp ANTENNA_479 (.A(_10077_));
 sg13g2_antennanp ANTENNA_480 (.A(_10077_));
 sg13g2_antennanp ANTENNA_481 (.A(_10085_));
 sg13g2_antennanp ANTENNA_482 (.A(_10085_));
 sg13g2_antennanp ANTENNA_483 (.A(_10085_));
 sg13g2_antennanp ANTENNA_484 (.A(_10085_));
 sg13g2_antennanp ANTENNA_485 (.A(_10085_));
 sg13g2_antennanp ANTENNA_486 (.A(_10085_));
 sg13g2_antennanp ANTENNA_487 (.A(_10085_));
 sg13g2_antennanp ANTENNA_488 (.A(_10085_));
 sg13g2_antennanp ANTENNA_489 (.A(_10085_));
 sg13g2_antennanp ANTENNA_490 (.A(_10092_));
 sg13g2_antennanp ANTENNA_491 (.A(_10092_));
 sg13g2_antennanp ANTENNA_492 (.A(_10092_));
 sg13g2_antennanp ANTENNA_493 (.A(_10092_));
 sg13g2_antennanp ANTENNA_494 (.A(_10092_));
 sg13g2_antennanp ANTENNA_495 (.A(_10107_));
 sg13g2_antennanp ANTENNA_496 (.A(_10107_));
 sg13g2_antennanp ANTENNA_497 (.A(_10107_));
 sg13g2_antennanp ANTENNA_498 (.A(_10107_));
 sg13g2_antennanp ANTENNA_499 (.A(_10151_));
 sg13g2_antennanp ANTENNA_500 (.A(_10151_));
 sg13g2_antennanp ANTENNA_501 (.A(_10151_));
 sg13g2_antennanp ANTENNA_502 (.A(_10404_));
 sg13g2_antennanp ANTENNA_503 (.A(_10404_));
 sg13g2_antennanp ANTENNA_504 (.A(_10404_));
 sg13g2_antennanp ANTENNA_505 (.A(_10404_));
 sg13g2_antennanp ANTENNA_506 (.A(_10435_));
 sg13g2_antennanp ANTENNA_507 (.A(_10435_));
 sg13g2_antennanp ANTENNA_508 (.A(_10435_));
 sg13g2_antennanp ANTENNA_509 (.A(_10435_));
 sg13g2_antennanp ANTENNA_510 (.A(_10439_));
 sg13g2_antennanp ANTENNA_511 (.A(_10439_));
 sg13g2_antennanp ANTENNA_512 (.A(_10439_));
 sg13g2_antennanp ANTENNA_513 (.A(_10439_));
 sg13g2_antennanp ANTENNA_514 (.A(_10441_));
 sg13g2_antennanp ANTENNA_515 (.A(_10441_));
 sg13g2_antennanp ANTENNA_516 (.A(_10441_));
 sg13g2_antennanp ANTENNA_517 (.A(_10441_));
 sg13g2_antennanp ANTENNA_518 (.A(_10460_));
 sg13g2_antennanp ANTENNA_519 (.A(_10460_));
 sg13g2_antennanp ANTENNA_520 (.A(_10460_));
 sg13g2_antennanp ANTENNA_521 (.A(_10460_));
 sg13g2_antennanp ANTENNA_522 (.A(_10831_));
 sg13g2_antennanp ANTENNA_523 (.A(_10831_));
 sg13g2_antennanp ANTENNA_524 (.A(_10831_));
 sg13g2_antennanp ANTENNA_525 (.A(_10831_));
 sg13g2_antennanp ANTENNA_526 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_527 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_528 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_529 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_530 (.A(\top_ihp.oisc.regs[2][10] ));
 sg13g2_antennanp ANTENNA_531 (.A(\top_ihp.oisc.regs[2][10] ));
 sg13g2_antennanp ANTENNA_532 (.A(\top_ihp.oisc.regs[2][10] ));
 sg13g2_antennanp ANTENNA_533 (.A(\top_ihp.oisc.regs[2][10] ));
 sg13g2_antennanp ANTENNA_534 (.A(\top_ihp.oisc.regs[2][10] ));
 sg13g2_antennanp ANTENNA_535 (.A(\top_ihp.oisc.regs[2][10] ));
 sg13g2_antennanp ANTENNA_536 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_537 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_538 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_539 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_540 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_541 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_542 (.A(\top_ihp.oisc.regs[32][13] ));
 sg13g2_antennanp ANTENNA_543 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_544 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_545 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_546 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_547 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_548 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_549 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_550 (.A(\top_ihp.oisc.regs[32][18] ));
 sg13g2_antennanp ANTENNA_551 (.A(\top_ihp.oisc.regs[32][18] ));
 sg13g2_antennanp ANTENNA_552 (.A(\top_ihp.oisc.regs[32][18] ));
 sg13g2_antennanp ANTENNA_553 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_554 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_555 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_556 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_557 (.A(\top_ihp.oisc.regs[32][22] ));
 sg13g2_antennanp ANTENNA_558 (.A(\top_ihp.oisc.regs[32][22] ));
 sg13g2_antennanp ANTENNA_559 (.A(\top_ihp.oisc.regs[32][22] ));
 sg13g2_antennanp ANTENNA_560 (.A(\top_ihp.oisc.regs[32][22] ));
 sg13g2_antennanp ANTENNA_561 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_562 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_563 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_564 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_565 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_566 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_567 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_568 (.A(\top_ihp.oisc.regs[32][26] ));
 sg13g2_antennanp ANTENNA_569 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_570 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_571 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_572 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_573 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_574 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_575 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_576 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_577 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_578 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_579 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_580 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_581 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_582 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_583 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_584 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_585 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_586 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_587 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_588 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_589 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_590 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_591 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_592 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_593 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_594 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_595 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_596 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_597 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_598 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_599 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_600 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_601 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_602 (.A(\top_ihp.ram_cs_o ));
 sg13g2_antennanp ANTENNA_603 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_604 (.A(net1));
 sg13g2_antennanp ANTENNA_605 (.A(net1));
 sg13g2_antennanp ANTENNA_606 (.A(net1));
 sg13g2_antennanp ANTENNA_607 (.A(net9));
 sg13g2_antennanp ANTENNA_608 (.A(net47));
 sg13g2_antennanp ANTENNA_609 (.A(net47));
 sg13g2_antennanp ANTENNA_610 (.A(net47));
 sg13g2_antennanp ANTENNA_611 (.A(net47));
 sg13g2_antennanp ANTENNA_612 (.A(net47));
 sg13g2_antennanp ANTENNA_613 (.A(net47));
 sg13g2_antennanp ANTENNA_614 (.A(net47));
 sg13g2_antennanp ANTENNA_615 (.A(net47));
 sg13g2_antennanp ANTENNA_616 (.A(net47));
 sg13g2_antennanp ANTENNA_617 (.A(net47));
 sg13g2_antennanp ANTENNA_618 (.A(net47));
 sg13g2_antennanp ANTENNA_619 (.A(net47));
 sg13g2_antennanp ANTENNA_620 (.A(net47));
 sg13g2_antennanp ANTENNA_621 (.A(net47));
 sg13g2_antennanp ANTENNA_622 (.A(net47));
 sg13g2_antennanp ANTENNA_623 (.A(net47));
 sg13g2_antennanp ANTENNA_624 (.A(net55));
 sg13g2_antennanp ANTENNA_625 (.A(net55));
 sg13g2_antennanp ANTENNA_626 (.A(net55));
 sg13g2_antennanp ANTENNA_627 (.A(net55));
 sg13g2_antennanp ANTENNA_628 (.A(net55));
 sg13g2_antennanp ANTENNA_629 (.A(net55));
 sg13g2_antennanp ANTENNA_630 (.A(net55));
 sg13g2_antennanp ANTENNA_631 (.A(net55));
 sg13g2_antennanp ANTENNA_632 (.A(net55));
 sg13g2_antennanp ANTENNA_633 (.A(net70));
 sg13g2_antennanp ANTENNA_634 (.A(net70));
 sg13g2_antennanp ANTENNA_635 (.A(net70));
 sg13g2_antennanp ANTENNA_636 (.A(net70));
 sg13g2_antennanp ANTENNA_637 (.A(net70));
 sg13g2_antennanp ANTENNA_638 (.A(net70));
 sg13g2_antennanp ANTENNA_639 (.A(net70));
 sg13g2_antennanp ANTENNA_640 (.A(net70));
 sg13g2_antennanp ANTENNA_641 (.A(net70));
 sg13g2_antennanp ANTENNA_642 (.A(net70));
 sg13g2_antennanp ANTENNA_643 (.A(net70));
 sg13g2_antennanp ANTENNA_644 (.A(net70));
 sg13g2_antennanp ANTENNA_645 (.A(net70));
 sg13g2_antennanp ANTENNA_646 (.A(net70));
 sg13g2_antennanp ANTENNA_647 (.A(net70));
 sg13g2_antennanp ANTENNA_648 (.A(net87));
 sg13g2_antennanp ANTENNA_649 (.A(net87));
 sg13g2_antennanp ANTENNA_650 (.A(net87));
 sg13g2_antennanp ANTENNA_651 (.A(net87));
 sg13g2_antennanp ANTENNA_652 (.A(net87));
 sg13g2_antennanp ANTENNA_653 (.A(net87));
 sg13g2_antennanp ANTENNA_654 (.A(net87));
 sg13g2_antennanp ANTENNA_655 (.A(net87));
 sg13g2_antennanp ANTENNA_656 (.A(net87));
 sg13g2_antennanp ANTENNA_657 (.A(net136));
 sg13g2_antennanp ANTENNA_658 (.A(net136));
 sg13g2_antennanp ANTENNA_659 (.A(net136));
 sg13g2_antennanp ANTENNA_660 (.A(net136));
 sg13g2_antennanp ANTENNA_661 (.A(net136));
 sg13g2_antennanp ANTENNA_662 (.A(net136));
 sg13g2_antennanp ANTENNA_663 (.A(net136));
 sg13g2_antennanp ANTENNA_664 (.A(net136));
 sg13g2_antennanp ANTENNA_665 (.A(net136));
 sg13g2_antennanp ANTENNA_666 (.A(net136));
 sg13g2_antennanp ANTENNA_667 (.A(net136));
 sg13g2_antennanp ANTENNA_668 (.A(net136));
 sg13g2_antennanp ANTENNA_669 (.A(net139));
 sg13g2_antennanp ANTENNA_670 (.A(net139));
 sg13g2_antennanp ANTENNA_671 (.A(net139));
 sg13g2_antennanp ANTENNA_672 (.A(net139));
 sg13g2_antennanp ANTENNA_673 (.A(net139));
 sg13g2_antennanp ANTENNA_674 (.A(net139));
 sg13g2_antennanp ANTENNA_675 (.A(net139));
 sg13g2_antennanp ANTENNA_676 (.A(net139));
 sg13g2_antennanp ANTENNA_677 (.A(net139));
 sg13g2_antennanp ANTENNA_678 (.A(net139));
 sg13g2_antennanp ANTENNA_679 (.A(net139));
 sg13g2_antennanp ANTENNA_680 (.A(net139));
 sg13g2_antennanp ANTENNA_681 (.A(net139));
 sg13g2_antennanp ANTENNA_682 (.A(net139));
 sg13g2_antennanp ANTENNA_683 (.A(net142));
 sg13g2_antennanp ANTENNA_684 (.A(net142));
 sg13g2_antennanp ANTENNA_685 (.A(net142));
 sg13g2_antennanp ANTENNA_686 (.A(net142));
 sg13g2_antennanp ANTENNA_687 (.A(net142));
 sg13g2_antennanp ANTENNA_688 (.A(net142));
 sg13g2_antennanp ANTENNA_689 (.A(net142));
 sg13g2_antennanp ANTENNA_690 (.A(net142));
 sg13g2_antennanp ANTENNA_691 (.A(net142));
 sg13g2_antennanp ANTENNA_692 (.A(net142));
 sg13g2_antennanp ANTENNA_693 (.A(net142));
 sg13g2_antennanp ANTENNA_694 (.A(net142));
 sg13g2_antennanp ANTENNA_695 (.A(net142));
 sg13g2_antennanp ANTENNA_696 (.A(net142));
 sg13g2_antennanp ANTENNA_697 (.A(net142));
 sg13g2_antennanp ANTENNA_698 (.A(net142));
 sg13g2_antennanp ANTENNA_699 (.A(net142));
 sg13g2_antennanp ANTENNA_700 (.A(net142));
 sg13g2_antennanp ANTENNA_701 (.A(net142));
 sg13g2_antennanp ANTENNA_702 (.A(net142));
 sg13g2_antennanp ANTENNA_703 (.A(net235));
 sg13g2_antennanp ANTENNA_704 (.A(net235));
 sg13g2_antennanp ANTENNA_705 (.A(net235));
 sg13g2_antennanp ANTENNA_706 (.A(net235));
 sg13g2_antennanp ANTENNA_707 (.A(net235));
 sg13g2_antennanp ANTENNA_708 (.A(net235));
 sg13g2_antennanp ANTENNA_709 (.A(net235));
 sg13g2_antennanp ANTENNA_710 (.A(net235));
 sg13g2_antennanp ANTENNA_711 (.A(net235));
 sg13g2_antennanp ANTENNA_712 (.A(net235));
 sg13g2_antennanp ANTENNA_713 (.A(net235));
 sg13g2_antennanp ANTENNA_714 (.A(net235));
 sg13g2_antennanp ANTENNA_715 (.A(net236));
 sg13g2_antennanp ANTENNA_716 (.A(net236));
 sg13g2_antennanp ANTENNA_717 (.A(net236));
 sg13g2_antennanp ANTENNA_718 (.A(net236));
 sg13g2_antennanp ANTENNA_719 (.A(net236));
 sg13g2_antennanp ANTENNA_720 (.A(net236));
 sg13g2_antennanp ANTENNA_721 (.A(net236));
 sg13g2_antennanp ANTENNA_722 (.A(net236));
 sg13g2_antennanp ANTENNA_723 (.A(net236));
 sg13g2_antennanp ANTENNA_724 (.A(net236));
 sg13g2_antennanp ANTENNA_725 (.A(net236));
 sg13g2_antennanp ANTENNA_726 (.A(net255));
 sg13g2_antennanp ANTENNA_727 (.A(net255));
 sg13g2_antennanp ANTENNA_728 (.A(net255));
 sg13g2_antennanp ANTENNA_729 (.A(net255));
 sg13g2_antennanp ANTENNA_730 (.A(net255));
 sg13g2_antennanp ANTENNA_731 (.A(net255));
 sg13g2_antennanp ANTENNA_732 (.A(net255));
 sg13g2_antennanp ANTENNA_733 (.A(net255));
 sg13g2_antennanp ANTENNA_734 (.A(net255));
 sg13g2_antennanp ANTENNA_735 (.A(net255));
 sg13g2_antennanp ANTENNA_736 (.A(net255));
 sg13g2_antennanp ANTENNA_737 (.A(net255));
 sg13g2_antennanp ANTENNA_738 (.A(net255));
 sg13g2_antennanp ANTENNA_739 (.A(net347));
 sg13g2_antennanp ANTENNA_740 (.A(net347));
 sg13g2_antennanp ANTENNA_741 (.A(net347));
 sg13g2_antennanp ANTENNA_742 (.A(net347));
 sg13g2_antennanp ANTENNA_743 (.A(net347));
 sg13g2_antennanp ANTENNA_744 (.A(net347));
 sg13g2_antennanp ANTENNA_745 (.A(net347));
 sg13g2_antennanp ANTENNA_746 (.A(net347));
 sg13g2_antennanp ANTENNA_747 (.A(net413));
 sg13g2_antennanp ANTENNA_748 (.A(net413));
 sg13g2_antennanp ANTENNA_749 (.A(net413));
 sg13g2_antennanp ANTENNA_750 (.A(net413));
 sg13g2_antennanp ANTENNA_751 (.A(net413));
 sg13g2_antennanp ANTENNA_752 (.A(net413));
 sg13g2_antennanp ANTENNA_753 (.A(net413));
 sg13g2_antennanp ANTENNA_754 (.A(net413));
 sg13g2_antennanp ANTENNA_755 (.A(net413));
 sg13g2_antennanp ANTENNA_756 (.A(net413));
 sg13g2_antennanp ANTENNA_757 (.A(net413));
 sg13g2_antennanp ANTENNA_758 (.A(net413));
 sg13g2_antennanp ANTENNA_759 (.A(net413));
 sg13g2_antennanp ANTENNA_760 (.A(net413));
 sg13g2_antennanp ANTENNA_761 (.A(net420));
 sg13g2_antennanp ANTENNA_762 (.A(net420));
 sg13g2_antennanp ANTENNA_763 (.A(net420));
 sg13g2_antennanp ANTENNA_764 (.A(net420));
 sg13g2_antennanp ANTENNA_765 (.A(net420));
 sg13g2_antennanp ANTENNA_766 (.A(net420));
 sg13g2_antennanp ANTENNA_767 (.A(net420));
 sg13g2_antennanp ANTENNA_768 (.A(net420));
 sg13g2_antennanp ANTENNA_769 (.A(net435));
 sg13g2_antennanp ANTENNA_770 (.A(net435));
 sg13g2_antennanp ANTENNA_771 (.A(net435));
 sg13g2_antennanp ANTENNA_772 (.A(net435));
 sg13g2_antennanp ANTENNA_773 (.A(net435));
 sg13g2_antennanp ANTENNA_774 (.A(net435));
 sg13g2_antennanp ANTENNA_775 (.A(net435));
 sg13g2_antennanp ANTENNA_776 (.A(net435));
 sg13g2_antennanp ANTENNA_777 (.A(net439));
 sg13g2_antennanp ANTENNA_778 (.A(net439));
 sg13g2_antennanp ANTENNA_779 (.A(net439));
 sg13g2_antennanp ANTENNA_780 (.A(net439));
 sg13g2_antennanp ANTENNA_781 (.A(net439));
 sg13g2_antennanp ANTENNA_782 (.A(net439));
 sg13g2_antennanp ANTENNA_783 (.A(net439));
 sg13g2_antennanp ANTENNA_784 (.A(net439));
 sg13g2_antennanp ANTENNA_785 (.A(net439));
 sg13g2_antennanp ANTENNA_786 (.A(net439));
 sg13g2_antennanp ANTENNA_787 (.A(net439));
 sg13g2_antennanp ANTENNA_788 (.A(net439));
 sg13g2_antennanp ANTENNA_789 (.A(net439));
 sg13g2_antennanp ANTENNA_790 (.A(net439));
 sg13g2_antennanp ANTENNA_791 (.A(net439));
 sg13g2_antennanp ANTENNA_792 (.A(net439));
 sg13g2_antennanp ANTENNA_793 (.A(net439));
 sg13g2_antennanp ANTENNA_794 (.A(net439));
 sg13g2_antennanp ANTENNA_795 (.A(net439));
 sg13g2_antennanp ANTENNA_796 (.A(net439));
 sg13g2_antennanp ANTENNA_797 (.A(net454));
 sg13g2_antennanp ANTENNA_798 (.A(net454));
 sg13g2_antennanp ANTENNA_799 (.A(net454));
 sg13g2_antennanp ANTENNA_800 (.A(net454));
 sg13g2_antennanp ANTENNA_801 (.A(net454));
 sg13g2_antennanp ANTENNA_802 (.A(net454));
 sg13g2_antennanp ANTENNA_803 (.A(net454));
 sg13g2_antennanp ANTENNA_804 (.A(net454));
 sg13g2_antennanp ANTENNA_805 (.A(net454));
 sg13g2_antennanp ANTENNA_806 (.A(net454));
 sg13g2_antennanp ANTENNA_807 (.A(net454));
 sg13g2_antennanp ANTENNA_808 (.A(net454));
 sg13g2_antennanp ANTENNA_809 (.A(net454));
 sg13g2_antennanp ANTENNA_810 (.A(net454));
 sg13g2_antennanp ANTENNA_811 (.A(net454));
 sg13g2_antennanp ANTENNA_812 (.A(net454));
 sg13g2_antennanp ANTENNA_813 (.A(net454));
 sg13g2_antennanp ANTENNA_814 (.A(net454));
 sg13g2_antennanp ANTENNA_815 (.A(net454));
 sg13g2_antennanp ANTENNA_816 (.A(net454));
 sg13g2_antennanp ANTENNA_817 (.A(net460));
 sg13g2_antennanp ANTENNA_818 (.A(net460));
 sg13g2_antennanp ANTENNA_819 (.A(net460));
 sg13g2_antennanp ANTENNA_820 (.A(net460));
 sg13g2_antennanp ANTENNA_821 (.A(net460));
 sg13g2_antennanp ANTENNA_822 (.A(net460));
 sg13g2_antennanp ANTENNA_823 (.A(net460));
 sg13g2_antennanp ANTENNA_824 (.A(net460));
 sg13g2_antennanp ANTENNA_825 (.A(net460));
 sg13g2_antennanp ANTENNA_826 (.A(net460));
 sg13g2_antennanp ANTENNA_827 (.A(net460));
 sg13g2_antennanp ANTENNA_828 (.A(net460));
 sg13g2_antennanp ANTENNA_829 (.A(net460));
 sg13g2_antennanp ANTENNA_830 (.A(net469));
 sg13g2_antennanp ANTENNA_831 (.A(net469));
 sg13g2_antennanp ANTENNA_832 (.A(net469));
 sg13g2_antennanp ANTENNA_833 (.A(net469));
 sg13g2_antennanp ANTENNA_834 (.A(net469));
 sg13g2_antennanp ANTENNA_835 (.A(net469));
 sg13g2_antennanp ANTENNA_836 (.A(net469));
 sg13g2_antennanp ANTENNA_837 (.A(net469));
 sg13g2_antennanp ANTENNA_838 (.A(net469));
 sg13g2_antennanp ANTENNA_839 (.A(net474));
 sg13g2_antennanp ANTENNA_840 (.A(net474));
 sg13g2_antennanp ANTENNA_841 (.A(net474));
 sg13g2_antennanp ANTENNA_842 (.A(net474));
 sg13g2_antennanp ANTENNA_843 (.A(net474));
 sg13g2_antennanp ANTENNA_844 (.A(net474));
 sg13g2_antennanp ANTENNA_845 (.A(net474));
 sg13g2_antennanp ANTENNA_846 (.A(net474));
 sg13g2_antennanp ANTENNA_847 (.A(net475));
 sg13g2_antennanp ANTENNA_848 (.A(net475));
 sg13g2_antennanp ANTENNA_849 (.A(net475));
 sg13g2_antennanp ANTENNA_850 (.A(net475));
 sg13g2_antennanp ANTENNA_851 (.A(net475));
 sg13g2_antennanp ANTENNA_852 (.A(net475));
 sg13g2_antennanp ANTENNA_853 (.A(net475));
 sg13g2_antennanp ANTENNA_854 (.A(net475));
 sg13g2_antennanp ANTENNA_855 (.A(net475));
 sg13g2_antennanp ANTENNA_856 (.A(net475));
 sg13g2_antennanp ANTENNA_857 (.A(net475));
 sg13g2_antennanp ANTENNA_858 (.A(net475));
 sg13g2_antennanp ANTENNA_859 (.A(net475));
 sg13g2_antennanp ANTENNA_860 (.A(net475));
 sg13g2_antennanp ANTENNA_861 (.A(net475));
 sg13g2_antennanp ANTENNA_862 (.A(net475));
 sg13g2_antennanp ANTENNA_863 (.A(net480));
 sg13g2_antennanp ANTENNA_864 (.A(net480));
 sg13g2_antennanp ANTENNA_865 (.A(net480));
 sg13g2_antennanp ANTENNA_866 (.A(net480));
 sg13g2_antennanp ANTENNA_867 (.A(net480));
 sg13g2_antennanp ANTENNA_868 (.A(net480));
 sg13g2_antennanp ANTENNA_869 (.A(net480));
 sg13g2_antennanp ANTENNA_870 (.A(net480));
 sg13g2_antennanp ANTENNA_871 (.A(net480));
 sg13g2_antennanp ANTENNA_872 (.A(net483));
 sg13g2_antennanp ANTENNA_873 (.A(net483));
 sg13g2_antennanp ANTENNA_874 (.A(net483));
 sg13g2_antennanp ANTENNA_875 (.A(net483));
 sg13g2_antennanp ANTENNA_876 (.A(net483));
 sg13g2_antennanp ANTENNA_877 (.A(net483));
 sg13g2_antennanp ANTENNA_878 (.A(net483));
 sg13g2_antennanp ANTENNA_879 (.A(net483));
 sg13g2_antennanp ANTENNA_880 (.A(net483));
 sg13g2_antennanp ANTENNA_881 (.A(net562));
 sg13g2_antennanp ANTENNA_882 (.A(net562));
 sg13g2_antennanp ANTENNA_883 (.A(net562));
 sg13g2_antennanp ANTENNA_884 (.A(net562));
 sg13g2_antennanp ANTENNA_885 (.A(net562));
 sg13g2_antennanp ANTENNA_886 (.A(net562));
 sg13g2_antennanp ANTENNA_887 (.A(net562));
 sg13g2_antennanp ANTENNA_888 (.A(net562));
 sg13g2_antennanp ANTENNA_889 (.A(net562));
 sg13g2_antennanp ANTENNA_890 (.A(net562));
 sg13g2_antennanp ANTENNA_891 (.A(net562));
 sg13g2_antennanp ANTENNA_892 (.A(net562));
 sg13g2_antennanp ANTENNA_893 (.A(net562));
 sg13g2_antennanp ANTENNA_894 (.A(net562));
 sg13g2_antennanp ANTENNA_895 (.A(net602));
 sg13g2_antennanp ANTENNA_896 (.A(net602));
 sg13g2_antennanp ANTENNA_897 (.A(net602));
 sg13g2_antennanp ANTENNA_898 (.A(net602));
 sg13g2_antennanp ANTENNA_899 (.A(net602));
 sg13g2_antennanp ANTENNA_900 (.A(net602));
 sg13g2_antennanp ANTENNA_901 (.A(net602));
 sg13g2_antennanp ANTENNA_902 (.A(net602));
 sg13g2_antennanp ANTENNA_903 (.A(net602));
 sg13g2_antennanp ANTENNA_904 (.A(net602));
 sg13g2_antennanp ANTENNA_905 (.A(net602));
 sg13g2_antennanp ANTENNA_906 (.A(net602));
 sg13g2_antennanp ANTENNA_907 (.A(net602));
 sg13g2_antennanp ANTENNA_908 (.A(net602));
 sg13g2_antennanp ANTENNA_909 (.A(net602));
 sg13g2_antennanp ANTENNA_910 (.A(net602));
 sg13g2_antennanp ANTENNA_911 (.A(net602));
 sg13g2_antennanp ANTENNA_912 (.A(net602));
 sg13g2_antennanp ANTENNA_913 (.A(net602));
 sg13g2_antennanp ANTENNA_914 (.A(net602));
 sg13g2_antennanp ANTENNA_915 (.A(net602));
 sg13g2_antennanp ANTENNA_916 (.A(net602));
 sg13g2_antennanp ANTENNA_917 (.A(net643));
 sg13g2_antennanp ANTENNA_918 (.A(net643));
 sg13g2_antennanp ANTENNA_919 (.A(net643));
 sg13g2_antennanp ANTENNA_920 (.A(net643));
 sg13g2_antennanp ANTENNA_921 (.A(net643));
 sg13g2_antennanp ANTENNA_922 (.A(net643));
 sg13g2_antennanp ANTENNA_923 (.A(net643));
 sg13g2_antennanp ANTENNA_924 (.A(net643));
 sg13g2_antennanp ANTENNA_925 (.A(net643));
 sg13g2_antennanp ANTENNA_926 (.A(net644));
 sg13g2_antennanp ANTENNA_927 (.A(net644));
 sg13g2_antennanp ANTENNA_928 (.A(net644));
 sg13g2_antennanp ANTENNA_929 (.A(net644));
 sg13g2_antennanp ANTENNA_930 (.A(net644));
 sg13g2_antennanp ANTENNA_931 (.A(net644));
 sg13g2_antennanp ANTENNA_932 (.A(net644));
 sg13g2_antennanp ANTENNA_933 (.A(net644));
 sg13g2_antennanp ANTENNA_934 (.A(net644));
 sg13g2_antennanp ANTENNA_935 (.A(net663));
 sg13g2_antennanp ANTENNA_936 (.A(net663));
 sg13g2_antennanp ANTENNA_937 (.A(net663));
 sg13g2_antennanp ANTENNA_938 (.A(net663));
 sg13g2_antennanp ANTENNA_939 (.A(net663));
 sg13g2_antennanp ANTENNA_940 (.A(net663));
 sg13g2_antennanp ANTENNA_941 (.A(net663));
 sg13g2_antennanp ANTENNA_942 (.A(net663));
 sg13g2_antennanp ANTENNA_943 (.A(net663));
 sg13g2_antennanp ANTENNA_944 (.A(net663));
 sg13g2_antennanp ANTENNA_945 (.A(net663));
 sg13g2_antennanp ANTENNA_946 (.A(net663));
 sg13g2_antennanp ANTENNA_947 (.A(net663));
 sg13g2_antennanp ANTENNA_948 (.A(net663));
 sg13g2_antennanp ANTENNA_949 (.A(net663));
 sg13g2_antennanp ANTENNA_950 (.A(net663));
 sg13g2_antennanp ANTENNA_951 (.A(net663));
 sg13g2_antennanp ANTENNA_952 (.A(net663));
 sg13g2_antennanp ANTENNA_953 (.A(net663));
 sg13g2_antennanp ANTENNA_954 (.A(net663));
 sg13g2_antennanp ANTENNA_955 (.A(net663));
 sg13g2_antennanp ANTENNA_956 (.A(net682));
 sg13g2_antennanp ANTENNA_957 (.A(net682));
 sg13g2_antennanp ANTENNA_958 (.A(net682));
 sg13g2_antennanp ANTENNA_959 (.A(net682));
 sg13g2_antennanp ANTENNA_960 (.A(net682));
 sg13g2_antennanp ANTENNA_961 (.A(net682));
 sg13g2_antennanp ANTENNA_962 (.A(net682));
 sg13g2_antennanp ANTENNA_963 (.A(net682));
 sg13g2_antennanp ANTENNA_964 (.A(net682));
 sg13g2_antennanp ANTENNA_965 (.A(net682));
 sg13g2_antennanp ANTENNA_966 (.A(net682));
 sg13g2_antennanp ANTENNA_967 (.A(net682));
 sg13g2_antennanp ANTENNA_968 (.A(net684));
 sg13g2_antennanp ANTENNA_969 (.A(net684));
 sg13g2_antennanp ANTENNA_970 (.A(net684));
 sg13g2_antennanp ANTENNA_971 (.A(net684));
 sg13g2_antennanp ANTENNA_972 (.A(net684));
 sg13g2_antennanp ANTENNA_973 (.A(net684));
 sg13g2_antennanp ANTENNA_974 (.A(net684));
 sg13g2_antennanp ANTENNA_975 (.A(net684));
 sg13g2_antennanp ANTENNA_976 (.A(net684));
 sg13g2_antennanp ANTENNA_977 (.A(net684));
 sg13g2_antennanp ANTENNA_978 (.A(net684));
 sg13g2_antennanp ANTENNA_979 (.A(net684));
 sg13g2_antennanp ANTENNA_980 (.A(net684));
 sg13g2_antennanp ANTENNA_981 (.A(net735));
 sg13g2_antennanp ANTENNA_982 (.A(net735));
 sg13g2_antennanp ANTENNA_983 (.A(net735));
 sg13g2_antennanp ANTENNA_984 (.A(net735));
 sg13g2_antennanp ANTENNA_985 (.A(net735));
 sg13g2_antennanp ANTENNA_986 (.A(net735));
 sg13g2_antennanp ANTENNA_987 (.A(net735));
 sg13g2_antennanp ANTENNA_988 (.A(net735));
 sg13g2_antennanp ANTENNA_989 (.A(net735));
 sg13g2_antennanp ANTENNA_990 (.A(_00294_));
 sg13g2_antennanp ANTENNA_991 (.A(_00294_));
 sg13g2_antennanp ANTENNA_992 (.A(_00296_));
 sg13g2_antennanp ANTENNA_993 (.A(_00299_));
 sg13g2_antennanp ANTENNA_994 (.A(_00299_));
 sg13g2_antennanp ANTENNA_995 (.A(_00299_));
 sg13g2_antennanp ANTENNA_996 (.A(_00300_));
 sg13g2_antennanp ANTENNA_997 (.A(_00305_));
 sg13g2_antennanp ANTENNA_998 (.A(_00307_));
 sg13g2_antennanp ANTENNA_999 (.A(_00307_));
 sg13g2_antennanp ANTENNA_1000 (.A(_00311_));
 sg13g2_antennanp ANTENNA_1001 (.A(_00311_));
 sg13g2_antennanp ANTENNA_1002 (.A(_00316_));
 sg13g2_antennanp ANTENNA_1003 (.A(_00319_));
 sg13g2_antennanp ANTENNA_1004 (.A(_00320_));
 sg13g2_antennanp ANTENNA_1005 (.A(_00322_));
 sg13g2_antennanp ANTENNA_1006 (.A(_00322_));
 sg13g2_antennanp ANTENNA_1007 (.A(_00323_));
 sg13g2_antennanp ANTENNA_1008 (.A(_00324_));
 sg13g2_antennanp ANTENNA_1009 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1010 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1011 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1012 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1013 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1014 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1015 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1016 (.A(_03014_));
 sg13g2_antennanp ANTENNA_1017 (.A(_03014_));
 sg13g2_antennanp ANTENNA_1018 (.A(_03014_));
 sg13g2_antennanp ANTENNA_1019 (.A(_03021_));
 sg13g2_antennanp ANTENNA_1020 (.A(_03021_));
 sg13g2_antennanp ANTENNA_1021 (.A(_03021_));
 sg13g2_antennanp ANTENNA_1022 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1023 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1024 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1025 (.A(_03108_));
 sg13g2_antennanp ANTENNA_1026 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1027 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1028 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1029 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1030 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1031 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1032 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1033 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1034 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1035 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1036 (.A(_03713_));
 sg13g2_antennanp ANTENNA_1037 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1038 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1039 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1040 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1041 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1042 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1043 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1044 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1045 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1046 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1047 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1048 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1049 (.A(_04857_));
 sg13g2_antennanp ANTENNA_1050 (.A(_04857_));
 sg13g2_antennanp ANTENNA_1051 (.A(_04871_));
 sg13g2_antennanp ANTENNA_1052 (.A(_04871_));
 sg13g2_antennanp ANTENNA_1053 (.A(_04871_));
 sg13g2_antennanp ANTENNA_1054 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1055 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1056 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1057 (.A(_04883_));
 sg13g2_antennanp ANTENNA_1058 (.A(_04912_));
 sg13g2_antennanp ANTENNA_1059 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1060 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1061 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1062 (.A(_04921_));
 sg13g2_antennanp ANTENNA_1063 (.A(_04921_));
 sg13g2_antennanp ANTENNA_1064 (.A(_04921_));
 sg13g2_antennanp ANTENNA_1065 (.A(_04932_));
 sg13g2_antennanp ANTENNA_1066 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1067 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1068 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1069 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1070 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1071 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1072 (.A(_05024_));
 sg13g2_antennanp ANTENNA_1073 (.A(_05100_));
 sg13g2_antennanp ANTENNA_1074 (.A(_05100_));
 sg13g2_antennanp ANTENNA_1075 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1076 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1077 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1078 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1079 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1080 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1081 (.A(_05102_));
 sg13g2_antennanp ANTENNA_1082 (.A(_05102_));
 sg13g2_antennanp ANTENNA_1083 (.A(_05118_));
 sg13g2_antennanp ANTENNA_1084 (.A(_05124_));
 sg13g2_antennanp ANTENNA_1085 (.A(_05124_));
 sg13g2_antennanp ANTENNA_1086 (.A(_05128_));
 sg13g2_antennanp ANTENNA_1087 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1088 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1089 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1090 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1091 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1092 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1093 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1094 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1095 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1096 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1097 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1098 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1099 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1100 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1101 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1102 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1103 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1104 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1105 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1106 (.A(_05136_));
 sg13g2_antennanp ANTENNA_1107 (.A(_05198_));
 sg13g2_antennanp ANTENNA_1108 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1109 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1110 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1111 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1112 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1113 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1114 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1115 (.A(_05205_));
 sg13g2_antennanp ANTENNA_1116 (.A(_05209_));
 sg13g2_antennanp ANTENNA_1117 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1118 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1119 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1120 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1121 (.A(_05250_));
 sg13g2_antennanp ANTENNA_1122 (.A(_05250_));
 sg13g2_antennanp ANTENNA_1123 (.A(_05250_));
 sg13g2_antennanp ANTENNA_1124 (.A(_05250_));
 sg13g2_antennanp ANTENNA_1125 (.A(_05252_));
 sg13g2_antennanp ANTENNA_1126 (.A(_05258_));
 sg13g2_antennanp ANTENNA_1127 (.A(_05286_));
 sg13g2_antennanp ANTENNA_1128 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1129 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1130 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1131 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1132 (.A(_05318_));
 sg13g2_antennanp ANTENNA_1133 (.A(_05328_));
 sg13g2_antennanp ANTENNA_1134 (.A(_05339_));
 sg13g2_antennanp ANTENNA_1135 (.A(_05342_));
 sg13g2_antennanp ANTENNA_1136 (.A(_05342_));
 sg13g2_antennanp ANTENNA_1137 (.A(_05342_));
 sg13g2_antennanp ANTENNA_1138 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1139 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1140 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1141 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1142 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1143 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1144 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1145 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1146 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1147 (.A(_05346_));
 sg13g2_antennanp ANTENNA_1148 (.A(_05350_));
 sg13g2_antennanp ANTENNA_1149 (.A(_05389_));
 sg13g2_antennanp ANTENNA_1150 (.A(_05390_));
 sg13g2_antennanp ANTENNA_1151 (.A(_05404_));
 sg13g2_antennanp ANTENNA_1152 (.A(_05415_));
 sg13g2_antennanp ANTENNA_1153 (.A(_05415_));
 sg13g2_antennanp ANTENNA_1154 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1155 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1156 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1157 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1158 (.A(_05442_));
 sg13g2_antennanp ANTENNA_1159 (.A(_05459_));
 sg13g2_antennanp ANTENNA_1160 (.A(_05477_));
 sg13g2_antennanp ANTENNA_1161 (.A(_05500_));
 sg13g2_antennanp ANTENNA_1162 (.A(_05576_));
 sg13g2_antennanp ANTENNA_1163 (.A(_05591_));
 sg13g2_antennanp ANTENNA_1164 (.A(_05591_));
 sg13g2_antennanp ANTENNA_1165 (.A(_05591_));
 sg13g2_antennanp ANTENNA_1166 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1167 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1168 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1169 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1170 (.A(_05611_));
 sg13g2_antennanp ANTENNA_1171 (.A(_05633_));
 sg13g2_antennanp ANTENNA_1172 (.A(_05681_));
 sg13g2_antennanp ANTENNA_1173 (.A(_05726_));
 sg13g2_antennanp ANTENNA_1174 (.A(_05750_));
 sg13g2_antennanp ANTENNA_1175 (.A(_05777_));
 sg13g2_antennanp ANTENNA_1176 (.A(_05814_));
 sg13g2_antennanp ANTENNA_1177 (.A(_05816_));
 sg13g2_antennanp ANTENNA_1178 (.A(_05818_));
 sg13g2_antennanp ANTENNA_1179 (.A(_05827_));
 sg13g2_antennanp ANTENNA_1180 (.A(_05829_));
 sg13g2_antennanp ANTENNA_1181 (.A(_05837_));
 sg13g2_antennanp ANTENNA_1182 (.A(_05874_));
 sg13g2_antennanp ANTENNA_1183 (.A(_05886_));
 sg13g2_antennanp ANTENNA_1184 (.A(_05886_));
 sg13g2_antennanp ANTENNA_1185 (.A(_05890_));
 sg13g2_antennanp ANTENNA_1186 (.A(_05897_));
 sg13g2_antennanp ANTENNA_1187 (.A(_05904_));
 sg13g2_antennanp ANTENNA_1188 (.A(_05924_));
 sg13g2_antennanp ANTENNA_1189 (.A(_05924_));
 sg13g2_antennanp ANTENNA_1190 (.A(_05939_));
 sg13g2_antennanp ANTENNA_1191 (.A(_05946_));
 sg13g2_antennanp ANTENNA_1192 (.A(_05951_));
 sg13g2_antennanp ANTENNA_1193 (.A(_05957_));
 sg13g2_antennanp ANTENNA_1194 (.A(_05998_));
 sg13g2_antennanp ANTENNA_1195 (.A(_06018_));
 sg13g2_antennanp ANTENNA_1196 (.A(_06023_));
 sg13g2_antennanp ANTENNA_1197 (.A(_06046_));
 sg13g2_antennanp ANTENNA_1198 (.A(_06050_));
 sg13g2_antennanp ANTENNA_1199 (.A(_06053_));
 sg13g2_antennanp ANTENNA_1200 (.A(_06064_));
 sg13g2_antennanp ANTENNA_1201 (.A(_06075_));
 sg13g2_antennanp ANTENNA_1202 (.A(_06091_));
 sg13g2_antennanp ANTENNA_1203 (.A(_06116_));
 sg13g2_antennanp ANTENNA_1204 (.A(_06134_));
 sg13g2_antennanp ANTENNA_1205 (.A(_06134_));
 sg13g2_antennanp ANTENNA_1206 (.A(_06139_));
 sg13g2_antennanp ANTENNA_1207 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1208 (.A(_06151_));
 sg13g2_antennanp ANTENNA_1209 (.A(_06167_));
 sg13g2_antennanp ANTENNA_1210 (.A(_06179_));
 sg13g2_antennanp ANTENNA_1211 (.A(_06182_));
 sg13g2_antennanp ANTENNA_1212 (.A(_06182_));
 sg13g2_antennanp ANTENNA_1213 (.A(_06196_));
 sg13g2_antennanp ANTENNA_1214 (.A(_06209_));
 sg13g2_antennanp ANTENNA_1215 (.A(_06225_));
 sg13g2_antennanp ANTENNA_1216 (.A(_06227_));
 sg13g2_antennanp ANTENNA_1217 (.A(_06244_));
 sg13g2_antennanp ANTENNA_1218 (.A(_06249_));
 sg13g2_antennanp ANTENNA_1219 (.A(_06250_));
 sg13g2_antennanp ANTENNA_1220 (.A(_06271_));
 sg13g2_antennanp ANTENNA_1221 (.A(_06271_));
 sg13g2_antennanp ANTENNA_1222 (.A(_06281_));
 sg13g2_antennanp ANTENNA_1223 (.A(_06290_));
 sg13g2_antennanp ANTENNA_1224 (.A(_06300_));
 sg13g2_antennanp ANTENNA_1225 (.A(_06322_));
 sg13g2_antennanp ANTENNA_1226 (.A(_06324_));
 sg13g2_antennanp ANTENNA_1227 (.A(_06328_));
 sg13g2_antennanp ANTENNA_1228 (.A(_06334_));
 sg13g2_antennanp ANTENNA_1229 (.A(_06335_));
 sg13g2_antennanp ANTENNA_1230 (.A(_06342_));
 sg13g2_antennanp ANTENNA_1231 (.A(_06347_));
 sg13g2_antennanp ANTENNA_1232 (.A(_06351_));
 sg13g2_antennanp ANTENNA_1233 (.A(_06361_));
 sg13g2_antennanp ANTENNA_1234 (.A(_06366_));
 sg13g2_antennanp ANTENNA_1235 (.A(_06372_));
 sg13g2_antennanp ANTENNA_1236 (.A(_06374_));
 sg13g2_antennanp ANTENNA_1237 (.A(_06391_));
 sg13g2_antennanp ANTENNA_1238 (.A(_06396_));
 sg13g2_antennanp ANTENNA_1239 (.A(_06397_));
 sg13g2_antennanp ANTENNA_1240 (.A(_06417_));
 sg13g2_antennanp ANTENNA_1241 (.A(_06417_));
 sg13g2_antennanp ANTENNA_1242 (.A(_06422_));
 sg13g2_antennanp ANTENNA_1243 (.A(_06440_));
 sg13g2_antennanp ANTENNA_1244 (.A(_06448_));
 sg13g2_antennanp ANTENNA_1245 (.A(_06467_));
 sg13g2_antennanp ANTENNA_1246 (.A(_06484_));
 sg13g2_antennanp ANTENNA_1247 (.A(_06492_));
 sg13g2_antennanp ANTENNA_1248 (.A(_06497_));
 sg13g2_antennanp ANTENNA_1249 (.A(_06504_));
 sg13g2_antennanp ANTENNA_1250 (.A(_06506_));
 sg13g2_antennanp ANTENNA_1251 (.A(_06512_));
 sg13g2_antennanp ANTENNA_1252 (.A(_06517_));
 sg13g2_antennanp ANTENNA_1253 (.A(_06522_));
 sg13g2_antennanp ANTENNA_1254 (.A(_06523_));
 sg13g2_antennanp ANTENNA_1255 (.A(_06546_));
 sg13g2_antennanp ANTENNA_1256 (.A(_06548_));
 sg13g2_antennanp ANTENNA_1257 (.A(_06559_));
 sg13g2_antennanp ANTENNA_1258 (.A(_06588_));
 sg13g2_antennanp ANTENNA_1259 (.A(_06589_));
 sg13g2_antennanp ANTENNA_1260 (.A(_06596_));
 sg13g2_antennanp ANTENNA_1261 (.A(_06621_));
 sg13g2_antennanp ANTENNA_1262 (.A(_06640_));
 sg13g2_antennanp ANTENNA_1263 (.A(_06658_));
 sg13g2_antennanp ANTENNA_1264 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1265 (.A(_06679_));
 sg13g2_antennanp ANTENNA_1266 (.A(_06680_));
 sg13g2_antennanp ANTENNA_1267 (.A(_06682_));
 sg13g2_antennanp ANTENNA_1268 (.A(_06684_));
 sg13g2_antennanp ANTENNA_1269 (.A(_06687_));
 sg13g2_antennanp ANTENNA_1270 (.A(_06688_));
 sg13g2_antennanp ANTENNA_1271 (.A(_06701_));
 sg13g2_antennanp ANTENNA_1272 (.A(_06712_));
 sg13g2_antennanp ANTENNA_1273 (.A(_06732_));
 sg13g2_antennanp ANTENNA_1274 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1275 (.A(_06758_));
 sg13g2_antennanp ANTENNA_1276 (.A(_06761_));
 sg13g2_antennanp ANTENNA_1277 (.A(_06761_));
 sg13g2_antennanp ANTENNA_1278 (.A(_06764_));
 sg13g2_antennanp ANTENNA_1279 (.A(_06768_));
 sg13g2_antennanp ANTENNA_1280 (.A(_06775_));
 sg13g2_antennanp ANTENNA_1281 (.A(_06796_));
 sg13g2_antennanp ANTENNA_1282 (.A(_06813_));
 sg13g2_antennanp ANTENNA_1283 (.A(_06830_));
 sg13g2_antennanp ANTENNA_1284 (.A(_06830_));
 sg13g2_antennanp ANTENNA_1285 (.A(_06834_));
 sg13g2_antennanp ANTENNA_1286 (.A(_06849_));
 sg13g2_antennanp ANTENNA_1287 (.A(_06905_));
 sg13g2_antennanp ANTENNA_1288 (.A(_06905_));
 sg13g2_antennanp ANTENNA_1289 (.A(_06905_));
 sg13g2_antennanp ANTENNA_1290 (.A(_06926_));
 sg13g2_antennanp ANTENNA_1291 (.A(_07022_));
 sg13g2_antennanp ANTENNA_1292 (.A(_07040_));
 sg13g2_antennanp ANTENNA_1293 (.A(_07040_));
 sg13g2_antennanp ANTENNA_1294 (.A(_07057_));
 sg13g2_antennanp ANTENNA_1295 (.A(_07071_));
 sg13g2_antennanp ANTENNA_1296 (.A(_07071_));
 sg13g2_antennanp ANTENNA_1297 (.A(_07085_));
 sg13g2_antennanp ANTENNA_1298 (.A(_07098_));
 sg13g2_antennanp ANTENNA_1299 (.A(_07154_));
 sg13g2_antennanp ANTENNA_1300 (.A(_07170_));
 sg13g2_antennanp ANTENNA_1301 (.A(_07243_));
 sg13g2_antennanp ANTENNA_1302 (.A(_07258_));
 sg13g2_antennanp ANTENNA_1303 (.A(_07273_));
 sg13g2_antennanp ANTENNA_1304 (.A(_07316_));
 sg13g2_antennanp ANTENNA_1305 (.A(_07316_));
 sg13g2_antennanp ANTENNA_1306 (.A(_07331_));
 sg13g2_antennanp ANTENNA_1307 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1308 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1309 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1310 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1311 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1312 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1313 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1314 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1315 (.A(_07534_));
 sg13g2_antennanp ANTENNA_1316 (.A(_07663_));
 sg13g2_antennanp ANTENNA_1317 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1318 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1319 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1320 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1321 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1322 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1323 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1324 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1325 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1326 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1327 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1328 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1329 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1330 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1331 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1332 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1333 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1334 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1335 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1336 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1337 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1338 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1339 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1340 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1341 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1342 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1343 (.A(_09301_));
 sg13g2_antennanp ANTENNA_1344 (.A(_09301_));
 sg13g2_antennanp ANTENNA_1345 (.A(_09301_));
 sg13g2_antennanp ANTENNA_1346 (.A(_09301_));
 sg13g2_antennanp ANTENNA_1347 (.A(_09301_));
 sg13g2_antennanp ANTENNA_1348 (.A(_09301_));
 sg13g2_antennanp ANTENNA_1349 (.A(_09573_));
 sg13g2_antennanp ANTENNA_1350 (.A(_09573_));
 sg13g2_antennanp ANTENNA_1351 (.A(_09573_));
 sg13g2_antennanp ANTENNA_1352 (.A(_09573_));
 sg13g2_antennanp ANTENNA_1353 (.A(_09599_));
 sg13g2_antennanp ANTENNA_1354 (.A(_09599_));
 sg13g2_antennanp ANTENNA_1355 (.A(_09599_));
 sg13g2_antennanp ANTENNA_1356 (.A(_09599_));
 sg13g2_antennanp ANTENNA_1357 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1358 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1359 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1360 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1361 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1362 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1363 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1364 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1365 (.A(_09910_));
 sg13g2_antennanp ANTENNA_1366 (.A(_09960_));
 sg13g2_antennanp ANTENNA_1367 (.A(_09960_));
 sg13g2_antennanp ANTENNA_1368 (.A(_09960_));
 sg13g2_antennanp ANTENNA_1369 (.A(_09960_));
 sg13g2_antennanp ANTENNA_1370 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1371 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1372 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1373 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1374 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1375 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1376 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1377 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1378 (.A(_10009_));
 sg13g2_antennanp ANTENNA_1379 (.A(_10032_));
 sg13g2_antennanp ANTENNA_1380 (.A(_10032_));
 sg13g2_antennanp ANTENNA_1381 (.A(_10032_));
 sg13g2_antennanp ANTENNA_1382 (.A(_10032_));
 sg13g2_antennanp ANTENNA_1383 (.A(_10074_));
 sg13g2_antennanp ANTENNA_1384 (.A(_10074_));
 sg13g2_antennanp ANTENNA_1385 (.A(_10074_));
 sg13g2_antennanp ANTENNA_1386 (.A(_10074_));
 sg13g2_antennanp ANTENNA_1387 (.A(_10077_));
 sg13g2_antennanp ANTENNA_1388 (.A(_10077_));
 sg13g2_antennanp ANTENNA_1389 (.A(_10077_));
 sg13g2_antennanp ANTENNA_1390 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1391 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1392 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1393 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1394 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1395 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1396 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1397 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1398 (.A(_10085_));
 sg13g2_antennanp ANTENNA_1399 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1400 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1401 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1402 (.A(_10092_));
 sg13g2_antennanp ANTENNA_1403 (.A(_10151_));
 sg13g2_antennanp ANTENNA_1404 (.A(_10151_));
 sg13g2_antennanp ANTENNA_1405 (.A(_10151_));
 sg13g2_antennanp ANTENNA_1406 (.A(_10151_));
 sg13g2_antennanp ANTENNA_1407 (.A(_10151_));
 sg13g2_antennanp ANTENNA_1408 (.A(_10151_));
 sg13g2_antennanp ANTENNA_1409 (.A(_10404_));
 sg13g2_antennanp ANTENNA_1410 (.A(_10404_));
 sg13g2_antennanp ANTENNA_1411 (.A(_10404_));
 sg13g2_antennanp ANTENNA_1412 (.A(_10404_));
 sg13g2_antennanp ANTENNA_1413 (.A(_10435_));
 sg13g2_antennanp ANTENNA_1414 (.A(_10435_));
 sg13g2_antennanp ANTENNA_1415 (.A(_10435_));
 sg13g2_antennanp ANTENNA_1416 (.A(_10435_));
 sg13g2_antennanp ANTENNA_1417 (.A(_10460_));
 sg13g2_antennanp ANTENNA_1418 (.A(_10460_));
 sg13g2_antennanp ANTENNA_1419 (.A(_10460_));
 sg13g2_antennanp ANTENNA_1420 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_1421 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_1422 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_1423 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_1424 (.A(\top_ihp.oisc.regs[2][4] ));
 sg13g2_antennanp ANTENNA_1425 (.A(\top_ihp.oisc.regs[2][4] ));
 sg13g2_antennanp ANTENNA_1426 (.A(\top_ihp.oisc.regs[2][4] ));
 sg13g2_antennanp ANTENNA_1427 (.A(\top_ihp.oisc.regs[2][4] ));
 sg13g2_antennanp ANTENNA_1428 (.A(\top_ihp.oisc.regs[2][4] ));
 sg13g2_antennanp ANTENNA_1429 (.A(\top_ihp.oisc.regs[2][4] ));
 sg13g2_antennanp ANTENNA_1430 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1431 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1432 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1433 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_1434 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_1435 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_1436 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_1437 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_1438 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1439 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1440 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1441 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1442 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1443 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1444 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1445 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1446 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1447 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1448 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1449 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1450 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1451 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_1452 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_1453 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_1454 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_1455 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_1456 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_1457 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_1458 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1459 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1460 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1461 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1462 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1463 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1464 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1465 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1466 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1467 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1468 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1469 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1470 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1471 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1472 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_1473 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_1474 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_1475 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_1476 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_1477 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_1478 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_1479 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_1480 (.A(\top_ihp.ram_cs_o ));
 sg13g2_antennanp ANTENNA_1481 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_1482 (.A(net1));
 sg13g2_antennanp ANTENNA_1483 (.A(net1));
 sg13g2_antennanp ANTENNA_1484 (.A(net1));
 sg13g2_antennanp ANTENNA_1485 (.A(net9));
 sg13g2_antennanp ANTENNA_1486 (.A(net47));
 sg13g2_antennanp ANTENNA_1487 (.A(net47));
 sg13g2_antennanp ANTENNA_1488 (.A(net47));
 sg13g2_antennanp ANTENNA_1489 (.A(net47));
 sg13g2_antennanp ANTENNA_1490 (.A(net47));
 sg13g2_antennanp ANTENNA_1491 (.A(net47));
 sg13g2_antennanp ANTENNA_1492 (.A(net47));
 sg13g2_antennanp ANTENNA_1493 (.A(net47));
 sg13g2_antennanp ANTENNA_1494 (.A(net47));
 sg13g2_antennanp ANTENNA_1495 (.A(net87));
 sg13g2_antennanp ANTENNA_1496 (.A(net87));
 sg13g2_antennanp ANTENNA_1497 (.A(net87));
 sg13g2_antennanp ANTENNA_1498 (.A(net87));
 sg13g2_antennanp ANTENNA_1499 (.A(net87));
 sg13g2_antennanp ANTENNA_1500 (.A(net87));
 sg13g2_antennanp ANTENNA_1501 (.A(net87));
 sg13g2_antennanp ANTENNA_1502 (.A(net87));
 sg13g2_antennanp ANTENNA_1503 (.A(net87));
 sg13g2_antennanp ANTENNA_1504 (.A(net136));
 sg13g2_antennanp ANTENNA_1505 (.A(net136));
 sg13g2_antennanp ANTENNA_1506 (.A(net136));
 sg13g2_antennanp ANTENNA_1507 (.A(net136));
 sg13g2_antennanp ANTENNA_1508 (.A(net136));
 sg13g2_antennanp ANTENNA_1509 (.A(net136));
 sg13g2_antennanp ANTENNA_1510 (.A(net136));
 sg13g2_antennanp ANTENNA_1511 (.A(net136));
 sg13g2_antennanp ANTENNA_1512 (.A(net136));
 sg13g2_antennanp ANTENNA_1513 (.A(net142));
 sg13g2_antennanp ANTENNA_1514 (.A(net142));
 sg13g2_antennanp ANTENNA_1515 (.A(net142));
 sg13g2_antennanp ANTENNA_1516 (.A(net142));
 sg13g2_antennanp ANTENNA_1517 (.A(net142));
 sg13g2_antennanp ANTENNA_1518 (.A(net142));
 sg13g2_antennanp ANTENNA_1519 (.A(net142));
 sg13g2_antennanp ANTENNA_1520 (.A(net142));
 sg13g2_antennanp ANTENNA_1521 (.A(net142));
 sg13g2_antennanp ANTENNA_1522 (.A(net235));
 sg13g2_antennanp ANTENNA_1523 (.A(net235));
 sg13g2_antennanp ANTENNA_1524 (.A(net235));
 sg13g2_antennanp ANTENNA_1525 (.A(net235));
 sg13g2_antennanp ANTENNA_1526 (.A(net235));
 sg13g2_antennanp ANTENNA_1527 (.A(net235));
 sg13g2_antennanp ANTENNA_1528 (.A(net235));
 sg13g2_antennanp ANTENNA_1529 (.A(net235));
 sg13g2_antennanp ANTENNA_1530 (.A(net235));
 sg13g2_antennanp ANTENNA_1531 (.A(net255));
 sg13g2_antennanp ANTENNA_1532 (.A(net255));
 sg13g2_antennanp ANTENNA_1533 (.A(net255));
 sg13g2_antennanp ANTENNA_1534 (.A(net255));
 sg13g2_antennanp ANTENNA_1535 (.A(net255));
 sg13g2_antennanp ANTENNA_1536 (.A(net255));
 sg13g2_antennanp ANTENNA_1537 (.A(net255));
 sg13g2_antennanp ANTENNA_1538 (.A(net255));
 sg13g2_antennanp ANTENNA_1539 (.A(net334));
 sg13g2_antennanp ANTENNA_1540 (.A(net334));
 sg13g2_antennanp ANTENNA_1541 (.A(net334));
 sg13g2_antennanp ANTENNA_1542 (.A(net334));
 sg13g2_antennanp ANTENNA_1543 (.A(net334));
 sg13g2_antennanp ANTENNA_1544 (.A(net334));
 sg13g2_antennanp ANTENNA_1545 (.A(net334));
 sg13g2_antennanp ANTENNA_1546 (.A(net334));
 sg13g2_antennanp ANTENNA_1547 (.A(net347));
 sg13g2_antennanp ANTENNA_1548 (.A(net347));
 sg13g2_antennanp ANTENNA_1549 (.A(net347));
 sg13g2_antennanp ANTENNA_1550 (.A(net347));
 sg13g2_antennanp ANTENNA_1551 (.A(net347));
 sg13g2_antennanp ANTENNA_1552 (.A(net347));
 sg13g2_antennanp ANTENNA_1553 (.A(net347));
 sg13g2_antennanp ANTENNA_1554 (.A(net347));
 sg13g2_antennanp ANTENNA_1555 (.A(net348));
 sg13g2_antennanp ANTENNA_1556 (.A(net348));
 sg13g2_antennanp ANTENNA_1557 (.A(net348));
 sg13g2_antennanp ANTENNA_1558 (.A(net348));
 sg13g2_antennanp ANTENNA_1559 (.A(net348));
 sg13g2_antennanp ANTENNA_1560 (.A(net348));
 sg13g2_antennanp ANTENNA_1561 (.A(net348));
 sg13g2_antennanp ANTENNA_1562 (.A(net348));
 sg13g2_antennanp ANTENNA_1563 (.A(net412));
 sg13g2_antennanp ANTENNA_1564 (.A(net412));
 sg13g2_antennanp ANTENNA_1565 (.A(net412));
 sg13g2_antennanp ANTENNA_1566 (.A(net412));
 sg13g2_antennanp ANTENNA_1567 (.A(net412));
 sg13g2_antennanp ANTENNA_1568 (.A(net412));
 sg13g2_antennanp ANTENNA_1569 (.A(net412));
 sg13g2_antennanp ANTENNA_1570 (.A(net412));
 sg13g2_antennanp ANTENNA_1571 (.A(net412));
 sg13g2_antennanp ANTENNA_1572 (.A(net413));
 sg13g2_antennanp ANTENNA_1573 (.A(net413));
 sg13g2_antennanp ANTENNA_1574 (.A(net413));
 sg13g2_antennanp ANTENNA_1575 (.A(net413));
 sg13g2_antennanp ANTENNA_1576 (.A(net413));
 sg13g2_antennanp ANTENNA_1577 (.A(net413));
 sg13g2_antennanp ANTENNA_1578 (.A(net413));
 sg13g2_antennanp ANTENNA_1579 (.A(net413));
 sg13g2_antennanp ANTENNA_1580 (.A(net413));
 sg13g2_antennanp ANTENNA_1581 (.A(net413));
 sg13g2_antennanp ANTENNA_1582 (.A(net413));
 sg13g2_antennanp ANTENNA_1583 (.A(net413));
 sg13g2_antennanp ANTENNA_1584 (.A(net413));
 sg13g2_antennanp ANTENNA_1585 (.A(net413));
 sg13g2_antennanp ANTENNA_1586 (.A(net413));
 sg13g2_antennanp ANTENNA_1587 (.A(net413));
 sg13g2_antennanp ANTENNA_1588 (.A(net413));
 sg13g2_antennanp ANTENNA_1589 (.A(net413));
 sg13g2_antennanp ANTENNA_1590 (.A(net413));
 sg13g2_antennanp ANTENNA_1591 (.A(net413));
 sg13g2_antennanp ANTENNA_1592 (.A(net413));
 sg13g2_antennanp ANTENNA_1593 (.A(net413));
 sg13g2_antennanp ANTENNA_1594 (.A(net413));
 sg13g2_antennanp ANTENNA_1595 (.A(net413));
 sg13g2_antennanp ANTENNA_1596 (.A(net413));
 sg13g2_antennanp ANTENNA_1597 (.A(net413));
 sg13g2_antennanp ANTENNA_1598 (.A(net413));
 sg13g2_antennanp ANTENNA_1599 (.A(net413));
 sg13g2_antennanp ANTENNA_1600 (.A(net413));
 sg13g2_antennanp ANTENNA_1601 (.A(net413));
 sg13g2_antennanp ANTENNA_1602 (.A(net420));
 sg13g2_antennanp ANTENNA_1603 (.A(net420));
 sg13g2_antennanp ANTENNA_1604 (.A(net420));
 sg13g2_antennanp ANTENNA_1605 (.A(net420));
 sg13g2_antennanp ANTENNA_1606 (.A(net420));
 sg13g2_antennanp ANTENNA_1607 (.A(net420));
 sg13g2_antennanp ANTENNA_1608 (.A(net420));
 sg13g2_antennanp ANTENNA_1609 (.A(net420));
 sg13g2_antennanp ANTENNA_1610 (.A(net454));
 sg13g2_antennanp ANTENNA_1611 (.A(net454));
 sg13g2_antennanp ANTENNA_1612 (.A(net454));
 sg13g2_antennanp ANTENNA_1613 (.A(net454));
 sg13g2_antennanp ANTENNA_1614 (.A(net454));
 sg13g2_antennanp ANTENNA_1615 (.A(net454));
 sg13g2_antennanp ANTENNA_1616 (.A(net454));
 sg13g2_antennanp ANTENNA_1617 (.A(net454));
 sg13g2_antennanp ANTENNA_1618 (.A(net454));
 sg13g2_antennanp ANTENNA_1619 (.A(net474));
 sg13g2_antennanp ANTENNA_1620 (.A(net474));
 sg13g2_antennanp ANTENNA_1621 (.A(net474));
 sg13g2_antennanp ANTENNA_1622 (.A(net474));
 sg13g2_antennanp ANTENNA_1623 (.A(net474));
 sg13g2_antennanp ANTENNA_1624 (.A(net474));
 sg13g2_antennanp ANTENNA_1625 (.A(net474));
 sg13g2_antennanp ANTENNA_1626 (.A(net474));
 sg13g2_antennanp ANTENNA_1627 (.A(net474));
 sg13g2_antennanp ANTENNA_1628 (.A(net474));
 sg13g2_antennanp ANTENNA_1629 (.A(net474));
 sg13g2_antennanp ANTENNA_1630 (.A(net474));
 sg13g2_antennanp ANTENNA_1631 (.A(net474));
 sg13g2_antennanp ANTENNA_1632 (.A(net475));
 sg13g2_antennanp ANTENNA_1633 (.A(net475));
 sg13g2_antennanp ANTENNA_1634 (.A(net475));
 sg13g2_antennanp ANTENNA_1635 (.A(net475));
 sg13g2_antennanp ANTENNA_1636 (.A(net475));
 sg13g2_antennanp ANTENNA_1637 (.A(net475));
 sg13g2_antennanp ANTENNA_1638 (.A(net475));
 sg13g2_antennanp ANTENNA_1639 (.A(net475));
 sg13g2_antennanp ANTENNA_1640 (.A(net480));
 sg13g2_antennanp ANTENNA_1641 (.A(net480));
 sg13g2_antennanp ANTENNA_1642 (.A(net480));
 sg13g2_antennanp ANTENNA_1643 (.A(net480));
 sg13g2_antennanp ANTENNA_1644 (.A(net480));
 sg13g2_antennanp ANTENNA_1645 (.A(net480));
 sg13g2_antennanp ANTENNA_1646 (.A(net480));
 sg13g2_antennanp ANTENNA_1647 (.A(net480));
 sg13g2_antennanp ANTENNA_1648 (.A(net480));
 sg13g2_antennanp ANTENNA_1649 (.A(net483));
 sg13g2_antennanp ANTENNA_1650 (.A(net483));
 sg13g2_antennanp ANTENNA_1651 (.A(net483));
 sg13g2_antennanp ANTENNA_1652 (.A(net483));
 sg13g2_antennanp ANTENNA_1653 (.A(net483));
 sg13g2_antennanp ANTENNA_1654 (.A(net483));
 sg13g2_antennanp ANTENNA_1655 (.A(net483));
 sg13g2_antennanp ANTENNA_1656 (.A(net483));
 sg13g2_antennanp ANTENNA_1657 (.A(net483));
 sg13g2_antennanp ANTENNA_1658 (.A(net595));
 sg13g2_antennanp ANTENNA_1659 (.A(net595));
 sg13g2_antennanp ANTENNA_1660 (.A(net595));
 sg13g2_antennanp ANTENNA_1661 (.A(net595));
 sg13g2_antennanp ANTENNA_1662 (.A(net595));
 sg13g2_antennanp ANTENNA_1663 (.A(net595));
 sg13g2_antennanp ANTENNA_1664 (.A(net595));
 sg13g2_antennanp ANTENNA_1665 (.A(net595));
 sg13g2_antennanp ANTENNA_1666 (.A(net595));
 sg13g2_antennanp ANTENNA_1667 (.A(net595));
 sg13g2_antennanp ANTENNA_1668 (.A(net595));
 sg13g2_antennanp ANTENNA_1669 (.A(net595));
 sg13g2_antennanp ANTENNA_1670 (.A(net643));
 sg13g2_antennanp ANTENNA_1671 (.A(net643));
 sg13g2_antennanp ANTENNA_1672 (.A(net643));
 sg13g2_antennanp ANTENNA_1673 (.A(net643));
 sg13g2_antennanp ANTENNA_1674 (.A(net643));
 sg13g2_antennanp ANTENNA_1675 (.A(net643));
 sg13g2_antennanp ANTENNA_1676 (.A(net643));
 sg13g2_antennanp ANTENNA_1677 (.A(net643));
 sg13g2_antennanp ANTENNA_1678 (.A(net643));
 sg13g2_antennanp ANTENNA_1679 (.A(net663));
 sg13g2_antennanp ANTENNA_1680 (.A(net663));
 sg13g2_antennanp ANTENNA_1681 (.A(net663));
 sg13g2_antennanp ANTENNA_1682 (.A(net663));
 sg13g2_antennanp ANTENNA_1683 (.A(net663));
 sg13g2_antennanp ANTENNA_1684 (.A(net663));
 sg13g2_antennanp ANTENNA_1685 (.A(net663));
 sg13g2_antennanp ANTENNA_1686 (.A(net663));
 sg13g2_antennanp ANTENNA_1687 (.A(net663));
 sg13g2_antennanp ANTENNA_1688 (.A(net663));
 sg13g2_antennanp ANTENNA_1689 (.A(net663));
 sg13g2_antennanp ANTENNA_1690 (.A(net663));
 sg13g2_antennanp ANTENNA_1691 (.A(net663));
 sg13g2_antennanp ANTENNA_1692 (.A(net663));
 sg13g2_antennanp ANTENNA_1693 (.A(net663));
 sg13g2_antennanp ANTENNA_1694 (.A(net663));
 sg13g2_antennanp ANTENNA_1695 (.A(net710));
 sg13g2_antennanp ANTENNA_1696 (.A(net710));
 sg13g2_antennanp ANTENNA_1697 (.A(net710));
 sg13g2_antennanp ANTENNA_1698 (.A(net710));
 sg13g2_antennanp ANTENNA_1699 (.A(net710));
 sg13g2_antennanp ANTENNA_1700 (.A(net710));
 sg13g2_antennanp ANTENNA_1701 (.A(net710));
 sg13g2_antennanp ANTENNA_1702 (.A(net710));
 sg13g2_antennanp ANTENNA_1703 (.A(net735));
 sg13g2_antennanp ANTENNA_1704 (.A(net735));
 sg13g2_antennanp ANTENNA_1705 (.A(net735));
 sg13g2_antennanp ANTENNA_1706 (.A(net735));
 sg13g2_antennanp ANTENNA_1707 (.A(net735));
 sg13g2_antennanp ANTENNA_1708 (.A(net735));
 sg13g2_antennanp ANTENNA_1709 (.A(net735));
 sg13g2_antennanp ANTENNA_1710 (.A(net735));
 sg13g2_antennanp ANTENNA_1711 (.A(net735));
 sg13g2_antennanp ANTENNA_1712 (.A(_00294_));
 sg13g2_antennanp ANTENNA_1713 (.A(_00294_));
 sg13g2_antennanp ANTENNA_1714 (.A(_00296_));
 sg13g2_antennanp ANTENNA_1715 (.A(_00299_));
 sg13g2_antennanp ANTENNA_1716 (.A(_00299_));
 sg13g2_antennanp ANTENNA_1717 (.A(_00300_));
 sg13g2_antennanp ANTENNA_1718 (.A(_00305_));
 sg13g2_antennanp ANTENNA_1719 (.A(_00307_));
 sg13g2_antennanp ANTENNA_1720 (.A(_00311_));
 sg13g2_antennanp ANTENNA_1721 (.A(_00311_));
 sg13g2_antennanp ANTENNA_1722 (.A(_00316_));
 sg13g2_antennanp ANTENNA_1723 (.A(_00319_));
 sg13g2_antennanp ANTENNA_1724 (.A(_00320_));
 sg13g2_antennanp ANTENNA_1725 (.A(_00322_));
 sg13g2_antennanp ANTENNA_1726 (.A(_00322_));
 sg13g2_antennanp ANTENNA_1727 (.A(_00324_));
 sg13g2_antennanp ANTENNA_1728 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1729 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1730 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1731 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1732 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1733 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1734 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1735 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1736 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1737 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1738 (.A(_03021_));
 sg13g2_antennanp ANTENNA_1739 (.A(_03021_));
 sg13g2_antennanp ANTENNA_1740 (.A(_03021_));
 sg13g2_antennanp ANTENNA_1741 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1742 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1743 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1744 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1745 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1746 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1747 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1748 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1749 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1750 (.A(_03492_));
 sg13g2_antennanp ANTENNA_1751 (.A(_03713_));
 sg13g2_antennanp ANTENNA_1752 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1753 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1754 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1755 (.A(_04741_));
 sg13g2_antennanp ANTENNA_1756 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1757 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1758 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1759 (.A(_04851_));
 sg13g2_antennanp ANTENNA_1760 (.A(_04857_));
 sg13g2_antennanp ANTENNA_1761 (.A(_04871_));
 sg13g2_antennanp ANTENNA_1762 (.A(_04871_));
 sg13g2_antennanp ANTENNA_1763 (.A(_04871_));
 sg13g2_antennanp ANTENNA_1764 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1765 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1766 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1767 (.A(_04873_));
 sg13g2_antennanp ANTENNA_1768 (.A(_04883_));
 sg13g2_antennanp ANTENNA_1769 (.A(_04912_));
 sg13g2_antennanp ANTENNA_1770 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1771 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1772 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1773 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1774 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1775 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1776 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1777 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1778 (.A(_04917_));
 sg13g2_antennanp ANTENNA_1779 (.A(_04921_));
 sg13g2_antennanp ANTENNA_1780 (.A(_04921_));
 sg13g2_antennanp ANTENNA_1781 (.A(_04921_));
 sg13g2_antennanp ANTENNA_1782 (.A(_04932_));
 sg13g2_antennanp ANTENNA_1783 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1784 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1785 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1786 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1787 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1788 (.A(_05012_));
 sg13g2_antennanp ANTENNA_1789 (.A(_05024_));
 sg13g2_antennanp ANTENNA_1790 (.A(_05072_));
 sg13g2_antennanp ANTENNA_1791 (.A(_05072_));
 sg13g2_antennanp ANTENNA_1792 (.A(_05072_));
 sg13g2_antennanp ANTENNA_1793 (.A(_05100_));
 sg13g2_antennanp ANTENNA_1794 (.A(_05100_));
 sg13g2_antennanp ANTENNA_1795 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1796 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1797 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1798 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1799 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1800 (.A(_05101_));
 sg13g2_antennanp ANTENNA_1801 (.A(_05102_));
 sg13g2_antennanp ANTENNA_1802 (.A(_05102_));
 sg13g2_antennanp ANTENNA_1803 (.A(_05118_));
 sg13g2_antennanp ANTENNA_1804 (.A(_05124_));
 sg13g2_antennanp ANTENNA_1805 (.A(_05128_));
 sg13g2_antennanp ANTENNA_1806 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1807 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1808 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1809 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1810 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1811 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1812 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1813 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1814 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1815 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1816 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1817 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1818 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1819 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1820 (.A(_05130_));
 sg13g2_antennanp ANTENNA_1821 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1822 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1823 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1824 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1825 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1826 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1827 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1828 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1829 (.A(_05134_));
 sg13g2_antennanp ANTENNA_1830 (.A(_05136_));
 sg13g2_antennanp ANTENNA_1831 (.A(_05198_));
 sg13g2_antennanp ANTENNA_1832 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1833 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1834 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1835 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1836 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1837 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1838 (.A(_05205_));
 sg13g2_antennanp ANTENNA_1839 (.A(_05209_));
 sg13g2_antennanp ANTENNA_1840 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1841 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1842 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1843 (.A(_05238_));
 sg13g2_antennanp ANTENNA_1844 (.A(_05252_));
 sg13g2_antennanp ANTENNA_1845 (.A(_05258_));
 sg13g2_antennanp ANTENNA_1846 (.A(_05286_));
 sg13g2_antennanp ANTENNA_1847 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1848 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1849 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1850 (.A(_05302_));
 sg13g2_antennanp ANTENNA_1851 (.A(_05318_));
 sg13g2_antennanp ANTENNA_1852 (.A(_05328_));
 sg13g2_antennanp ANTENNA_1853 (.A(_05339_));
 sg13g2_antennanp ANTENNA_1854 (.A(_05342_));
 sg13g2_antennanp ANTENNA_1855 (.A(_05342_));
 sg13g2_antennanp ANTENNA_1856 (.A(_05342_));
 sg13g2_antennanp ANTENNA_1857 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1858 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1859 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1860 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1861 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1862 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1863 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1864 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1865 (.A(_05344_));
 sg13g2_antennanp ANTENNA_1866 (.A(_05346_));
 sg13g2_antennanp ANTENNA_1867 (.A(_05350_));
 sg13g2_antennanp ANTENNA_1868 (.A(_05389_));
 sg13g2_antennanp ANTENNA_1869 (.A(_05404_));
 sg13g2_antennanp ANTENNA_1870 (.A(_05415_));
 sg13g2_antennanp ANTENNA_1871 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1872 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1873 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1874 (.A(_05459_));
 sg13g2_antennanp ANTENNA_1875 (.A(_05477_));
 sg13g2_antennanp ANTENNA_1876 (.A(_05500_));
 sg13g2_antennanp ANTENNA_1877 (.A(_05576_));
 sg13g2_antennanp ANTENNA_1878 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1879 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1880 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1881 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1882 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1883 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1884 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1885 (.A(_05609_));
 sg13g2_antennanp ANTENNA_1886 (.A(_05611_));
 sg13g2_antennanp ANTENNA_1887 (.A(_05633_));
 sg13g2_antennanp ANTENNA_1888 (.A(_05681_));
 sg13g2_antennanp ANTENNA_1889 (.A(_05726_));
 sg13g2_antennanp ANTENNA_1890 (.A(_05750_));
 sg13g2_antennanp ANTENNA_1891 (.A(_05777_));
 sg13g2_antennanp ANTENNA_1892 (.A(_05814_));
 sg13g2_antennanp ANTENNA_1893 (.A(_05816_));
 sg13g2_antennanp ANTENNA_1894 (.A(_05818_));
 sg13g2_antennanp ANTENNA_1895 (.A(_05827_));
 sg13g2_antennanp ANTENNA_1896 (.A(_05829_));
 sg13g2_antennanp ANTENNA_1897 (.A(_05874_));
 sg13g2_antennanp ANTENNA_1898 (.A(_05886_));
 sg13g2_antennanp ANTENNA_1899 (.A(_05890_));
 sg13g2_antennanp ANTENNA_1900 (.A(_05904_));
 sg13g2_antennanp ANTENNA_1901 (.A(_05924_));
 sg13g2_antennanp ANTENNA_1902 (.A(_05924_));
 sg13g2_antennanp ANTENNA_1903 (.A(_05939_));
 sg13g2_antennanp ANTENNA_1904 (.A(_05946_));
 sg13g2_antennanp ANTENNA_1905 (.A(_05951_));
 sg13g2_antennanp ANTENNA_1906 (.A(_05957_));
 sg13g2_antennanp ANTENNA_1907 (.A(_05998_));
 sg13g2_antennanp ANTENNA_1908 (.A(_05998_));
 sg13g2_antennanp ANTENNA_1909 (.A(_06018_));
 sg13g2_antennanp ANTENNA_1910 (.A(_06023_));
 sg13g2_antennanp ANTENNA_1911 (.A(_06046_));
 sg13g2_antennanp ANTENNA_1912 (.A(_06050_));
 sg13g2_antennanp ANTENNA_1913 (.A(_06053_));
 sg13g2_antennanp ANTENNA_1914 (.A(_06053_));
 sg13g2_antennanp ANTENNA_1915 (.A(_06064_));
 sg13g2_antennanp ANTENNA_1916 (.A(_06075_));
 sg13g2_antennanp ANTENNA_1917 (.A(_06083_));
 sg13g2_antennanp ANTENNA_1918 (.A(_06091_));
 sg13g2_antennanp ANTENNA_1919 (.A(_06116_));
 sg13g2_antennanp ANTENNA_1920 (.A(_06134_));
 sg13g2_antennanp ANTENNA_1921 (.A(_06134_));
 sg13g2_antennanp ANTENNA_1922 (.A(_06139_));
 sg13g2_antennanp ANTENNA_1923 (.A(_06146_));
 sg13g2_antennanp ANTENNA_1924 (.A(_06151_));
 sg13g2_antennanp ANTENNA_1925 (.A(_06167_));
 sg13g2_antennanp ANTENNA_1926 (.A(_06179_));
 sg13g2_antennanp ANTENNA_1927 (.A(_06196_));
 sg13g2_antennanp ANTENNA_1928 (.A(_06209_));
 sg13g2_antennanp ANTENNA_1929 (.A(_06225_));
 sg13g2_antennanp ANTENNA_1930 (.A(_06227_));
 sg13g2_antennanp ANTENNA_1931 (.A(_06244_));
 sg13g2_antennanp ANTENNA_1932 (.A(_06249_));
 sg13g2_antennanp ANTENNA_1933 (.A(_06250_));
 sg13g2_antennanp ANTENNA_1934 (.A(_06271_));
 sg13g2_antennanp ANTENNA_1935 (.A(_06271_));
 sg13g2_antennanp ANTENNA_1936 (.A(_06281_));
 sg13g2_antennanp ANTENNA_1937 (.A(_06290_));
 sg13g2_antennanp ANTENNA_1938 (.A(_06300_));
 sg13g2_antennanp ANTENNA_1939 (.A(_06322_));
 sg13g2_antennanp ANTENNA_1940 (.A(_06324_));
 sg13g2_antennanp ANTENNA_1941 (.A(_06328_));
 sg13g2_antennanp ANTENNA_1942 (.A(_06334_));
 sg13g2_antennanp ANTENNA_1943 (.A(_06342_));
 sg13g2_antennanp ANTENNA_1944 (.A(_06347_));
 sg13g2_antennanp ANTENNA_1945 (.A(_06351_));
 sg13g2_antennanp ANTENNA_1946 (.A(_06361_));
 sg13g2_antennanp ANTENNA_1947 (.A(_06366_));
 sg13g2_antennanp ANTENNA_1948 (.A(_06372_));
 sg13g2_antennanp ANTENNA_1949 (.A(_06374_));
 sg13g2_antennanp ANTENNA_1950 (.A(_06391_));
 sg13g2_antennanp ANTENNA_1951 (.A(_06396_));
 sg13g2_antennanp ANTENNA_1952 (.A(_06397_));
 sg13g2_antennanp ANTENNA_1953 (.A(_06417_));
 sg13g2_antennanp ANTENNA_1954 (.A(_06417_));
 sg13g2_antennanp ANTENNA_1955 (.A(_06422_));
 sg13g2_antennanp ANTENNA_1956 (.A(_06440_));
 sg13g2_antennanp ANTENNA_1957 (.A(_06448_));
 sg13g2_antennanp ANTENNA_1958 (.A(_06463_));
 sg13g2_antennanp ANTENNA_1959 (.A(_06467_));
 sg13g2_antennanp ANTENNA_1960 (.A(_06467_));
 sg13g2_antennanp ANTENNA_1961 (.A(_06484_));
 sg13g2_antennanp ANTENNA_1962 (.A(_06492_));
 sg13g2_antennanp ANTENNA_1963 (.A(_06497_));
 sg13g2_antennanp ANTENNA_1964 (.A(_06504_));
 sg13g2_antennanp ANTENNA_1965 (.A(_06506_));
 sg13g2_antennanp ANTENNA_1966 (.A(_06512_));
 sg13g2_antennanp ANTENNA_1967 (.A(_06517_));
 sg13g2_antennanp ANTENNA_1968 (.A(_06522_));
 sg13g2_antennanp ANTENNA_1969 (.A(_06523_));
 sg13g2_antennanp ANTENNA_1970 (.A(_06546_));
 sg13g2_antennanp ANTENNA_1971 (.A(_06548_));
 sg13g2_antennanp ANTENNA_1972 (.A(_06559_));
 sg13g2_antennanp ANTENNA_1973 (.A(_06588_));
 sg13g2_antennanp ANTENNA_1974 (.A(_06589_));
 sg13g2_antennanp ANTENNA_1975 (.A(_06596_));
 sg13g2_antennanp ANTENNA_1976 (.A(_06621_));
 sg13g2_antennanp ANTENNA_1977 (.A(_06640_));
 sg13g2_antennanp ANTENNA_1978 (.A(_06658_));
 sg13g2_antennanp ANTENNA_1979 (.A(_06667_));
 sg13g2_antennanp ANTENNA_1980 (.A(_06679_));
 sg13g2_antennanp ANTENNA_1981 (.A(_06679_));
 sg13g2_antennanp ANTENNA_1982 (.A(_06680_));
 sg13g2_antennanp ANTENNA_1983 (.A(_06682_));
 sg13g2_antennanp ANTENNA_1984 (.A(_06684_));
 sg13g2_antennanp ANTENNA_1985 (.A(_06687_));
 sg13g2_antennanp ANTENNA_1986 (.A(_06688_));
 sg13g2_antennanp ANTENNA_1987 (.A(_06701_));
 sg13g2_antennanp ANTENNA_1988 (.A(_06712_));
 sg13g2_antennanp ANTENNA_1989 (.A(_06732_));
 sg13g2_antennanp ANTENNA_1990 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1991 (.A(_06758_));
 sg13g2_antennanp ANTENNA_1992 (.A(_06761_));
 sg13g2_antennanp ANTENNA_1993 (.A(_06761_));
 sg13g2_antennanp ANTENNA_1994 (.A(_06764_));
 sg13g2_antennanp ANTENNA_1995 (.A(_06768_));
 sg13g2_antennanp ANTENNA_1996 (.A(_06775_));
 sg13g2_antennanp ANTENNA_1997 (.A(_06813_));
 sg13g2_antennanp ANTENNA_1998 (.A(_06830_));
 sg13g2_antennanp ANTENNA_1999 (.A(_06830_));
 sg13g2_antennanp ANTENNA_2000 (.A(_06834_));
 sg13g2_antennanp ANTENNA_2001 (.A(_06849_));
 sg13g2_antennanp ANTENNA_2002 (.A(_06926_));
 sg13g2_antennanp ANTENNA_2003 (.A(_06926_));
 sg13g2_antennanp ANTENNA_2004 (.A(_07040_));
 sg13g2_antennanp ANTENNA_2005 (.A(_07040_));
 sg13g2_antennanp ANTENNA_2006 (.A(_07057_));
 sg13g2_antennanp ANTENNA_2007 (.A(_07071_));
 sg13g2_antennanp ANTENNA_2008 (.A(_07085_));
 sg13g2_antennanp ANTENNA_2009 (.A(_07098_));
 sg13g2_antennanp ANTENNA_2010 (.A(_07154_));
 sg13g2_antennanp ANTENNA_2011 (.A(_07170_));
 sg13g2_antennanp ANTENNA_2012 (.A(_07243_));
 sg13g2_antennanp ANTENNA_2013 (.A(_07258_));
 sg13g2_antennanp ANTENNA_2014 (.A(_07273_));
 sg13g2_antennanp ANTENNA_2015 (.A(_07301_));
 sg13g2_antennanp ANTENNA_2016 (.A(_07301_));
 sg13g2_antennanp ANTENNA_2017 (.A(_07316_));
 sg13g2_antennanp ANTENNA_2018 (.A(_07331_));
 sg13g2_antennanp ANTENNA_2019 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2020 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2021 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2022 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2023 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2024 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2025 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2026 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2027 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2028 (.A(_07663_));
 sg13g2_antennanp ANTENNA_2029 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2030 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2031 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2032 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2033 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2034 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2035 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2036 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2037 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2038 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2039 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2040 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2041 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2042 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2043 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2044 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2045 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2046 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2047 (.A(_09894_));
 sg13g2_antennanp ANTENNA_2048 (.A(_09894_));
 sg13g2_antennanp ANTENNA_2049 (.A(_09894_));
 sg13g2_antennanp ANTENNA_2050 (.A(_09894_));
 sg13g2_antennanp ANTENNA_2051 (.A(_09894_));
 sg13g2_antennanp ANTENNA_2052 (.A(_09894_));
 sg13g2_antennanp ANTENNA_2053 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2054 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2055 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2056 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2057 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2058 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2059 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2060 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2061 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2062 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2063 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2064 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2065 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2066 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2067 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2068 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2069 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2070 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2071 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2072 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2073 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2074 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2075 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2076 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2077 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2078 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2079 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2080 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2081 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2082 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2083 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2084 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2085 (.A(_10077_));
 sg13g2_antennanp ANTENNA_2086 (.A(_10077_));
 sg13g2_antennanp ANTENNA_2087 (.A(_10077_));
 sg13g2_antennanp ANTENNA_2088 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2089 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2090 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2091 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2092 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2093 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2094 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2095 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2096 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2097 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2098 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2099 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2100 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2101 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2102 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2103 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2104 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2105 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2106 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2107 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2108 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2109 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2110 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2111 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2112 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2113 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2114 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2115 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2116 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2117 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2118 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2119 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2120 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2121 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2122 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2123 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2124 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2125 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2126 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2127 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2128 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2129 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2130 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2131 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2132 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2133 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2134 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2135 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2136 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2137 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2138 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2139 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2140 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_2141 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_2142 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_2143 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_2144 (.A(\top_ihp.oisc.regs[32][3] ));
 sg13g2_antennanp ANTENNA_2145 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2146 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2147 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2148 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2149 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2150 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2151 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2152 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2153 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2154 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2155 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2156 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2157 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2158 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2159 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2160 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_2161 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_2162 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_2163 (.A(\top_ihp.ram_cs_o ));
 sg13g2_antennanp ANTENNA_2164 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_2165 (.A(net1));
 sg13g2_antennanp ANTENNA_2166 (.A(net1));
 sg13g2_antennanp ANTENNA_2167 (.A(net1));
 sg13g2_antennanp ANTENNA_2168 (.A(net9));
 sg13g2_antennanp ANTENNA_2169 (.A(net47));
 sg13g2_antennanp ANTENNA_2170 (.A(net47));
 sg13g2_antennanp ANTENNA_2171 (.A(net47));
 sg13g2_antennanp ANTENNA_2172 (.A(net47));
 sg13g2_antennanp ANTENNA_2173 (.A(net47));
 sg13g2_antennanp ANTENNA_2174 (.A(net47));
 sg13g2_antennanp ANTENNA_2175 (.A(net47));
 sg13g2_antennanp ANTENNA_2176 (.A(net47));
 sg13g2_antennanp ANTENNA_2177 (.A(net47));
 sg13g2_antennanp ANTENNA_2178 (.A(net87));
 sg13g2_antennanp ANTENNA_2179 (.A(net87));
 sg13g2_antennanp ANTENNA_2180 (.A(net87));
 sg13g2_antennanp ANTENNA_2181 (.A(net87));
 sg13g2_antennanp ANTENNA_2182 (.A(net87));
 sg13g2_antennanp ANTENNA_2183 (.A(net87));
 sg13g2_antennanp ANTENNA_2184 (.A(net87));
 sg13g2_antennanp ANTENNA_2185 (.A(net87));
 sg13g2_antennanp ANTENNA_2186 (.A(net87));
 sg13g2_antennanp ANTENNA_2187 (.A(net136));
 sg13g2_antennanp ANTENNA_2188 (.A(net136));
 sg13g2_antennanp ANTENNA_2189 (.A(net136));
 sg13g2_antennanp ANTENNA_2190 (.A(net136));
 sg13g2_antennanp ANTENNA_2191 (.A(net136));
 sg13g2_antennanp ANTENNA_2192 (.A(net136));
 sg13g2_antennanp ANTENNA_2193 (.A(net136));
 sg13g2_antennanp ANTENNA_2194 (.A(net136));
 sg13g2_antennanp ANTENNA_2195 (.A(net136));
 sg13g2_antennanp ANTENNA_2196 (.A(net142));
 sg13g2_antennanp ANTENNA_2197 (.A(net142));
 sg13g2_antennanp ANTENNA_2198 (.A(net142));
 sg13g2_antennanp ANTENNA_2199 (.A(net142));
 sg13g2_antennanp ANTENNA_2200 (.A(net142));
 sg13g2_antennanp ANTENNA_2201 (.A(net142));
 sg13g2_antennanp ANTENNA_2202 (.A(net142));
 sg13g2_antennanp ANTENNA_2203 (.A(net142));
 sg13g2_antennanp ANTENNA_2204 (.A(net142));
 sg13g2_antennanp ANTENNA_2205 (.A(net142));
 sg13g2_antennanp ANTENNA_2206 (.A(net142));
 sg13g2_antennanp ANTENNA_2207 (.A(net142));
 sg13g2_antennanp ANTENNA_2208 (.A(net235));
 sg13g2_antennanp ANTENNA_2209 (.A(net235));
 sg13g2_antennanp ANTENNA_2210 (.A(net235));
 sg13g2_antennanp ANTENNA_2211 (.A(net235));
 sg13g2_antennanp ANTENNA_2212 (.A(net235));
 sg13g2_antennanp ANTENNA_2213 (.A(net235));
 sg13g2_antennanp ANTENNA_2214 (.A(net235));
 sg13g2_antennanp ANTENNA_2215 (.A(net235));
 sg13g2_antennanp ANTENNA_2216 (.A(net235));
 sg13g2_antennanp ANTENNA_2217 (.A(net235));
 sg13g2_antennanp ANTENNA_2218 (.A(net235));
 sg13g2_antennanp ANTENNA_2219 (.A(net235));
 sg13g2_antennanp ANTENNA_2220 (.A(net255));
 sg13g2_antennanp ANTENNA_2221 (.A(net255));
 sg13g2_antennanp ANTENNA_2222 (.A(net255));
 sg13g2_antennanp ANTENNA_2223 (.A(net255));
 sg13g2_antennanp ANTENNA_2224 (.A(net255));
 sg13g2_antennanp ANTENNA_2225 (.A(net255));
 sg13g2_antennanp ANTENNA_2226 (.A(net255));
 sg13g2_antennanp ANTENNA_2227 (.A(net255));
 sg13g2_antennanp ANTENNA_2228 (.A(net255));
 sg13g2_antennanp ANTENNA_2229 (.A(net255));
 sg13g2_antennanp ANTENNA_2230 (.A(net255));
 sg13g2_antennanp ANTENNA_2231 (.A(net255));
 sg13g2_antennanp ANTENNA_2232 (.A(net255));
 sg13g2_antennanp ANTENNA_2233 (.A(net334));
 sg13g2_antennanp ANTENNA_2234 (.A(net334));
 sg13g2_antennanp ANTENNA_2235 (.A(net334));
 sg13g2_antennanp ANTENNA_2236 (.A(net334));
 sg13g2_antennanp ANTENNA_2237 (.A(net334));
 sg13g2_antennanp ANTENNA_2238 (.A(net334));
 sg13g2_antennanp ANTENNA_2239 (.A(net334));
 sg13g2_antennanp ANTENNA_2240 (.A(net334));
 sg13g2_antennanp ANTENNA_2241 (.A(net334));
 sg13g2_antennanp ANTENNA_2242 (.A(net347));
 sg13g2_antennanp ANTENNA_2243 (.A(net347));
 sg13g2_antennanp ANTENNA_2244 (.A(net347));
 sg13g2_antennanp ANTENNA_2245 (.A(net347));
 sg13g2_antennanp ANTENNA_2246 (.A(net347));
 sg13g2_antennanp ANTENNA_2247 (.A(net347));
 sg13g2_antennanp ANTENNA_2248 (.A(net347));
 sg13g2_antennanp ANTENNA_2249 (.A(net347));
 sg13g2_antennanp ANTENNA_2250 (.A(net412));
 sg13g2_antennanp ANTENNA_2251 (.A(net412));
 sg13g2_antennanp ANTENNA_2252 (.A(net412));
 sg13g2_antennanp ANTENNA_2253 (.A(net412));
 sg13g2_antennanp ANTENNA_2254 (.A(net412));
 sg13g2_antennanp ANTENNA_2255 (.A(net412));
 sg13g2_antennanp ANTENNA_2256 (.A(net412));
 sg13g2_antennanp ANTENNA_2257 (.A(net412));
 sg13g2_antennanp ANTENNA_2258 (.A(net413));
 sg13g2_antennanp ANTENNA_2259 (.A(net413));
 sg13g2_antennanp ANTENNA_2260 (.A(net413));
 sg13g2_antennanp ANTENNA_2261 (.A(net413));
 sg13g2_antennanp ANTENNA_2262 (.A(net413));
 sg13g2_antennanp ANTENNA_2263 (.A(net413));
 sg13g2_antennanp ANTENNA_2264 (.A(net413));
 sg13g2_antennanp ANTENNA_2265 (.A(net413));
 sg13g2_antennanp ANTENNA_2266 (.A(net413));
 sg13g2_antennanp ANTENNA_2267 (.A(net420));
 sg13g2_antennanp ANTENNA_2268 (.A(net420));
 sg13g2_antennanp ANTENNA_2269 (.A(net420));
 sg13g2_antennanp ANTENNA_2270 (.A(net420));
 sg13g2_antennanp ANTENNA_2271 (.A(net420));
 sg13g2_antennanp ANTENNA_2272 (.A(net420));
 sg13g2_antennanp ANTENNA_2273 (.A(net420));
 sg13g2_antennanp ANTENNA_2274 (.A(net420));
 sg13g2_antennanp ANTENNA_2275 (.A(net454));
 sg13g2_antennanp ANTENNA_2276 (.A(net454));
 sg13g2_antennanp ANTENNA_2277 (.A(net454));
 sg13g2_antennanp ANTENNA_2278 (.A(net454));
 sg13g2_antennanp ANTENNA_2279 (.A(net454));
 sg13g2_antennanp ANTENNA_2280 (.A(net454));
 sg13g2_antennanp ANTENNA_2281 (.A(net454));
 sg13g2_antennanp ANTENNA_2282 (.A(net454));
 sg13g2_antennanp ANTENNA_2283 (.A(net454));
 sg13g2_antennanp ANTENNA_2284 (.A(net474));
 sg13g2_antennanp ANTENNA_2285 (.A(net474));
 sg13g2_antennanp ANTENNA_2286 (.A(net474));
 sg13g2_antennanp ANTENNA_2287 (.A(net474));
 sg13g2_antennanp ANTENNA_2288 (.A(net474));
 sg13g2_antennanp ANTENNA_2289 (.A(net474));
 sg13g2_antennanp ANTENNA_2290 (.A(net474));
 sg13g2_antennanp ANTENNA_2291 (.A(net474));
 sg13g2_antennanp ANTENNA_2292 (.A(net474));
 sg13g2_antennanp ANTENNA_2293 (.A(net474));
 sg13g2_antennanp ANTENNA_2294 (.A(net474));
 sg13g2_antennanp ANTENNA_2295 (.A(net474));
 sg13g2_antennanp ANTENNA_2296 (.A(net474));
 sg13g2_antennanp ANTENNA_2297 (.A(net480));
 sg13g2_antennanp ANTENNA_2298 (.A(net480));
 sg13g2_antennanp ANTENNA_2299 (.A(net480));
 sg13g2_antennanp ANTENNA_2300 (.A(net480));
 sg13g2_antennanp ANTENNA_2301 (.A(net480));
 sg13g2_antennanp ANTENNA_2302 (.A(net480));
 sg13g2_antennanp ANTENNA_2303 (.A(net480));
 sg13g2_antennanp ANTENNA_2304 (.A(net480));
 sg13g2_antennanp ANTENNA_2305 (.A(net480));
 sg13g2_antennanp ANTENNA_2306 (.A(net595));
 sg13g2_antennanp ANTENNA_2307 (.A(net595));
 sg13g2_antennanp ANTENNA_2308 (.A(net595));
 sg13g2_antennanp ANTENNA_2309 (.A(net595));
 sg13g2_antennanp ANTENNA_2310 (.A(net595));
 sg13g2_antennanp ANTENNA_2311 (.A(net595));
 sg13g2_antennanp ANTENNA_2312 (.A(net595));
 sg13g2_antennanp ANTENNA_2313 (.A(net595));
 sg13g2_antennanp ANTENNA_2314 (.A(net595));
 sg13g2_antennanp ANTENNA_2315 (.A(net663));
 sg13g2_antennanp ANTENNA_2316 (.A(net663));
 sg13g2_antennanp ANTENNA_2317 (.A(net663));
 sg13g2_antennanp ANTENNA_2318 (.A(net663));
 sg13g2_antennanp ANTENNA_2319 (.A(net663));
 sg13g2_antennanp ANTENNA_2320 (.A(net663));
 sg13g2_antennanp ANTENNA_2321 (.A(net663));
 sg13g2_antennanp ANTENNA_2322 (.A(net663));
 sg13g2_antennanp ANTENNA_2323 (.A(net663));
 sg13g2_antennanp ANTENNA_2324 (.A(net735));
 sg13g2_antennanp ANTENNA_2325 (.A(net735));
 sg13g2_antennanp ANTENNA_2326 (.A(net735));
 sg13g2_antennanp ANTENNA_2327 (.A(net735));
 sg13g2_antennanp ANTENNA_2328 (.A(net735));
 sg13g2_antennanp ANTENNA_2329 (.A(net735));
 sg13g2_antennanp ANTENNA_2330 (.A(net735));
 sg13g2_antennanp ANTENNA_2331 (.A(net735));
 sg13g2_antennanp ANTENNA_2332 (.A(net735));
 sg13g2_antennanp ANTENNA_2333 (.A(_00294_));
 sg13g2_antennanp ANTENNA_2334 (.A(_00294_));
 sg13g2_antennanp ANTENNA_2335 (.A(_00296_));
 sg13g2_antennanp ANTENNA_2336 (.A(_00299_));
 sg13g2_antennanp ANTENNA_2337 (.A(_00300_));
 sg13g2_antennanp ANTENNA_2338 (.A(_00305_));
 sg13g2_antennanp ANTENNA_2339 (.A(_00307_));
 sg13g2_antennanp ANTENNA_2340 (.A(_00307_));
 sg13g2_antennanp ANTENNA_2341 (.A(_00311_));
 sg13g2_antennanp ANTENNA_2342 (.A(_00311_));
 sg13g2_antennanp ANTENNA_2343 (.A(_00316_));
 sg13g2_antennanp ANTENNA_2344 (.A(_00319_));
 sg13g2_antennanp ANTENNA_2345 (.A(_00320_));
 sg13g2_antennanp ANTENNA_2346 (.A(_00322_));
 sg13g2_antennanp ANTENNA_2347 (.A(_00322_));
 sg13g2_antennanp ANTENNA_2348 (.A(_00324_));
 sg13g2_antennanp ANTENNA_2349 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2350 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2351 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2352 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2353 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2354 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2355 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2356 (.A(_03021_));
 sg13g2_antennanp ANTENNA_2357 (.A(_03021_));
 sg13g2_antennanp ANTENNA_2358 (.A(_03021_));
 sg13g2_antennanp ANTENNA_2359 (.A(_03492_));
 sg13g2_antennanp ANTENNA_2360 (.A(_03492_));
 sg13g2_antennanp ANTENNA_2361 (.A(_03492_));
 sg13g2_antennanp ANTENNA_2362 (.A(_03492_));
 sg13g2_antennanp ANTENNA_2363 (.A(_03713_));
 sg13g2_antennanp ANTENNA_2364 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2365 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2366 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2367 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2368 (.A(_04847_));
 sg13g2_antennanp ANTENNA_2369 (.A(_04847_));
 sg13g2_antennanp ANTENNA_2370 (.A(_04847_));
 sg13g2_antennanp ANTENNA_2371 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2372 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2373 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2374 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2375 (.A(_04857_));
 sg13g2_antennanp ANTENNA_2376 (.A(_04871_));
 sg13g2_antennanp ANTENNA_2377 (.A(_04871_));
 sg13g2_antennanp ANTENNA_2378 (.A(_04871_));
 sg13g2_antennanp ANTENNA_2379 (.A(_04873_));
 sg13g2_antennanp ANTENNA_2380 (.A(_04873_));
 sg13g2_antennanp ANTENNA_2381 (.A(_04873_));
 sg13g2_antennanp ANTENNA_2382 (.A(_04883_));
 sg13g2_antennanp ANTENNA_2383 (.A(_04912_));
 sg13g2_antennanp ANTENNA_2384 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2385 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2386 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2387 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2388 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2389 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2390 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2391 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2392 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2393 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2394 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2395 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2396 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2397 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2398 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2399 (.A(_04932_));
 sg13g2_antennanp ANTENNA_2400 (.A(_05100_));
 sg13g2_antennanp ANTENNA_2401 (.A(_05100_));
 sg13g2_antennanp ANTENNA_2402 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2403 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2404 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2405 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2406 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2407 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2408 (.A(_05102_));
 sg13g2_antennanp ANTENNA_2409 (.A(_05118_));
 sg13g2_antennanp ANTENNA_2410 (.A(_05124_));
 sg13g2_antennanp ANTENNA_2411 (.A(_05128_));
 sg13g2_antennanp ANTENNA_2412 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2413 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2414 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2415 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2416 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2417 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2418 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2419 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2420 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2421 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2422 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2423 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2424 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2425 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2426 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2427 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2428 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2429 (.A(_05130_));
 sg13g2_antennanp ANTENNA_2430 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2431 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2432 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2433 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2434 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2435 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2436 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2437 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2438 (.A(_05134_));
 sg13g2_antennanp ANTENNA_2439 (.A(_05136_));
 sg13g2_antennanp ANTENNA_2440 (.A(_05198_));
 sg13g2_antennanp ANTENNA_2441 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2442 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2443 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2444 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2445 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2446 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2447 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2448 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2449 (.A(_05205_));
 sg13g2_antennanp ANTENNA_2450 (.A(_05209_));
 sg13g2_antennanp ANTENNA_2451 (.A(_05238_));
 sg13g2_antennanp ANTENNA_2452 (.A(_05238_));
 sg13g2_antennanp ANTENNA_2453 (.A(_05238_));
 sg13g2_antennanp ANTENNA_2454 (.A(_05238_));
 sg13g2_antennanp ANTENNA_2455 (.A(_05252_));
 sg13g2_antennanp ANTENNA_2456 (.A(_05258_));
 sg13g2_antennanp ANTENNA_2457 (.A(_05286_));
 sg13g2_antennanp ANTENNA_2458 (.A(_05302_));
 sg13g2_antennanp ANTENNA_2459 (.A(_05302_));
 sg13g2_antennanp ANTENNA_2460 (.A(_05302_));
 sg13g2_antennanp ANTENNA_2461 (.A(_05302_));
 sg13g2_antennanp ANTENNA_2462 (.A(_05302_));
 sg13g2_antennanp ANTENNA_2463 (.A(_05302_));
 sg13g2_antennanp ANTENNA_2464 (.A(_05318_));
 sg13g2_antennanp ANTENNA_2465 (.A(_05328_));
 sg13g2_antennanp ANTENNA_2466 (.A(_05339_));
 sg13g2_antennanp ANTENNA_2467 (.A(_05342_));
 sg13g2_antennanp ANTENNA_2468 (.A(_05342_));
 sg13g2_antennanp ANTENNA_2469 (.A(_05342_));
 sg13g2_antennanp ANTENNA_2470 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2471 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2472 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2473 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2474 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2475 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2476 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2477 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2478 (.A(_05344_));
 sg13g2_antennanp ANTENNA_2479 (.A(_05350_));
 sg13g2_antennanp ANTENNA_2480 (.A(_05389_));
 sg13g2_antennanp ANTENNA_2481 (.A(_05404_));
 sg13g2_antennanp ANTENNA_2482 (.A(_05415_));
 sg13g2_antennanp ANTENNA_2483 (.A(_05424_));
 sg13g2_antennanp ANTENNA_2484 (.A(_05424_));
 sg13g2_antennanp ANTENNA_2485 (.A(_05424_));
 sg13g2_antennanp ANTENNA_2486 (.A(_05424_));
 sg13g2_antennanp ANTENNA_2487 (.A(_05459_));
 sg13g2_antennanp ANTENNA_2488 (.A(_05500_));
 sg13g2_antennanp ANTENNA_2489 (.A(_05576_));
 sg13g2_antennanp ANTENNA_2490 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2491 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2492 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2493 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2494 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2495 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2496 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2497 (.A(_05609_));
 sg13g2_antennanp ANTENNA_2498 (.A(_05611_));
 sg13g2_antennanp ANTENNA_2499 (.A(_05633_));
 sg13g2_antennanp ANTENNA_2500 (.A(_05681_));
 sg13g2_antennanp ANTENNA_2501 (.A(_05681_));
 sg13g2_antennanp ANTENNA_2502 (.A(_05726_));
 sg13g2_antennanp ANTENNA_2503 (.A(_05750_));
 sg13g2_antennanp ANTENNA_2504 (.A(_05777_));
 sg13g2_antennanp ANTENNA_2505 (.A(_05814_));
 sg13g2_antennanp ANTENNA_2506 (.A(_05816_));
 sg13g2_antennanp ANTENNA_2507 (.A(_05818_));
 sg13g2_antennanp ANTENNA_2508 (.A(_05827_));
 sg13g2_antennanp ANTENNA_2509 (.A(_05829_));
 sg13g2_antennanp ANTENNA_2510 (.A(_05874_));
 sg13g2_antennanp ANTENNA_2511 (.A(_05886_));
 sg13g2_antennanp ANTENNA_2512 (.A(_05890_));
 sg13g2_antennanp ANTENNA_2513 (.A(_05904_));
 sg13g2_antennanp ANTENNA_2514 (.A(_05924_));
 sg13g2_antennanp ANTENNA_2515 (.A(_05939_));
 sg13g2_antennanp ANTENNA_2516 (.A(_05946_));
 sg13g2_antennanp ANTENNA_2517 (.A(_05951_));
 sg13g2_antennanp ANTENNA_2518 (.A(_05957_));
 sg13g2_antennanp ANTENNA_2519 (.A(_05997_));
 sg13g2_antennanp ANTENNA_2520 (.A(_05998_));
 sg13g2_antennanp ANTENNA_2521 (.A(_05998_));
 sg13g2_antennanp ANTENNA_2522 (.A(_06018_));
 sg13g2_antennanp ANTENNA_2523 (.A(_06023_));
 sg13g2_antennanp ANTENNA_2524 (.A(_06046_));
 sg13g2_antennanp ANTENNA_2525 (.A(_06050_));
 sg13g2_antennanp ANTENNA_2526 (.A(_06050_));
 sg13g2_antennanp ANTENNA_2527 (.A(_06053_));
 sg13g2_antennanp ANTENNA_2528 (.A(_06064_));
 sg13g2_antennanp ANTENNA_2529 (.A(_06075_));
 sg13g2_antennanp ANTENNA_2530 (.A(_06091_));
 sg13g2_antennanp ANTENNA_2531 (.A(_06116_));
 sg13g2_antennanp ANTENNA_2532 (.A(_06134_));
 sg13g2_antennanp ANTENNA_2533 (.A(_06139_));
 sg13g2_antennanp ANTENNA_2534 (.A(_06146_));
 sg13g2_antennanp ANTENNA_2535 (.A(_06151_));
 sg13g2_antennanp ANTENNA_2536 (.A(_06167_));
 sg13g2_antennanp ANTENNA_2537 (.A(_06179_));
 sg13g2_antennanp ANTENNA_2538 (.A(_06196_));
 sg13g2_antennanp ANTENNA_2539 (.A(_06209_));
 sg13g2_antennanp ANTENNA_2540 (.A(_06225_));
 sg13g2_antennanp ANTENNA_2541 (.A(_06227_));
 sg13g2_antennanp ANTENNA_2542 (.A(_06244_));
 sg13g2_antennanp ANTENNA_2543 (.A(_06249_));
 sg13g2_antennanp ANTENNA_2544 (.A(_06250_));
 sg13g2_antennanp ANTENNA_2545 (.A(_06271_));
 sg13g2_antennanp ANTENNA_2546 (.A(_06271_));
 sg13g2_antennanp ANTENNA_2547 (.A(_06281_));
 sg13g2_antennanp ANTENNA_2548 (.A(_06290_));
 sg13g2_antennanp ANTENNA_2549 (.A(_06300_));
 sg13g2_antennanp ANTENNA_2550 (.A(_06322_));
 sg13g2_antennanp ANTENNA_2551 (.A(_06324_));
 sg13g2_antennanp ANTENNA_2552 (.A(_06328_));
 sg13g2_antennanp ANTENNA_2553 (.A(_06334_));
 sg13g2_antennanp ANTENNA_2554 (.A(_06335_));
 sg13g2_antennanp ANTENNA_2555 (.A(_06342_));
 sg13g2_antennanp ANTENNA_2556 (.A(_06347_));
 sg13g2_antennanp ANTENNA_2557 (.A(_06361_));
 sg13g2_antennanp ANTENNA_2558 (.A(_06366_));
 sg13g2_antennanp ANTENNA_2559 (.A(_06372_));
 sg13g2_antennanp ANTENNA_2560 (.A(_06374_));
 sg13g2_antennanp ANTENNA_2561 (.A(_06391_));
 sg13g2_antennanp ANTENNA_2562 (.A(_06396_));
 sg13g2_antennanp ANTENNA_2563 (.A(_06397_));
 sg13g2_antennanp ANTENNA_2564 (.A(_06417_));
 sg13g2_antennanp ANTENNA_2565 (.A(_06422_));
 sg13g2_antennanp ANTENNA_2566 (.A(_06440_));
 sg13g2_antennanp ANTENNA_2567 (.A(_06448_));
 sg13g2_antennanp ANTENNA_2568 (.A(_06463_));
 sg13g2_antennanp ANTENNA_2569 (.A(_06463_));
 sg13g2_antennanp ANTENNA_2570 (.A(_06467_));
 sg13g2_antennanp ANTENNA_2571 (.A(_06484_));
 sg13g2_antennanp ANTENNA_2572 (.A(_06492_));
 sg13g2_antennanp ANTENNA_2573 (.A(_06497_));
 sg13g2_antennanp ANTENNA_2574 (.A(_06504_));
 sg13g2_antennanp ANTENNA_2575 (.A(_06506_));
 sg13g2_antennanp ANTENNA_2576 (.A(_06512_));
 sg13g2_antennanp ANTENNA_2577 (.A(_06517_));
 sg13g2_antennanp ANTENNA_2578 (.A(_06522_));
 sg13g2_antennanp ANTENNA_2579 (.A(_06523_));
 sg13g2_antennanp ANTENNA_2580 (.A(_06546_));
 sg13g2_antennanp ANTENNA_2581 (.A(_06548_));
 sg13g2_antennanp ANTENNA_2582 (.A(_06559_));
 sg13g2_antennanp ANTENNA_2583 (.A(_06588_));
 sg13g2_antennanp ANTENNA_2584 (.A(_06589_));
 sg13g2_antennanp ANTENNA_2585 (.A(_06596_));
 sg13g2_antennanp ANTENNA_2586 (.A(_06621_));
 sg13g2_antennanp ANTENNA_2587 (.A(_06640_));
 sg13g2_antennanp ANTENNA_2588 (.A(_06658_));
 sg13g2_antennanp ANTENNA_2589 (.A(_06667_));
 sg13g2_antennanp ANTENNA_2590 (.A(_06679_));
 sg13g2_antennanp ANTENNA_2591 (.A(_06679_));
 sg13g2_antennanp ANTENNA_2592 (.A(_06682_));
 sg13g2_antennanp ANTENNA_2593 (.A(_06684_));
 sg13g2_antennanp ANTENNA_2594 (.A(_06687_));
 sg13g2_antennanp ANTENNA_2595 (.A(_06688_));
 sg13g2_antennanp ANTENNA_2596 (.A(_06701_));
 sg13g2_antennanp ANTENNA_2597 (.A(_06712_));
 sg13g2_antennanp ANTENNA_2598 (.A(_06732_));
 sg13g2_antennanp ANTENNA_2599 (.A(_06745_));
 sg13g2_antennanp ANTENNA_2600 (.A(_06758_));
 sg13g2_antennanp ANTENNA_2601 (.A(_06761_));
 sg13g2_antennanp ANTENNA_2602 (.A(_06761_));
 sg13g2_antennanp ANTENNA_2603 (.A(_06764_));
 sg13g2_antennanp ANTENNA_2604 (.A(_06768_));
 sg13g2_antennanp ANTENNA_2605 (.A(_06775_));
 sg13g2_antennanp ANTENNA_2606 (.A(_06813_));
 sg13g2_antennanp ANTENNA_2607 (.A(_06830_));
 sg13g2_antennanp ANTENNA_2608 (.A(_06830_));
 sg13g2_antennanp ANTENNA_2609 (.A(_06834_));
 sg13g2_antennanp ANTENNA_2610 (.A(_06844_));
 sg13g2_antennanp ANTENNA_2611 (.A(_06849_));
 sg13g2_antennanp ANTENNA_2612 (.A(_06926_));
 sg13g2_antennanp ANTENNA_2613 (.A(_06926_));
 sg13g2_antennanp ANTENNA_2614 (.A(_07040_));
 sg13g2_antennanp ANTENNA_2615 (.A(_07040_));
 sg13g2_antennanp ANTENNA_2616 (.A(_07057_));
 sg13g2_antennanp ANTENNA_2617 (.A(_07085_));
 sg13g2_antennanp ANTENNA_2618 (.A(_07098_));
 sg13g2_antennanp ANTENNA_2619 (.A(_07154_));
 sg13g2_antennanp ANTENNA_2620 (.A(_07170_));
 sg13g2_antennanp ANTENNA_2621 (.A(_07243_));
 sg13g2_antennanp ANTENNA_2622 (.A(_07258_));
 sg13g2_antennanp ANTENNA_2623 (.A(_07273_));
 sg13g2_antennanp ANTENNA_2624 (.A(_07316_));
 sg13g2_antennanp ANTENNA_2625 (.A(_07331_));
 sg13g2_antennanp ANTENNA_2626 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2627 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2628 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2629 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2630 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2631 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2632 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2633 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2634 (.A(_07534_));
 sg13g2_antennanp ANTENNA_2635 (.A(_07663_));
 sg13g2_antennanp ANTENNA_2636 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2637 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2638 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2639 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2640 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2641 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2642 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2643 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2644 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2645 (.A(_09301_));
 sg13g2_antennanp ANTENNA_2646 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2647 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2648 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2649 (.A(_09573_));
 sg13g2_antennanp ANTENNA_2650 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2651 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2652 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2653 (.A(_09599_));
 sg13g2_antennanp ANTENNA_2654 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2655 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2656 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2657 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2658 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2659 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2660 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2661 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2662 (.A(_09910_));
 sg13g2_antennanp ANTENNA_2663 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2664 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2665 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2666 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2667 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2668 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2669 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2670 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2671 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2672 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2673 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2674 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2675 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2676 (.A(_09960_));
 sg13g2_antennanp ANTENNA_2677 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2678 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2679 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2680 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2681 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2682 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2683 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2684 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2685 (.A(_10009_));
 sg13g2_antennanp ANTENNA_2686 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2687 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2688 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2689 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2690 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2691 (.A(_10032_));
 sg13g2_antennanp ANTENNA_2692 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2693 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2694 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2695 (.A(_10074_));
 sg13g2_antennanp ANTENNA_2696 (.A(_10077_));
 sg13g2_antennanp ANTENNA_2697 (.A(_10077_));
 sg13g2_antennanp ANTENNA_2698 (.A(_10077_));
 sg13g2_antennanp ANTENNA_2699 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2700 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2701 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2702 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2703 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2704 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2705 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2706 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2707 (.A(_10085_));
 sg13g2_antennanp ANTENNA_2708 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2709 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2710 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2711 (.A(_10092_));
 sg13g2_antennanp ANTENNA_2712 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2713 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2714 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2715 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2716 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2717 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2718 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2719 (.A(_10151_));
 sg13g2_antennanp ANTENNA_2720 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2721 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2722 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2723 (.A(_10404_));
 sg13g2_antennanp ANTENNA_2724 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2725 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2726 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2727 (.A(_10435_));
 sg13g2_antennanp ANTENNA_2728 (.A(_10460_));
 sg13g2_antennanp ANTENNA_2729 (.A(_10460_));
 sg13g2_antennanp ANTENNA_2730 (.A(_10460_));
 sg13g2_antennanp ANTENNA_2731 (.A(_10460_));
 sg13g2_antennanp ANTENNA_2732 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2733 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2734 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2735 (.A(\top_ihp.oisc.regs[2][0] ));
 sg13g2_antennanp ANTENNA_2736 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2737 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2738 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2739 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_2740 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2741 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2742 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2743 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_2744 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2745 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2746 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2747 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2748 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2749 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2750 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2751 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2752 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_2753 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2754 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2755 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2756 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2757 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2758 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2759 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2760 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2761 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2762 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2763 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2764 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2765 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2766 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2767 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_2768 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_2769 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_2770 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_2771 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_2772 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_2773 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_2774 (.A(\top_ihp.oisc.regs[32][9] ));
 sg13g2_antennanp ANTENNA_2775 (.A(\top_ihp.ram_cs_o ));
 sg13g2_antennanp ANTENNA_2776 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_2777 (.A(net1));
 sg13g2_antennanp ANTENNA_2778 (.A(net1));
 sg13g2_antennanp ANTENNA_2779 (.A(net1));
 sg13g2_antennanp ANTENNA_2780 (.A(net9));
 sg13g2_antennanp ANTENNA_2781 (.A(net47));
 sg13g2_antennanp ANTENNA_2782 (.A(net47));
 sg13g2_antennanp ANTENNA_2783 (.A(net47));
 sg13g2_antennanp ANTENNA_2784 (.A(net47));
 sg13g2_antennanp ANTENNA_2785 (.A(net47));
 sg13g2_antennanp ANTENNA_2786 (.A(net47));
 sg13g2_antennanp ANTENNA_2787 (.A(net47));
 sg13g2_antennanp ANTENNA_2788 (.A(net47));
 sg13g2_antennanp ANTENNA_2789 (.A(net47));
 sg13g2_antennanp ANTENNA_2790 (.A(net47));
 sg13g2_antennanp ANTENNA_2791 (.A(net47));
 sg13g2_antennanp ANTENNA_2792 (.A(net47));
 sg13g2_antennanp ANTENNA_2793 (.A(net47));
 sg13g2_antennanp ANTENNA_2794 (.A(net47));
 sg13g2_antennanp ANTENNA_2795 (.A(net47));
 sg13g2_antennanp ANTENNA_2796 (.A(net47));
 sg13g2_antennanp ANTENNA_2797 (.A(net47));
 sg13g2_antennanp ANTENNA_2798 (.A(net62));
 sg13g2_antennanp ANTENNA_2799 (.A(net62));
 sg13g2_antennanp ANTENNA_2800 (.A(net62));
 sg13g2_antennanp ANTENNA_2801 (.A(net62));
 sg13g2_antennanp ANTENNA_2802 (.A(net62));
 sg13g2_antennanp ANTENNA_2803 (.A(net62));
 sg13g2_antennanp ANTENNA_2804 (.A(net62));
 sg13g2_antennanp ANTENNA_2805 (.A(net62));
 sg13g2_antennanp ANTENNA_2806 (.A(net62));
 sg13g2_antennanp ANTENNA_2807 (.A(net136));
 sg13g2_antennanp ANTENNA_2808 (.A(net136));
 sg13g2_antennanp ANTENNA_2809 (.A(net136));
 sg13g2_antennanp ANTENNA_2810 (.A(net136));
 sg13g2_antennanp ANTENNA_2811 (.A(net136));
 sg13g2_antennanp ANTENNA_2812 (.A(net136));
 sg13g2_antennanp ANTENNA_2813 (.A(net136));
 sg13g2_antennanp ANTENNA_2814 (.A(net136));
 sg13g2_antennanp ANTENNA_2815 (.A(net136));
 sg13g2_antennanp ANTENNA_2816 (.A(net136));
 sg13g2_antennanp ANTENNA_2817 (.A(net136));
 sg13g2_antennanp ANTENNA_2818 (.A(net136));
 sg13g2_antennanp ANTENNA_2819 (.A(net136));
 sg13g2_antennanp ANTENNA_2820 (.A(net136));
 sg13g2_antennanp ANTENNA_2821 (.A(net136));
 sg13g2_antennanp ANTENNA_2822 (.A(net136));
 sg13g2_antennanp ANTENNA_2823 (.A(net142));
 sg13g2_antennanp ANTENNA_2824 (.A(net142));
 sg13g2_antennanp ANTENNA_2825 (.A(net142));
 sg13g2_antennanp ANTENNA_2826 (.A(net142));
 sg13g2_antennanp ANTENNA_2827 (.A(net142));
 sg13g2_antennanp ANTENNA_2828 (.A(net142));
 sg13g2_antennanp ANTENNA_2829 (.A(net142));
 sg13g2_antennanp ANTENNA_2830 (.A(net142));
 sg13g2_antennanp ANTENNA_2831 (.A(net142));
 sg13g2_antennanp ANTENNA_2832 (.A(net235));
 sg13g2_antennanp ANTENNA_2833 (.A(net235));
 sg13g2_antennanp ANTENNA_2834 (.A(net235));
 sg13g2_antennanp ANTENNA_2835 (.A(net235));
 sg13g2_antennanp ANTENNA_2836 (.A(net235));
 sg13g2_antennanp ANTENNA_2837 (.A(net235));
 sg13g2_antennanp ANTENNA_2838 (.A(net235));
 sg13g2_antennanp ANTENNA_2839 (.A(net235));
 sg13g2_antennanp ANTENNA_2840 (.A(net235));
 sg13g2_antennanp ANTENNA_2841 (.A(net235));
 sg13g2_antennanp ANTENNA_2842 (.A(net235));
 sg13g2_antennanp ANTENNA_2843 (.A(net235));
 sg13g2_antennanp ANTENNA_2844 (.A(net334));
 sg13g2_antennanp ANTENNA_2845 (.A(net334));
 sg13g2_antennanp ANTENNA_2846 (.A(net334));
 sg13g2_antennanp ANTENNA_2847 (.A(net334));
 sg13g2_antennanp ANTENNA_2848 (.A(net334));
 sg13g2_antennanp ANTENNA_2849 (.A(net334));
 sg13g2_antennanp ANTENNA_2850 (.A(net334));
 sg13g2_antennanp ANTENNA_2851 (.A(net334));
 sg13g2_antennanp ANTENNA_2852 (.A(net334));
 sg13g2_antennanp ANTENNA_2853 (.A(net347));
 sg13g2_antennanp ANTENNA_2854 (.A(net347));
 sg13g2_antennanp ANTENNA_2855 (.A(net347));
 sg13g2_antennanp ANTENNA_2856 (.A(net347));
 sg13g2_antennanp ANTENNA_2857 (.A(net347));
 sg13g2_antennanp ANTENNA_2858 (.A(net347));
 sg13g2_antennanp ANTENNA_2859 (.A(net347));
 sg13g2_antennanp ANTENNA_2860 (.A(net347));
 sg13g2_antennanp ANTENNA_2861 (.A(net412));
 sg13g2_antennanp ANTENNA_2862 (.A(net412));
 sg13g2_antennanp ANTENNA_2863 (.A(net412));
 sg13g2_antennanp ANTENNA_2864 (.A(net412));
 sg13g2_antennanp ANTENNA_2865 (.A(net412));
 sg13g2_antennanp ANTENNA_2866 (.A(net412));
 sg13g2_antennanp ANTENNA_2867 (.A(net412));
 sg13g2_antennanp ANTENNA_2868 (.A(net412));
 sg13g2_antennanp ANTENNA_2869 (.A(net412));
 sg13g2_antennanp ANTENNA_2870 (.A(net420));
 sg13g2_antennanp ANTENNA_2871 (.A(net420));
 sg13g2_antennanp ANTENNA_2872 (.A(net420));
 sg13g2_antennanp ANTENNA_2873 (.A(net420));
 sg13g2_antennanp ANTENNA_2874 (.A(net420));
 sg13g2_antennanp ANTENNA_2875 (.A(net420));
 sg13g2_antennanp ANTENNA_2876 (.A(net420));
 sg13g2_antennanp ANTENNA_2877 (.A(net420));
 sg13g2_antennanp ANTENNA_2878 (.A(net420));
 sg13g2_antennanp ANTENNA_2879 (.A(net420));
 sg13g2_antennanp ANTENNA_2880 (.A(net420));
 sg13g2_antennanp ANTENNA_2881 (.A(net420));
 sg13g2_antennanp ANTENNA_2882 (.A(net420));
 sg13g2_antennanp ANTENNA_2883 (.A(net420));
 sg13g2_antennanp ANTENNA_2884 (.A(net420));
 sg13g2_antennanp ANTENNA_2885 (.A(net420));
 sg13g2_antennanp ANTENNA_2886 (.A(net420));
 sg13g2_antennanp ANTENNA_2887 (.A(net420));
 sg13g2_antennanp ANTENNA_2888 (.A(net420));
 sg13g2_antennanp ANTENNA_2889 (.A(net420));
 sg13g2_antennanp ANTENNA_2890 (.A(net420));
 sg13g2_antennanp ANTENNA_2891 (.A(net420));
 sg13g2_antennanp ANTENNA_2892 (.A(net454));
 sg13g2_antennanp ANTENNA_2893 (.A(net454));
 sg13g2_antennanp ANTENNA_2894 (.A(net454));
 sg13g2_antennanp ANTENNA_2895 (.A(net454));
 sg13g2_antennanp ANTENNA_2896 (.A(net454));
 sg13g2_antennanp ANTENNA_2897 (.A(net454));
 sg13g2_antennanp ANTENNA_2898 (.A(net454));
 sg13g2_antennanp ANTENNA_2899 (.A(net454));
 sg13g2_antennanp ANTENNA_2900 (.A(net454));
 sg13g2_antennanp ANTENNA_2901 (.A(net474));
 sg13g2_antennanp ANTENNA_2902 (.A(net474));
 sg13g2_antennanp ANTENNA_2903 (.A(net474));
 sg13g2_antennanp ANTENNA_2904 (.A(net474));
 sg13g2_antennanp ANTENNA_2905 (.A(net474));
 sg13g2_antennanp ANTENNA_2906 (.A(net474));
 sg13g2_antennanp ANTENNA_2907 (.A(net474));
 sg13g2_antennanp ANTENNA_2908 (.A(net474));
 sg13g2_antennanp ANTENNA_2909 (.A(net480));
 sg13g2_antennanp ANTENNA_2910 (.A(net480));
 sg13g2_antennanp ANTENNA_2911 (.A(net480));
 sg13g2_antennanp ANTENNA_2912 (.A(net480));
 sg13g2_antennanp ANTENNA_2913 (.A(net480));
 sg13g2_antennanp ANTENNA_2914 (.A(net480));
 sg13g2_antennanp ANTENNA_2915 (.A(net480));
 sg13g2_antennanp ANTENNA_2916 (.A(net480));
 sg13g2_antennanp ANTENNA_2917 (.A(net480));
 sg13g2_antennanp ANTENNA_2918 (.A(net663));
 sg13g2_antennanp ANTENNA_2919 (.A(net663));
 sg13g2_antennanp ANTENNA_2920 (.A(net663));
 sg13g2_antennanp ANTENNA_2921 (.A(net663));
 sg13g2_antennanp ANTENNA_2922 (.A(net663));
 sg13g2_antennanp ANTENNA_2923 (.A(net663));
 sg13g2_antennanp ANTENNA_2924 (.A(net663));
 sg13g2_antennanp ANTENNA_2925 (.A(net663));
 sg13g2_antennanp ANTENNA_2926 (.A(net663));
 sg13g2_antennanp ANTENNA_2927 (.A(net735));
 sg13g2_antennanp ANTENNA_2928 (.A(net735));
 sg13g2_antennanp ANTENNA_2929 (.A(net735));
 sg13g2_antennanp ANTENNA_2930 (.A(net735));
 sg13g2_antennanp ANTENNA_2931 (.A(net735));
 sg13g2_antennanp ANTENNA_2932 (.A(net735));
 sg13g2_antennanp ANTENNA_2933 (.A(net735));
 sg13g2_antennanp ANTENNA_2934 (.A(net735));
 sg13g2_antennanp ANTENNA_2935 (.A(net735));
 sg13g2_antennanp ANTENNA_2936 (.A(_00294_));
 sg13g2_antennanp ANTENNA_2937 (.A(_00294_));
 sg13g2_antennanp ANTENNA_2938 (.A(_00296_));
 sg13g2_antennanp ANTENNA_2939 (.A(_00299_));
 sg13g2_antennanp ANTENNA_2940 (.A(_00300_));
 sg13g2_antennanp ANTENNA_2941 (.A(_00305_));
 sg13g2_antennanp ANTENNA_2942 (.A(_00307_));
 sg13g2_antennanp ANTENNA_2943 (.A(_00311_));
 sg13g2_antennanp ANTENNA_2944 (.A(_00311_));
 sg13g2_antennanp ANTENNA_2945 (.A(_00316_));
 sg13g2_antennanp ANTENNA_2946 (.A(_00319_));
 sg13g2_antennanp ANTENNA_2947 (.A(_00320_));
 sg13g2_antennanp ANTENNA_2948 (.A(_00322_));
 sg13g2_antennanp ANTENNA_2949 (.A(_00322_));
 sg13g2_antennanp ANTENNA_2950 (.A(_00324_));
 sg13g2_antennanp ANTENNA_2951 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2952 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2953 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2954 (.A(_02777_));
 sg13g2_antennanp ANTENNA_2955 (.A(_03021_));
 sg13g2_antennanp ANTENNA_2956 (.A(_03021_));
 sg13g2_antennanp ANTENNA_2957 (.A(_03021_));
 sg13g2_antennanp ANTENNA_2958 (.A(_03713_));
 sg13g2_antennanp ANTENNA_2959 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2960 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2961 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2962 (.A(_04741_));
 sg13g2_antennanp ANTENNA_2963 (.A(_04847_));
 sg13g2_antennanp ANTENNA_2964 (.A(_04847_));
 sg13g2_antennanp ANTENNA_2965 (.A(_04847_));
 sg13g2_antennanp ANTENNA_2966 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2967 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2968 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2969 (.A(_04851_));
 sg13g2_antennanp ANTENNA_2970 (.A(_04857_));
 sg13g2_antennanp ANTENNA_2971 (.A(_04873_));
 sg13g2_antennanp ANTENNA_2972 (.A(_04873_));
 sg13g2_antennanp ANTENNA_2973 (.A(_04873_));
 sg13g2_antennanp ANTENNA_2974 (.A(_04883_));
 sg13g2_antennanp ANTENNA_2975 (.A(_04912_));
 sg13g2_antennanp ANTENNA_2976 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2977 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2978 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2979 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2980 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2981 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2982 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2983 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2984 (.A(_04917_));
 sg13g2_antennanp ANTENNA_2985 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2986 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2987 (.A(_04921_));
 sg13g2_antennanp ANTENNA_2988 (.A(_04932_));
 sg13g2_antennanp ANTENNA_2989 (.A(_05012_));
 sg13g2_antennanp ANTENNA_2990 (.A(_05012_));
 sg13g2_antennanp ANTENNA_2991 (.A(_05012_));
 sg13g2_antennanp ANTENNA_2992 (.A(_05012_));
 sg13g2_antennanp ANTENNA_2993 (.A(_05012_));
 sg13g2_antennanp ANTENNA_2994 (.A(_05012_));
 sg13g2_antennanp ANTENNA_2995 (.A(_05024_));
 sg13g2_antennanp ANTENNA_2996 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2997 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2998 (.A(_05101_));
 sg13g2_antennanp ANTENNA_2999 (.A(_05101_));
 sg13g2_antennanp ANTENNA_3000 (.A(_05101_));
 sg13g2_antennanp ANTENNA_3001 (.A(_05101_));
 sg13g2_antennanp ANTENNA_3002 (.A(_05102_));
 sg13g2_antennanp ANTENNA_3003 (.A(_05102_));
 sg13g2_antennanp ANTENNA_3004 (.A(_05118_));
 sg13g2_antennanp ANTENNA_3005 (.A(_05124_));
 sg13g2_antennanp ANTENNA_3006 (.A(_05128_));
 sg13g2_antennanp ANTENNA_3007 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3008 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3009 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3010 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3011 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3012 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3013 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3014 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3015 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3016 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3017 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3018 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3019 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3020 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3021 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3022 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3023 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3024 (.A(_05130_));
 sg13g2_antennanp ANTENNA_3025 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3026 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3027 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3028 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3029 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3030 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3031 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3032 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3033 (.A(_05134_));
 sg13g2_antennanp ANTENNA_3034 (.A(_05136_));
 sg13g2_antennanp ANTENNA_3035 (.A(_05198_));
 sg13g2_antennanp ANTENNA_3036 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3037 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3038 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3039 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3040 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3041 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3042 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3043 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3044 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3045 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3046 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3047 (.A(_05201_));
 sg13g2_antennanp ANTENNA_3048 (.A(_05205_));
 sg13g2_antennanp ANTENNA_3049 (.A(_05209_));
 sg13g2_antennanp ANTENNA_3050 (.A(_05238_));
 sg13g2_antennanp ANTENNA_3051 (.A(_05238_));
 sg13g2_antennanp ANTENNA_3052 (.A(_05238_));
 sg13g2_antennanp ANTENNA_3053 (.A(_05238_));
 sg13g2_antennanp ANTENNA_3054 (.A(_05252_));
 sg13g2_antennanp ANTENNA_3055 (.A(_05258_));
 sg13g2_antennanp ANTENNA_3056 (.A(_05286_));
 sg13g2_antennanp ANTENNA_3057 (.A(_05302_));
 sg13g2_antennanp ANTENNA_3058 (.A(_05302_));
 sg13g2_antennanp ANTENNA_3059 (.A(_05302_));
 sg13g2_antennanp ANTENNA_3060 (.A(_05318_));
 sg13g2_antennanp ANTENNA_3061 (.A(_05318_));
 sg13g2_antennanp ANTENNA_3062 (.A(_05328_));
 sg13g2_antennanp ANTENNA_3063 (.A(_05339_));
 sg13g2_antennanp ANTENNA_3064 (.A(_05342_));
 sg13g2_antennanp ANTENNA_3065 (.A(_05342_));
 sg13g2_antennanp ANTENNA_3066 (.A(_05342_));
 sg13g2_antennanp ANTENNA_3067 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3068 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3069 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3070 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3071 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3072 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3073 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3074 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3075 (.A(_05344_));
 sg13g2_antennanp ANTENNA_3076 (.A(_05350_));
 sg13g2_antennanp ANTENNA_3077 (.A(_05389_));
 sg13g2_antennanp ANTENNA_3078 (.A(_05404_));
 sg13g2_antennanp ANTENNA_3079 (.A(_05415_));
 sg13g2_antennanp ANTENNA_3080 (.A(_05424_));
 sg13g2_antennanp ANTENNA_3081 (.A(_05424_));
 sg13g2_antennanp ANTENNA_3082 (.A(_05424_));
 sg13g2_antennanp ANTENNA_3083 (.A(_05424_));
 sg13g2_antennanp ANTENNA_3084 (.A(_05459_));
 sg13g2_antennanp ANTENNA_3085 (.A(_05500_));
 sg13g2_antennanp ANTENNA_3086 (.A(_05576_));
 sg13g2_antennanp ANTENNA_3087 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3088 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3089 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3090 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3091 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3092 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3093 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3094 (.A(_05609_));
 sg13g2_antennanp ANTENNA_3095 (.A(_05611_));
 sg13g2_antennanp ANTENNA_3096 (.A(_05633_));
 sg13g2_antennanp ANTENNA_3097 (.A(_05657_));
 sg13g2_antennanp ANTENNA_3098 (.A(_05681_));
 sg13g2_antennanp ANTENNA_3099 (.A(_05681_));
 sg13g2_antennanp ANTENNA_3100 (.A(_05726_));
 sg13g2_antennanp ANTENNA_3101 (.A(_05750_));
 sg13g2_antennanp ANTENNA_3102 (.A(_05750_));
 sg13g2_antennanp ANTENNA_3103 (.A(_05777_));
 sg13g2_antennanp ANTENNA_3104 (.A(_05814_));
 sg13g2_antennanp ANTENNA_3105 (.A(_05816_));
 sg13g2_antennanp ANTENNA_3106 (.A(_05818_));
 sg13g2_antennanp ANTENNA_3107 (.A(_05827_));
 sg13g2_antennanp ANTENNA_3108 (.A(_05829_));
 sg13g2_antennanp ANTENNA_3109 (.A(_05874_));
 sg13g2_antennanp ANTENNA_3110 (.A(_05886_));
 sg13g2_antennanp ANTENNA_3111 (.A(_05890_));
 sg13g2_antennanp ANTENNA_3112 (.A(_05904_));
 sg13g2_antennanp ANTENNA_3113 (.A(_05924_));
 sg13g2_antennanp ANTENNA_3114 (.A(_05939_));
 sg13g2_antennanp ANTENNA_3115 (.A(_05946_));
 sg13g2_antennanp ANTENNA_3116 (.A(_05951_));
 sg13g2_antennanp ANTENNA_3117 (.A(_05957_));
 sg13g2_antennanp ANTENNA_3118 (.A(_05998_));
 sg13g2_antennanp ANTENNA_3119 (.A(_05998_));
 sg13g2_antennanp ANTENNA_3120 (.A(_06018_));
 sg13g2_antennanp ANTENNA_3121 (.A(_06023_));
 sg13g2_antennanp ANTENNA_3122 (.A(_06046_));
 sg13g2_antennanp ANTENNA_3123 (.A(_06050_));
 sg13g2_antennanp ANTENNA_3124 (.A(_06053_));
 sg13g2_antennanp ANTENNA_3125 (.A(_06064_));
 sg13g2_antennanp ANTENNA_3126 (.A(_06075_));
 sg13g2_antennanp ANTENNA_3127 (.A(_06091_));
 sg13g2_antennanp ANTENNA_3128 (.A(_06116_));
 sg13g2_antennanp ANTENNA_3129 (.A(_06134_));
 sg13g2_antennanp ANTENNA_3130 (.A(_06134_));
 sg13g2_antennanp ANTENNA_3131 (.A(_06139_));
 sg13g2_antennanp ANTENNA_3132 (.A(_06146_));
 sg13g2_antennanp ANTENNA_3133 (.A(_06146_));
 sg13g2_antennanp ANTENNA_3134 (.A(_06151_));
 sg13g2_antennanp ANTENNA_3135 (.A(_06167_));
 sg13g2_antennanp ANTENNA_3136 (.A(_06179_));
 sg13g2_antennanp ANTENNA_3137 (.A(_06196_));
 sg13g2_antennanp ANTENNA_3138 (.A(_06209_));
 sg13g2_antennanp ANTENNA_3139 (.A(_06225_));
 sg13g2_antennanp ANTENNA_3140 (.A(_06227_));
 sg13g2_antennanp ANTENNA_3141 (.A(_06244_));
 sg13g2_antennanp ANTENNA_3142 (.A(_06249_));
 sg13g2_antennanp ANTENNA_3143 (.A(_06250_));
 sg13g2_antennanp ANTENNA_3144 (.A(_06271_));
 sg13g2_antennanp ANTENNA_3145 (.A(_06271_));
 sg13g2_antennanp ANTENNA_3146 (.A(_06281_));
 sg13g2_antennanp ANTENNA_3147 (.A(_06290_));
 sg13g2_antennanp ANTENNA_3148 (.A(_06300_));
 sg13g2_antennanp ANTENNA_3149 (.A(_06322_));
 sg13g2_antennanp ANTENNA_3150 (.A(_06324_));
 sg13g2_antennanp ANTENNA_3151 (.A(_06328_));
 sg13g2_antennanp ANTENNA_3152 (.A(_06334_));
 sg13g2_antennanp ANTENNA_3153 (.A(_06347_));
 sg13g2_antennanp ANTENNA_3154 (.A(_06351_));
 sg13g2_antennanp ANTENNA_3155 (.A(_06361_));
 sg13g2_antennanp ANTENNA_3156 (.A(_06366_));
 sg13g2_antennanp ANTENNA_3157 (.A(_06372_));
 sg13g2_antennanp ANTENNA_3158 (.A(_06372_));
 sg13g2_antennanp ANTENNA_3159 (.A(_06374_));
 sg13g2_antennanp ANTENNA_3160 (.A(_06391_));
 sg13g2_antennanp ANTENNA_3161 (.A(_06396_));
 sg13g2_antennanp ANTENNA_3162 (.A(_06397_));
 sg13g2_antennanp ANTENNA_3163 (.A(_06417_));
 sg13g2_antennanp ANTENNA_3164 (.A(_06422_));
 sg13g2_antennanp ANTENNA_3165 (.A(_06440_));
 sg13g2_antennanp ANTENNA_3166 (.A(_06448_));
 sg13g2_antennanp ANTENNA_3167 (.A(_06463_));
 sg13g2_antennanp ANTENNA_3168 (.A(_06463_));
 sg13g2_antennanp ANTENNA_3169 (.A(_06467_));
 sg13g2_antennanp ANTENNA_3170 (.A(_06484_));
 sg13g2_antennanp ANTENNA_3171 (.A(_06492_));
 sg13g2_antennanp ANTENNA_3172 (.A(_06497_));
 sg13g2_antennanp ANTENNA_3173 (.A(_06504_));
 sg13g2_antennanp ANTENNA_3174 (.A(_06506_));
 sg13g2_antennanp ANTENNA_3175 (.A(_06512_));
 sg13g2_antennanp ANTENNA_3176 (.A(_06522_));
 sg13g2_antennanp ANTENNA_3177 (.A(_06523_));
 sg13g2_antennanp ANTENNA_3178 (.A(_06546_));
 sg13g2_antennanp ANTENNA_3179 (.A(_06548_));
 sg13g2_antennanp ANTENNA_3180 (.A(_06588_));
 sg13g2_antennanp ANTENNA_3181 (.A(_06589_));
 sg13g2_antennanp ANTENNA_3182 (.A(_06596_));
 sg13g2_antennanp ANTENNA_3183 (.A(_06621_));
 sg13g2_antennanp ANTENNA_3184 (.A(_06640_));
 sg13g2_antennanp ANTENNA_3185 (.A(_06658_));
 sg13g2_antennanp ANTENNA_3186 (.A(_06667_));
 sg13g2_antennanp ANTENNA_3187 (.A(_06679_));
 sg13g2_antennanp ANTENNA_3188 (.A(_06679_));
 sg13g2_antennanp ANTENNA_3189 (.A(_06682_));
 sg13g2_antennanp ANTENNA_3190 (.A(_06684_));
 sg13g2_antennanp ANTENNA_3191 (.A(_06687_));
 sg13g2_antennanp ANTENNA_3192 (.A(_06688_));
 sg13g2_antennanp ANTENNA_3193 (.A(_06701_));
 sg13g2_antennanp ANTENNA_3194 (.A(_06712_));
 sg13g2_antennanp ANTENNA_3195 (.A(_06732_));
 sg13g2_antennanp ANTENNA_3196 (.A(_06745_));
 sg13g2_antennanp ANTENNA_3197 (.A(_06758_));
 sg13g2_antennanp ANTENNA_3198 (.A(_06761_));
 sg13g2_antennanp ANTENNA_3199 (.A(_06761_));
 sg13g2_antennanp ANTENNA_3200 (.A(_06764_));
 sg13g2_antennanp ANTENNA_3201 (.A(_06768_));
 sg13g2_antennanp ANTENNA_3202 (.A(_06775_));
 sg13g2_antennanp ANTENNA_3203 (.A(_06813_));
 sg13g2_antennanp ANTENNA_3204 (.A(_06830_));
 sg13g2_antennanp ANTENNA_3205 (.A(_06830_));
 sg13g2_antennanp ANTENNA_3206 (.A(_06834_));
 sg13g2_antennanp ANTENNA_3207 (.A(_06844_));
 sg13g2_antennanp ANTENNA_3208 (.A(_06849_));
 sg13g2_antennanp ANTENNA_3209 (.A(_06926_));
 sg13g2_antennanp ANTENNA_3210 (.A(_06926_));
 sg13g2_antennanp ANTENNA_3211 (.A(_07040_));
 sg13g2_antennanp ANTENNA_3212 (.A(_07040_));
 sg13g2_antennanp ANTENNA_3213 (.A(_07057_));
 sg13g2_antennanp ANTENNA_3214 (.A(_07085_));
 sg13g2_antennanp ANTENNA_3215 (.A(_07098_));
 sg13g2_antennanp ANTENNA_3216 (.A(_07154_));
 sg13g2_antennanp ANTENNA_3217 (.A(_07170_));
 sg13g2_antennanp ANTENNA_3218 (.A(_07243_));
 sg13g2_antennanp ANTENNA_3219 (.A(_07258_));
 sg13g2_antennanp ANTENNA_3220 (.A(_07316_));
 sg13g2_antennanp ANTENNA_3221 (.A(_07331_));
 sg13g2_antennanp ANTENNA_3222 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3223 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3224 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3225 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3226 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3227 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3228 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3229 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3230 (.A(_07534_));
 sg13g2_antennanp ANTENNA_3231 (.A(_07663_));
 sg13g2_antennanp ANTENNA_3232 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3233 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3234 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3235 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3236 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3237 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3238 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3239 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3240 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3241 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3242 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3243 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3244 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3245 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3246 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3247 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3248 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3249 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3250 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3251 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3252 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3253 (.A(_09082_));
 sg13g2_antennanp ANTENNA_3254 (.A(_09104_));
 sg13g2_antennanp ANTENNA_3255 (.A(_09104_));
 sg13g2_antennanp ANTENNA_3256 (.A(_09104_));
 sg13g2_antennanp ANTENNA_3257 (.A(_09104_));
 sg13g2_antennanp ANTENNA_3258 (.A(_09301_));
 sg13g2_antennanp ANTENNA_3259 (.A(_09301_));
 sg13g2_antennanp ANTENNA_3260 (.A(_09301_));
 sg13g2_antennanp ANTENNA_3261 (.A(_09301_));
 sg13g2_antennanp ANTENNA_3262 (.A(_09301_));
 sg13g2_antennanp ANTENNA_3263 (.A(_09301_));
 sg13g2_antennanp ANTENNA_3264 (.A(_09573_));
 sg13g2_antennanp ANTENNA_3265 (.A(_09573_));
 sg13g2_antennanp ANTENNA_3266 (.A(_09573_));
 sg13g2_antennanp ANTENNA_3267 (.A(_09573_));
 sg13g2_antennanp ANTENNA_3268 (.A(_09599_));
 sg13g2_antennanp ANTENNA_3269 (.A(_09599_));
 sg13g2_antennanp ANTENNA_3270 (.A(_09599_));
 sg13g2_antennanp ANTENNA_3271 (.A(_09599_));
 sg13g2_antennanp ANTENNA_3272 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3273 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3274 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3275 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3276 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3277 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3278 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3279 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3280 (.A(_09910_));
 sg13g2_antennanp ANTENNA_3281 (.A(_09960_));
 sg13g2_antennanp ANTENNA_3282 (.A(_09960_));
 sg13g2_antennanp ANTENNA_3283 (.A(_09960_));
 sg13g2_antennanp ANTENNA_3284 (.A(_09960_));
 sg13g2_antennanp ANTENNA_3285 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3286 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3287 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3288 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3289 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3290 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3291 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3292 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3293 (.A(_10009_));
 sg13g2_antennanp ANTENNA_3294 (.A(_10032_));
 sg13g2_antennanp ANTENNA_3295 (.A(_10032_));
 sg13g2_antennanp ANTENNA_3296 (.A(_10032_));
 sg13g2_antennanp ANTENNA_3297 (.A(_10032_));
 sg13g2_antennanp ANTENNA_3298 (.A(_10074_));
 sg13g2_antennanp ANTENNA_3299 (.A(_10074_));
 sg13g2_antennanp ANTENNA_3300 (.A(_10074_));
 sg13g2_antennanp ANTENNA_3301 (.A(_10074_));
 sg13g2_antennanp ANTENNA_3302 (.A(_10077_));
 sg13g2_antennanp ANTENNA_3303 (.A(_10077_));
 sg13g2_antennanp ANTENNA_3304 (.A(_10077_));
 sg13g2_antennanp ANTENNA_3305 (.A(_10077_));
 sg13g2_antennanp ANTENNA_3306 (.A(_10077_));
 sg13g2_antennanp ANTENNA_3307 (.A(_10077_));
 sg13g2_antennanp ANTENNA_3308 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3309 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3310 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3311 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3312 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3313 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3314 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3315 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3316 (.A(_10085_));
 sg13g2_antennanp ANTENNA_3317 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3318 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3319 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3320 (.A(_10092_));
 sg13g2_antennanp ANTENNA_3321 (.A(_10151_));
 sg13g2_antennanp ANTENNA_3322 (.A(_10151_));
 sg13g2_antennanp ANTENNA_3323 (.A(_10151_));
 sg13g2_antennanp ANTENNA_3324 (.A(_10151_));
 sg13g2_antennanp ANTENNA_3325 (.A(_10404_));
 sg13g2_antennanp ANTENNA_3326 (.A(_10404_));
 sg13g2_antennanp ANTENNA_3327 (.A(_10404_));
 sg13g2_antennanp ANTENNA_3328 (.A(_10404_));
 sg13g2_antennanp ANTENNA_3329 (.A(_10435_));
 sg13g2_antennanp ANTENNA_3330 (.A(_10435_));
 sg13g2_antennanp ANTENNA_3331 (.A(_10435_));
 sg13g2_antennanp ANTENNA_3332 (.A(_10435_));
 sg13g2_antennanp ANTENNA_3333 (.A(_10460_));
 sg13g2_antennanp ANTENNA_3334 (.A(_10460_));
 sg13g2_antennanp ANTENNA_3335 (.A(_10460_));
 sg13g2_antennanp ANTENNA_3336 (.A(_10460_));
 sg13g2_antennanp ANTENNA_3337 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_3338 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_3339 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_3340 (.A(\top_ihp.oisc.regs[32][15] ));
 sg13g2_antennanp ANTENNA_3341 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_3342 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_3343 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_3344 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_3345 (.A(\top_ihp.oisc.regs[32][17] ));
 sg13g2_antennanp ANTENNA_3346 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_3347 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_3348 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_3349 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_3350 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_3351 (.A(\top_ihp.oisc.regs[32][28] ));
 sg13g2_antennanp ANTENNA_3352 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_3353 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_3354 (.A(\top_ihp.oisc.regs[32][4] ));
 sg13g2_antennanp ANTENNA_3355 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3356 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3357 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3358 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3359 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3360 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3361 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3362 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3363 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3364 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3365 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3366 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3367 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3368 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3369 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3370 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3371 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3372 (.A(\top_ihp.oisc.regs[32][7] ));
 sg13g2_antennanp ANTENNA_3373 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_3374 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_3375 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_3376 (.A(\top_ihp.oisc.regs[32][8] ));
 sg13g2_antennanp ANTENNA_3377 (.A(\top_ihp.ram_cs_o ));
 sg13g2_antennanp ANTENNA_3378 (.A(\top_ihp.tx ));
 sg13g2_antennanp ANTENNA_3379 (.A(net1));
 sg13g2_antennanp ANTENNA_3380 (.A(net1));
 sg13g2_antennanp ANTENNA_3381 (.A(net1));
 sg13g2_antennanp ANTENNA_3382 (.A(net9));
 sg13g2_antennanp ANTENNA_3383 (.A(net47));
 sg13g2_antennanp ANTENNA_3384 (.A(net47));
 sg13g2_antennanp ANTENNA_3385 (.A(net47));
 sg13g2_antennanp ANTENNA_3386 (.A(net47));
 sg13g2_antennanp ANTENNA_3387 (.A(net47));
 sg13g2_antennanp ANTENNA_3388 (.A(net47));
 sg13g2_antennanp ANTENNA_3389 (.A(net47));
 sg13g2_antennanp ANTENNA_3390 (.A(net47));
 sg13g2_antennanp ANTENNA_3391 (.A(net47));
 sg13g2_antennanp ANTENNA_3392 (.A(net47));
 sg13g2_antennanp ANTENNA_3393 (.A(net47));
 sg13g2_antennanp ANTENNA_3394 (.A(net47));
 sg13g2_antennanp ANTENNA_3395 (.A(net47));
 sg13g2_antennanp ANTENNA_3396 (.A(net47));
 sg13g2_antennanp ANTENNA_3397 (.A(net47));
 sg13g2_antennanp ANTENNA_3398 (.A(net47));
 sg13g2_antennanp ANTENNA_3399 (.A(net62));
 sg13g2_antennanp ANTENNA_3400 (.A(net62));
 sg13g2_antennanp ANTENNA_3401 (.A(net62));
 sg13g2_antennanp ANTENNA_3402 (.A(net62));
 sg13g2_antennanp ANTENNA_3403 (.A(net62));
 sg13g2_antennanp ANTENNA_3404 (.A(net62));
 sg13g2_antennanp ANTENNA_3405 (.A(net62));
 sg13g2_antennanp ANTENNA_3406 (.A(net62));
 sg13g2_antennanp ANTENNA_3407 (.A(net62));
 sg13g2_antennanp ANTENNA_3408 (.A(net87));
 sg13g2_antennanp ANTENNA_3409 (.A(net87));
 sg13g2_antennanp ANTENNA_3410 (.A(net87));
 sg13g2_antennanp ANTENNA_3411 (.A(net87));
 sg13g2_antennanp ANTENNA_3412 (.A(net87));
 sg13g2_antennanp ANTENNA_3413 (.A(net87));
 sg13g2_antennanp ANTENNA_3414 (.A(net87));
 sg13g2_antennanp ANTENNA_3415 (.A(net87));
 sg13g2_antennanp ANTENNA_3416 (.A(net87));
 sg13g2_antennanp ANTENNA_3417 (.A(net136));
 sg13g2_antennanp ANTENNA_3418 (.A(net136));
 sg13g2_antennanp ANTENNA_3419 (.A(net136));
 sg13g2_antennanp ANTENNA_3420 (.A(net136));
 sg13g2_antennanp ANTENNA_3421 (.A(net136));
 sg13g2_antennanp ANTENNA_3422 (.A(net136));
 sg13g2_antennanp ANTENNA_3423 (.A(net136));
 sg13g2_antennanp ANTENNA_3424 (.A(net136));
 sg13g2_antennanp ANTENNA_3425 (.A(net136));
 sg13g2_antennanp ANTENNA_3426 (.A(net136));
 sg13g2_antennanp ANTENNA_3427 (.A(net136));
 sg13g2_antennanp ANTENNA_3428 (.A(net136));
 sg13g2_antennanp ANTENNA_3429 (.A(net136));
 sg13g2_antennanp ANTENNA_3430 (.A(net136));
 sg13g2_antennanp ANTENNA_3431 (.A(net136));
 sg13g2_antennanp ANTENNA_3432 (.A(net136));
 sg13g2_antennanp ANTENNA_3433 (.A(net136));
 sg13g2_antennanp ANTENNA_3434 (.A(net142));
 sg13g2_antennanp ANTENNA_3435 (.A(net142));
 sg13g2_antennanp ANTENNA_3436 (.A(net142));
 sg13g2_antennanp ANTENNA_3437 (.A(net142));
 sg13g2_antennanp ANTENNA_3438 (.A(net142));
 sg13g2_antennanp ANTENNA_3439 (.A(net142));
 sg13g2_antennanp ANTENNA_3440 (.A(net142));
 sg13g2_antennanp ANTENNA_3441 (.A(net142));
 sg13g2_antennanp ANTENNA_3442 (.A(net142));
 sg13g2_antennanp ANTENNA_3443 (.A(net334));
 sg13g2_antennanp ANTENNA_3444 (.A(net334));
 sg13g2_antennanp ANTENNA_3445 (.A(net334));
 sg13g2_antennanp ANTENNA_3446 (.A(net334));
 sg13g2_antennanp ANTENNA_3447 (.A(net334));
 sg13g2_antennanp ANTENNA_3448 (.A(net334));
 sg13g2_antennanp ANTENNA_3449 (.A(net334));
 sg13g2_antennanp ANTENNA_3450 (.A(net334));
 sg13g2_antennanp ANTENNA_3451 (.A(net334));
 sg13g2_antennanp ANTENNA_3452 (.A(net347));
 sg13g2_antennanp ANTENNA_3453 (.A(net347));
 sg13g2_antennanp ANTENNA_3454 (.A(net347));
 sg13g2_antennanp ANTENNA_3455 (.A(net347));
 sg13g2_antennanp ANTENNA_3456 (.A(net347));
 sg13g2_antennanp ANTENNA_3457 (.A(net347));
 sg13g2_antennanp ANTENNA_3458 (.A(net347));
 sg13g2_antennanp ANTENNA_3459 (.A(net347));
 sg13g2_antennanp ANTENNA_3460 (.A(net412));
 sg13g2_antennanp ANTENNA_3461 (.A(net412));
 sg13g2_antennanp ANTENNA_3462 (.A(net412));
 sg13g2_antennanp ANTENNA_3463 (.A(net412));
 sg13g2_antennanp ANTENNA_3464 (.A(net412));
 sg13g2_antennanp ANTENNA_3465 (.A(net412));
 sg13g2_antennanp ANTENNA_3466 (.A(net412));
 sg13g2_antennanp ANTENNA_3467 (.A(net412));
 sg13g2_antennanp ANTENNA_3468 (.A(net412));
 sg13g2_antennanp ANTENNA_3469 (.A(net420));
 sg13g2_antennanp ANTENNA_3470 (.A(net420));
 sg13g2_antennanp ANTENNA_3471 (.A(net420));
 sg13g2_antennanp ANTENNA_3472 (.A(net420));
 sg13g2_antennanp ANTENNA_3473 (.A(net420));
 sg13g2_antennanp ANTENNA_3474 (.A(net420));
 sg13g2_antennanp ANTENNA_3475 (.A(net420));
 sg13g2_antennanp ANTENNA_3476 (.A(net420));
 sg13g2_antennanp ANTENNA_3477 (.A(net454));
 sg13g2_antennanp ANTENNA_3478 (.A(net454));
 sg13g2_antennanp ANTENNA_3479 (.A(net454));
 sg13g2_antennanp ANTENNA_3480 (.A(net454));
 sg13g2_antennanp ANTENNA_3481 (.A(net454));
 sg13g2_antennanp ANTENNA_3482 (.A(net454));
 sg13g2_antennanp ANTENNA_3483 (.A(net454));
 sg13g2_antennanp ANTENNA_3484 (.A(net454));
 sg13g2_antennanp ANTENNA_3485 (.A(net454));
 sg13g2_antennanp ANTENNA_3486 (.A(net474));
 sg13g2_antennanp ANTENNA_3487 (.A(net474));
 sg13g2_antennanp ANTENNA_3488 (.A(net474));
 sg13g2_antennanp ANTENNA_3489 (.A(net474));
 sg13g2_antennanp ANTENNA_3490 (.A(net474));
 sg13g2_antennanp ANTENNA_3491 (.A(net474));
 sg13g2_antennanp ANTENNA_3492 (.A(net474));
 sg13g2_antennanp ANTENNA_3493 (.A(net474));
 sg13g2_antennanp ANTENNA_3494 (.A(net480));
 sg13g2_antennanp ANTENNA_3495 (.A(net480));
 sg13g2_antennanp ANTENNA_3496 (.A(net480));
 sg13g2_antennanp ANTENNA_3497 (.A(net480));
 sg13g2_antennanp ANTENNA_3498 (.A(net480));
 sg13g2_antennanp ANTENNA_3499 (.A(net480));
 sg13g2_antennanp ANTENNA_3500 (.A(net480));
 sg13g2_antennanp ANTENNA_3501 (.A(net480));
 sg13g2_antennanp ANTENNA_3502 (.A(net480));
 sg13g2_antennanp ANTENNA_3503 (.A(net663));
 sg13g2_antennanp ANTENNA_3504 (.A(net663));
 sg13g2_antennanp ANTENNA_3505 (.A(net663));
 sg13g2_antennanp ANTENNA_3506 (.A(net663));
 sg13g2_antennanp ANTENNA_3507 (.A(net663));
 sg13g2_antennanp ANTENNA_3508 (.A(net663));
 sg13g2_antennanp ANTENNA_3509 (.A(net663));
 sg13g2_antennanp ANTENNA_3510 (.A(net663));
 sg13g2_antennanp ANTENNA_3511 (.A(net663));
 sg13g2_antennanp ANTENNA_3512 (.A(net735));
 sg13g2_antennanp ANTENNA_3513 (.A(net735));
 sg13g2_antennanp ANTENNA_3514 (.A(net735));
 sg13g2_antennanp ANTENNA_3515 (.A(net735));
 sg13g2_antennanp ANTENNA_3516 (.A(net735));
 sg13g2_antennanp ANTENNA_3517 (.A(net735));
 sg13g2_antennanp ANTENNA_3518 (.A(net735));
 sg13g2_antennanp ANTENNA_3519 (.A(net735));
 sg13g2_antennanp ANTENNA_3520 (.A(net735));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_4 FILLER_0_84 ();
 sg13g2_fill_1 FILLER_0_88 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_8 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_130 ();
 sg13g2_decap_8 FILLER_0_137 ();
 sg13g2_decap_8 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_fill_2 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_4 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_8 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_0_433 ();
 sg13g2_decap_8 FILLER_0_440 ();
 sg13g2_decap_8 FILLER_0_447 ();
 sg13g2_decap_8 FILLER_0_454 ();
 sg13g2_decap_8 FILLER_0_461 ();
 sg13g2_decap_8 FILLER_0_468 ();
 sg13g2_decap_8 FILLER_0_475 ();
 sg13g2_decap_8 FILLER_0_482 ();
 sg13g2_decap_8 FILLER_0_489 ();
 sg13g2_decap_8 FILLER_0_496 ();
 sg13g2_decap_8 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_524 ();
 sg13g2_decap_8 FILLER_0_531 ();
 sg13g2_decap_8 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_545 ();
 sg13g2_decap_8 FILLER_0_552 ();
 sg13g2_decap_8 FILLER_0_559 ();
 sg13g2_decap_8 FILLER_0_566 ();
 sg13g2_decap_8 FILLER_0_573 ();
 sg13g2_decap_8 FILLER_0_580 ();
 sg13g2_decap_8 FILLER_0_587 ();
 sg13g2_decap_8 FILLER_0_594 ();
 sg13g2_decap_8 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_608 ();
 sg13g2_decap_8 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_8 FILLER_0_678 ();
 sg13g2_decap_4 FILLER_0_685 ();
 sg13g2_fill_2 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_699 ();
 sg13g2_decap_8 FILLER_0_706 ();
 sg13g2_decap_4 FILLER_0_713 ();
 sg13g2_fill_2 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_decap_4 FILLER_0_737 ();
 sg13g2_fill_2 FILLER_0_741 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_754 ();
 sg13g2_decap_8 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_4 FILLER_0_775 ();
 sg13g2_fill_1 FILLER_0_779 ();
 sg13g2_fill_1 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_862 ();
 sg13g2_decap_8 FILLER_0_869 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_decap_4 FILLER_0_883 ();
 sg13g2_decap_8 FILLER_0_900 ();
 sg13g2_decap_8 FILLER_0_937 ();
 sg13g2_decap_8 FILLER_0_944 ();
 sg13g2_decap_8 FILLER_0_951 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_fill_1 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_decap_8 FILLER_0_1010 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_8 FILLER_0_1024 ();
 sg13g2_fill_2 FILLER_0_1031 ();
 sg13g2_fill_1 FILLER_0_1033 ();
 sg13g2_fill_1 FILLER_0_1038 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_4 FILLER_0_1050 ();
 sg13g2_fill_1 FILLER_0_1054 ();
 sg13g2_decap_8 FILLER_0_1063 ();
 sg13g2_decap_8 FILLER_0_1070 ();
 sg13g2_decap_8 FILLER_0_1077 ();
 sg13g2_decap_8 FILLER_0_1084 ();
 sg13g2_decap_8 FILLER_0_1091 ();
 sg13g2_fill_2 FILLER_0_1098 ();
 sg13g2_fill_1 FILLER_0_1100 ();
 sg13g2_decap_8 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_8 FILLER_0_1158 ();
 sg13g2_decap_4 FILLER_0_1165 ();
 sg13g2_decap_4 FILLER_0_1198 ();
 sg13g2_fill_2 FILLER_0_1202 ();
 sg13g2_decap_8 FILLER_0_1234 ();
 sg13g2_fill_1 FILLER_0_1241 ();
 sg13g2_decap_8 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1279 ();
 sg13g2_decap_4 FILLER_0_1286 ();
 sg13g2_fill_2 FILLER_0_1290 ();
 sg13g2_fill_2 FILLER_0_1296 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1309 ();
 sg13g2_decap_8 FILLER_0_1316 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_4 FILLER_0_1337 ();
 sg13g2_fill_1 FILLER_0_1341 ();
 sg13g2_fill_2 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1363 ();
 sg13g2_decap_8 FILLER_0_1370 ();
 sg13g2_decap_8 FILLER_0_1377 ();
 sg13g2_decap_8 FILLER_0_1384 ();
 sg13g2_decap_8 FILLER_0_1391 ();
 sg13g2_decap_8 FILLER_0_1398 ();
 sg13g2_decap_8 FILLER_0_1405 ();
 sg13g2_decap_8 FILLER_0_1412 ();
 sg13g2_fill_2 FILLER_0_1419 ();
 sg13g2_decap_4 FILLER_0_1447 ();
 sg13g2_fill_2 FILLER_0_1451 ();
 sg13g2_fill_2 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1486 ();
 sg13g2_decap_8 FILLER_0_1493 ();
 sg13g2_decap_8 FILLER_0_1500 ();
 sg13g2_decap_8 FILLER_0_1507 ();
 sg13g2_decap_8 FILLER_0_1514 ();
 sg13g2_decap_8 FILLER_0_1521 ();
 sg13g2_decap_8 FILLER_0_1528 ();
 sg13g2_decap_8 FILLER_0_1535 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_8 FILLER_0_1549 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_decap_8 FILLER_0_1563 ();
 sg13g2_decap_8 FILLER_0_1570 ();
 sg13g2_decap_8 FILLER_0_1577 ();
 sg13g2_decap_8 FILLER_0_1584 ();
 sg13g2_decap_8 FILLER_0_1591 ();
 sg13g2_decap_8 FILLER_0_1598 ();
 sg13g2_decap_8 FILLER_0_1605 ();
 sg13g2_decap_8 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1619 ();
 sg13g2_decap_8 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1633 ();
 sg13g2_decap_8 FILLER_0_1640 ();
 sg13g2_decap_8 FILLER_0_1647 ();
 sg13g2_fill_2 FILLER_0_1654 ();
 sg13g2_fill_1 FILLER_0_1656 ();
 sg13g2_decap_8 FILLER_0_1662 ();
 sg13g2_decap_8 FILLER_0_1669 ();
 sg13g2_decap_8 FILLER_0_1676 ();
 sg13g2_decap_8 FILLER_0_1683 ();
 sg13g2_decap_8 FILLER_0_1690 ();
 sg13g2_decap_8 FILLER_0_1697 ();
 sg13g2_decap_8 FILLER_0_1704 ();
 sg13g2_decap_8 FILLER_0_1711 ();
 sg13g2_decap_8 FILLER_0_1718 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_decap_8 FILLER_0_1739 ();
 sg13g2_decap_8 FILLER_0_1746 ();
 sg13g2_decap_4 FILLER_0_1753 ();
 sg13g2_fill_2 FILLER_0_1757 ();
 sg13g2_fill_1 FILLER_0_1777 ();
 sg13g2_fill_2 FILLER_0_1810 ();
 sg13g2_decap_8 FILLER_0_1817 ();
 sg13g2_decap_8 FILLER_0_1824 ();
 sg13g2_decap_8 FILLER_0_1831 ();
 sg13g2_decap_8 FILLER_0_1838 ();
 sg13g2_decap_8 FILLER_0_1849 ();
 sg13g2_decap_8 FILLER_0_1856 ();
 sg13g2_decap_8 FILLER_0_1863 ();
 sg13g2_decap_8 FILLER_0_1870 ();
 sg13g2_decap_8 FILLER_0_1877 ();
 sg13g2_decap_8 FILLER_0_1884 ();
 sg13g2_decap_8 FILLER_0_1891 ();
 sg13g2_decap_8 FILLER_0_1898 ();
 sg13g2_decap_8 FILLER_0_1905 ();
 sg13g2_decap_8 FILLER_0_1912 ();
 sg13g2_decap_8 FILLER_0_1919 ();
 sg13g2_decap_8 FILLER_0_1926 ();
 sg13g2_decap_8 FILLER_0_1959 ();
 sg13g2_decap_4 FILLER_0_1966 ();
 sg13g2_fill_1 FILLER_0_1970 ();
 sg13g2_decap_8 FILLER_0_2001 ();
 sg13g2_decap_8 FILLER_0_2008 ();
 sg13g2_decap_8 FILLER_0_2015 ();
 sg13g2_decap_8 FILLER_0_2022 ();
 sg13g2_decap_8 FILLER_0_2029 ();
 sg13g2_decap_8 FILLER_0_2036 ();
 sg13g2_decap_8 FILLER_0_2043 ();
 sg13g2_decap_8 FILLER_0_2050 ();
 sg13g2_decap_8 FILLER_0_2057 ();
 sg13g2_decap_8 FILLER_0_2064 ();
 sg13g2_decap_8 FILLER_0_2071 ();
 sg13g2_decap_8 FILLER_0_2078 ();
 sg13g2_decap_8 FILLER_0_2085 ();
 sg13g2_decap_8 FILLER_0_2092 ();
 sg13g2_decap_8 FILLER_0_2099 ();
 sg13g2_decap_4 FILLER_0_2106 ();
 sg13g2_fill_1 FILLER_0_2110 ();
 sg13g2_decap_8 FILLER_0_2115 ();
 sg13g2_decap_8 FILLER_0_2122 ();
 sg13g2_decap_8 FILLER_0_2129 ();
 sg13g2_decap_8 FILLER_0_2136 ();
 sg13g2_decap_8 FILLER_0_2143 ();
 sg13g2_decap_8 FILLER_0_2150 ();
 sg13g2_decap_8 FILLER_0_2157 ();
 sg13g2_decap_8 FILLER_0_2164 ();
 sg13g2_decap_8 FILLER_0_2171 ();
 sg13g2_decap_8 FILLER_0_2178 ();
 sg13g2_decap_8 FILLER_0_2185 ();
 sg13g2_decap_8 FILLER_0_2192 ();
 sg13g2_decap_8 FILLER_0_2199 ();
 sg13g2_decap_8 FILLER_0_2206 ();
 sg13g2_decap_8 FILLER_0_2213 ();
 sg13g2_decap_8 FILLER_0_2220 ();
 sg13g2_decap_8 FILLER_0_2227 ();
 sg13g2_decap_4 FILLER_0_2234 ();
 sg13g2_fill_1 FILLER_0_2238 ();
 sg13g2_decap_8 FILLER_0_2265 ();
 sg13g2_decap_8 FILLER_0_2272 ();
 sg13g2_fill_1 FILLER_0_2279 ();
 sg13g2_decap_8 FILLER_0_2284 ();
 sg13g2_decap_8 FILLER_0_2291 ();
 sg13g2_decap_8 FILLER_0_2298 ();
 sg13g2_decap_8 FILLER_0_2305 ();
 sg13g2_decap_8 FILLER_0_2312 ();
 sg13g2_decap_8 FILLER_0_2319 ();
 sg13g2_decap_8 FILLER_0_2326 ();
 sg13g2_decap_8 FILLER_0_2333 ();
 sg13g2_decap_8 FILLER_0_2340 ();
 sg13g2_decap_8 FILLER_0_2347 ();
 sg13g2_decap_4 FILLER_0_2354 ();
 sg13g2_fill_2 FILLER_0_2358 ();
 sg13g2_decap_8 FILLER_0_2386 ();
 sg13g2_decap_8 FILLER_0_2393 ();
 sg13g2_decap_8 FILLER_0_2400 ();
 sg13g2_decap_8 FILLER_0_2407 ();
 sg13g2_decap_8 FILLER_0_2414 ();
 sg13g2_decap_8 FILLER_0_2421 ();
 sg13g2_decap_8 FILLER_0_2428 ();
 sg13g2_decap_8 FILLER_0_2435 ();
 sg13g2_decap_8 FILLER_0_2442 ();
 sg13g2_decap_8 FILLER_0_2449 ();
 sg13g2_decap_8 FILLER_0_2456 ();
 sg13g2_decap_8 FILLER_0_2463 ();
 sg13g2_decap_8 FILLER_0_2470 ();
 sg13g2_decap_8 FILLER_0_2477 ();
 sg13g2_decap_8 FILLER_0_2484 ();
 sg13g2_decap_8 FILLER_0_2491 ();
 sg13g2_decap_8 FILLER_0_2498 ();
 sg13g2_decap_8 FILLER_0_2505 ();
 sg13g2_decap_8 FILLER_0_2512 ();
 sg13g2_decap_8 FILLER_0_2519 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_8 FILLER_0_2540 ();
 sg13g2_decap_8 FILLER_0_2547 ();
 sg13g2_decap_8 FILLER_0_2554 ();
 sg13g2_decap_8 FILLER_0_2561 ();
 sg13g2_decap_8 FILLER_0_2568 ();
 sg13g2_decap_8 FILLER_0_2575 ();
 sg13g2_decap_8 FILLER_0_2582 ();
 sg13g2_decap_8 FILLER_0_2589 ();
 sg13g2_decap_8 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2603 ();
 sg13g2_decap_8 FILLER_0_2610 ();
 sg13g2_decap_8 FILLER_0_2617 ();
 sg13g2_decap_8 FILLER_0_2624 ();
 sg13g2_decap_8 FILLER_0_2631 ();
 sg13g2_decap_8 FILLER_0_2638 ();
 sg13g2_decap_8 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2652 ();
 sg13g2_decap_8 FILLER_0_2659 ();
 sg13g2_decap_4 FILLER_0_2666 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_49 ();
 sg13g2_decap_4 FILLER_1_89 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_139 ();
 sg13g2_decap_4 FILLER_1_144 ();
 sg13g2_decap_8 FILLER_1_174 ();
 sg13g2_fill_2 FILLER_1_181 ();
 sg13g2_fill_1 FILLER_1_183 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_fill_2 FILLER_1_217 ();
 sg13g2_fill_1 FILLER_1_219 ();
 sg13g2_decap_8 FILLER_1_250 ();
 sg13g2_decap_4 FILLER_1_257 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_decap_4 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_292 ();
 sg13g2_decap_8 FILLER_1_320 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_341 ();
 sg13g2_decap_4 FILLER_1_348 ();
 sg13g2_fill_2 FILLER_1_352 ();
 sg13g2_fill_2 FILLER_1_380 ();
 sg13g2_fill_1 FILLER_1_382 ();
 sg13g2_fill_2 FILLER_1_409 ();
 sg13g2_fill_1 FILLER_1_411 ();
 sg13g2_fill_2 FILLER_1_438 ();
 sg13g2_fill_1 FILLER_1_474 ();
 sg13g2_fill_1 FILLER_1_480 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_fill_2 FILLER_1_646 ();
 sg13g2_fill_1 FILLER_1_678 ();
 sg13g2_fill_2 FILLER_1_726 ();
 sg13g2_fill_2 FILLER_1_732 ();
 sg13g2_fill_2 FILLER_1_760 ();
 sg13g2_fill_1 FILLER_1_762 ();
 sg13g2_fill_2 FILLER_1_789 ();
 sg13g2_fill_1 FILLER_1_821 ();
 sg13g2_decap_8 FILLER_1_904 ();
 sg13g2_decap_4 FILLER_1_911 ();
 sg13g2_fill_2 FILLER_1_915 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_8 FILLER_1_1010 ();
 sg13g2_fill_1 FILLER_1_1017 ();
 sg13g2_fill_2 FILLER_1_1065 ();
 sg13g2_fill_1 FILLER_1_1067 ();
 sg13g2_decap_4 FILLER_1_1094 ();
 sg13g2_fill_2 FILLER_1_1098 ();
 sg13g2_fill_1 FILLER_1_1130 ();
 sg13g2_fill_1 FILLER_1_1165 ();
 sg13g2_decap_8 FILLER_1_1173 ();
 sg13g2_decap_4 FILLER_1_1180 ();
 sg13g2_fill_1 FILLER_1_1184 ();
 sg13g2_decap_4 FILLER_1_1211 ();
 sg13g2_fill_2 FILLER_1_1215 ();
 sg13g2_fill_2 FILLER_1_1251 ();
 sg13g2_decap_8 FILLER_1_1265 ();
 sg13g2_decap_8 FILLER_1_1272 ();
 sg13g2_decap_8 FILLER_1_1279 ();
 sg13g2_fill_1 FILLER_1_1286 ();
 sg13g2_decap_4 FILLER_1_1325 ();
 sg13g2_fill_1 FILLER_1_1329 ();
 sg13g2_fill_2 FILLER_1_1372 ();
 sg13g2_fill_2 FILLER_1_1400 ();
 sg13g2_fill_1 FILLER_1_1402 ();
 sg13g2_fill_1 FILLER_1_1429 ();
 sg13g2_decap_4 FILLER_1_1489 ();
 sg13g2_fill_2 FILLER_1_1519 ();
 sg13g2_fill_1 FILLER_1_1521 ();
 sg13g2_fill_2 FILLER_1_1552 ();
 sg13g2_fill_1 FILLER_1_1554 ();
 sg13g2_decap_8 FILLER_1_1581 ();
 sg13g2_decap_4 FILLER_1_1614 ();
 sg13g2_fill_1 FILLER_1_1618 ();
 sg13g2_fill_1 FILLER_1_1645 ();
 sg13g2_fill_2 FILLER_1_1676 ();
 sg13g2_fill_2 FILLER_1_1718 ();
 sg13g2_decap_8 FILLER_1_1724 ();
 sg13g2_decap_8 FILLER_1_1731 ();
 sg13g2_decap_4 FILLER_1_1738 ();
 sg13g2_fill_1 FILLER_1_1742 ();
 sg13g2_fill_1 FILLER_1_1780 ();
 sg13g2_fill_2 FILLER_1_1828 ();
 sg13g2_fill_1 FILLER_1_1830 ();
 sg13g2_fill_2 FILLER_1_1836 ();
 sg13g2_decap_8 FILLER_1_1864 ();
 sg13g2_decap_8 FILLER_1_1871 ();
 sg13g2_decap_8 FILLER_1_1878 ();
 sg13g2_fill_2 FILLER_1_1885 ();
 sg13g2_fill_1 FILLER_1_1887 ();
 sg13g2_decap_8 FILLER_1_1948 ();
 sg13g2_decap_8 FILLER_1_1955 ();
 sg13g2_decap_8 FILLER_1_1962 ();
 sg13g2_fill_2 FILLER_1_1969 ();
 sg13g2_decap_8 FILLER_1_2001 ();
 sg13g2_decap_8 FILLER_1_2008 ();
 sg13g2_fill_1 FILLER_1_2015 ();
 sg13g2_decap_8 FILLER_1_2025 ();
 sg13g2_fill_2 FILLER_1_2032 ();
 sg13g2_fill_1 FILLER_1_2039 ();
 sg13g2_decap_4 FILLER_1_2092 ();
 sg13g2_fill_2 FILLER_1_2122 ();
 sg13g2_fill_1 FILLER_1_2124 ();
 sg13g2_decap_8 FILLER_1_2151 ();
 sg13g2_decap_4 FILLER_1_2158 ();
 sg13g2_fill_2 FILLER_1_2162 ();
 sg13g2_decap_8 FILLER_1_2169 ();
 sg13g2_decap_8 FILLER_1_2202 ();
 sg13g2_fill_2 FILLER_1_2209 ();
 sg13g2_fill_1 FILLER_1_2211 ();
 sg13g2_fill_1 FILLER_1_2238 ();
 sg13g2_decap_8 FILLER_1_2273 ();
 sg13g2_fill_1 FILLER_1_2285 ();
 sg13g2_fill_1 FILLER_1_2312 ();
 sg13g2_fill_2 FILLER_1_2317 ();
 sg13g2_fill_1 FILLER_1_2345 ();
 sg13g2_fill_2 FILLER_1_2372 ();
 sg13g2_decap_8 FILLER_1_2378 ();
 sg13g2_decap_8 FILLER_1_2385 ();
 sg13g2_decap_8 FILLER_1_2392 ();
 sg13g2_decap_8 FILLER_1_2399 ();
 sg13g2_decap_8 FILLER_1_2406 ();
 sg13g2_decap_8 FILLER_1_2413 ();
 sg13g2_decap_8 FILLER_1_2420 ();
 sg13g2_decap_8 FILLER_1_2427 ();
 sg13g2_decap_8 FILLER_1_2434 ();
 sg13g2_decap_8 FILLER_1_2441 ();
 sg13g2_decap_8 FILLER_1_2448 ();
 sg13g2_decap_8 FILLER_1_2455 ();
 sg13g2_decap_8 FILLER_1_2462 ();
 sg13g2_decap_8 FILLER_1_2469 ();
 sg13g2_decap_8 FILLER_1_2476 ();
 sg13g2_decap_8 FILLER_1_2483 ();
 sg13g2_decap_8 FILLER_1_2490 ();
 sg13g2_decap_8 FILLER_1_2497 ();
 sg13g2_decap_8 FILLER_1_2504 ();
 sg13g2_decap_8 FILLER_1_2511 ();
 sg13g2_decap_8 FILLER_1_2518 ();
 sg13g2_decap_8 FILLER_1_2525 ();
 sg13g2_decap_8 FILLER_1_2532 ();
 sg13g2_decap_8 FILLER_1_2539 ();
 sg13g2_decap_8 FILLER_1_2546 ();
 sg13g2_decap_8 FILLER_1_2553 ();
 sg13g2_decap_8 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2567 ();
 sg13g2_decap_8 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2581 ();
 sg13g2_decap_8 FILLER_1_2588 ();
 sg13g2_decap_8 FILLER_1_2595 ();
 sg13g2_decap_8 FILLER_1_2602 ();
 sg13g2_decap_8 FILLER_1_2609 ();
 sg13g2_decap_8 FILLER_1_2616 ();
 sg13g2_decap_8 FILLER_1_2623 ();
 sg13g2_decap_8 FILLER_1_2630 ();
 sg13g2_decap_8 FILLER_1_2637 ();
 sg13g2_decap_8 FILLER_1_2644 ();
 sg13g2_decap_8 FILLER_1_2651 ();
 sg13g2_decap_8 FILLER_1_2658 ();
 sg13g2_decap_4 FILLER_1_2665 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_93 ();
 sg13g2_fill_1 FILLER_2_120 ();
 sg13g2_fill_1 FILLER_2_129 ();
 sg13g2_fill_1 FILLER_2_134 ();
 sg13g2_fill_2 FILLER_2_143 ();
 sg13g2_fill_1 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_176 ();
 sg13g2_decap_8 FILLER_2_183 ();
 sg13g2_fill_1 FILLER_2_199 ();
 sg13g2_decap_4 FILLER_2_228 ();
 sg13g2_fill_1 FILLER_2_232 ();
 sg13g2_fill_2 FILLER_2_246 ();
 sg13g2_decap_4 FILLER_2_258 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_fill_2 FILLER_2_332 ();
 sg13g2_fill_1 FILLER_2_360 ();
 sg13g2_fill_1 FILLER_2_370 ();
 sg13g2_fill_1 FILLER_2_375 ();
 sg13g2_fill_2 FILLER_2_380 ();
 sg13g2_fill_1 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_2_447 ();
 sg13g2_decap_8 FILLER_2_454 ();
 sg13g2_decap_4 FILLER_2_461 ();
 sg13g2_fill_1 FILLER_2_465 ();
 sg13g2_fill_2 FILLER_2_492 ();
 sg13g2_fill_2 FILLER_2_520 ();
 sg13g2_decap_8 FILLER_2_526 ();
 sg13g2_decap_8 FILLER_2_533 ();
 sg13g2_decap_8 FILLER_2_540 ();
 sg13g2_decap_8 FILLER_2_547 ();
 sg13g2_decap_8 FILLER_2_554 ();
 sg13g2_decap_8 FILLER_2_561 ();
 sg13g2_decap_8 FILLER_2_568 ();
 sg13g2_decap_8 FILLER_2_575 ();
 sg13g2_decap_8 FILLER_2_582 ();
 sg13g2_decap_8 FILLER_2_589 ();
 sg13g2_decap_8 FILLER_2_596 ();
 sg13g2_decap_8 FILLER_2_603 ();
 sg13g2_decap_4 FILLER_2_610 ();
 sg13g2_fill_1 FILLER_2_614 ();
 sg13g2_decap_8 FILLER_2_619 ();
 sg13g2_fill_1 FILLER_2_626 ();
 sg13g2_decap_4 FILLER_2_631 ();
 sg13g2_fill_1 FILLER_2_635 ();
 sg13g2_decap_8 FILLER_2_722 ();
 sg13g2_decap_4 FILLER_2_814 ();
 sg13g2_fill_1 FILLER_2_818 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_4 FILLER_2_830 ();
 sg13g2_fill_1 FILLER_2_834 ();
 sg13g2_decap_4 FILLER_2_839 ();
 sg13g2_fill_1 FILLER_2_851 ();
 sg13g2_fill_2 FILLER_2_856 ();
 sg13g2_decap_8 FILLER_2_918 ();
 sg13g2_decap_4 FILLER_2_925 ();
 sg13g2_fill_2 FILLER_2_933 ();
 sg13g2_fill_2 FILLER_2_965 ();
 sg13g2_fill_1 FILLER_2_996 ();
 sg13g2_fill_2 FILLER_2_1023 ();
 sg13g2_fill_1 FILLER_2_1025 ();
 sg13g2_fill_1 FILLER_2_1104 ();
 sg13g2_fill_1 FILLER_2_1109 ();
 sg13g2_fill_1 FILLER_2_1136 ();
 sg13g2_fill_1 FILLER_2_1163 ();
 sg13g2_decap_8 FILLER_2_1220 ();
 sg13g2_decap_4 FILLER_2_1227 ();
 sg13g2_decap_4 FILLER_2_1248 ();
 sg13g2_fill_2 FILLER_2_1278 ();
 sg13g2_fill_2 FILLER_2_1306 ();
 sg13g2_fill_2 FILLER_2_1312 ();
 sg13g2_decap_4 FILLER_2_1344 ();
 sg13g2_fill_2 FILLER_2_1348 ();
 sg13g2_fill_2 FILLER_2_1384 ();
 sg13g2_fill_1 FILLER_2_1419 ();
 sg13g2_decap_4 FILLER_2_1455 ();
 sg13g2_fill_1 FILLER_2_1459 ();
 sg13g2_fill_1 FILLER_2_1577 ();
 sg13g2_decap_4 FILLER_2_1604 ();
 sg13g2_fill_2 FILLER_2_1608 ();
 sg13g2_decap_8 FILLER_2_1615 ();
 sg13g2_fill_2 FILLER_2_1622 ();
 sg13g2_fill_2 FILLER_2_1629 ();
 sg13g2_fill_1 FILLER_2_1657 ();
 sg13g2_fill_2 FILLER_2_1684 ();
 sg13g2_fill_1 FILLER_2_1686 ();
 sg13g2_fill_2 FILLER_2_1769 ();
 sg13g2_fill_1 FILLER_2_1797 ();
 sg13g2_fill_1 FILLER_2_1803 ();
 sg13g2_fill_1 FILLER_2_1830 ();
 sg13g2_fill_1 FILLER_2_1857 ();
 sg13g2_fill_2 FILLER_2_1884 ();
 sg13g2_fill_1 FILLER_2_1912 ();
 sg13g2_fill_2 FILLER_2_1939 ();
 sg13g2_decap_8 FILLER_2_1945 ();
 sg13g2_decap_8 FILLER_2_1952 ();
 sg13g2_decap_8 FILLER_2_1959 ();
 sg13g2_fill_2 FILLER_2_1966 ();
 sg13g2_decap_4 FILLER_2_1978 ();
 sg13g2_decap_8 FILLER_2_1990 ();
 sg13g2_decap_4 FILLER_2_1997 ();
 sg13g2_decap_8 FILLER_2_2062 ();
 sg13g2_fill_2 FILLER_2_2095 ();
 sg13g2_fill_2 FILLER_2_2106 ();
 sg13g2_decap_4 FILLER_2_2217 ();
 sg13g2_fill_1 FILLER_2_2221 ();
 sg13g2_fill_2 FILLER_2_2227 ();
 sg13g2_decap_4 FILLER_2_2264 ();
 sg13g2_fill_1 FILLER_2_2268 ();
 sg13g2_decap_4 FILLER_2_2274 ();
 sg13g2_fill_2 FILLER_2_2278 ();
 sg13g2_fill_2 FILLER_2_2389 ();
 sg13g2_fill_1 FILLER_2_2391 ();
 sg13g2_decap_8 FILLER_2_2426 ();
 sg13g2_decap_8 FILLER_2_2433 ();
 sg13g2_decap_8 FILLER_2_2440 ();
 sg13g2_decap_8 FILLER_2_2447 ();
 sg13g2_decap_8 FILLER_2_2454 ();
 sg13g2_decap_8 FILLER_2_2461 ();
 sg13g2_decap_8 FILLER_2_2468 ();
 sg13g2_decap_8 FILLER_2_2475 ();
 sg13g2_decap_8 FILLER_2_2482 ();
 sg13g2_decap_8 FILLER_2_2489 ();
 sg13g2_decap_8 FILLER_2_2496 ();
 sg13g2_decap_8 FILLER_2_2503 ();
 sg13g2_decap_8 FILLER_2_2510 ();
 sg13g2_decap_8 FILLER_2_2517 ();
 sg13g2_decap_8 FILLER_2_2524 ();
 sg13g2_decap_8 FILLER_2_2531 ();
 sg13g2_decap_8 FILLER_2_2538 ();
 sg13g2_decap_8 FILLER_2_2545 ();
 sg13g2_decap_8 FILLER_2_2552 ();
 sg13g2_decap_8 FILLER_2_2559 ();
 sg13g2_decap_8 FILLER_2_2566 ();
 sg13g2_decap_8 FILLER_2_2573 ();
 sg13g2_decap_8 FILLER_2_2580 ();
 sg13g2_decap_8 FILLER_2_2587 ();
 sg13g2_decap_8 FILLER_2_2594 ();
 sg13g2_decap_8 FILLER_2_2601 ();
 sg13g2_decap_8 FILLER_2_2608 ();
 sg13g2_decap_8 FILLER_2_2615 ();
 sg13g2_decap_8 FILLER_2_2622 ();
 sg13g2_decap_8 FILLER_2_2629 ();
 sg13g2_decap_8 FILLER_2_2636 ();
 sg13g2_decap_8 FILLER_2_2643 ();
 sg13g2_decap_8 FILLER_2_2650 ();
 sg13g2_decap_8 FILLER_2_2657 ();
 sg13g2_decap_4 FILLER_2_2664 ();
 sg13g2_fill_2 FILLER_2_2668 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_104 ();
 sg13g2_decap_4 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_120 ();
 sg13g2_fill_2 FILLER_3_159 ();
 sg13g2_decap_4 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_173 ();
 sg13g2_decap_4 FILLER_3_180 ();
 sg13g2_fill_2 FILLER_3_184 ();
 sg13g2_decap_4 FILLER_3_224 ();
 sg13g2_fill_1 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_255 ();
 sg13g2_fill_2 FILLER_3_262 ();
 sg13g2_fill_1 FILLER_3_264 ();
 sg13g2_decap_4 FILLER_3_291 ();
 sg13g2_fill_1 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_fill_2 FILLER_3_329 ();
 sg13g2_fill_1 FILLER_3_331 ();
 sg13g2_fill_2 FILLER_3_358 ();
 sg13g2_fill_1 FILLER_3_370 ();
 sg13g2_fill_1 FILLER_3_376 ();
 sg13g2_fill_1 FILLER_3_381 ();
 sg13g2_fill_1 FILLER_3_387 ();
 sg13g2_decap_4 FILLER_3_414 ();
 sg13g2_fill_2 FILLER_3_418 ();
 sg13g2_decap_4 FILLER_3_425 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_4 FILLER_3_435 ();
 sg13g2_decap_8 FILLER_3_443 ();
 sg13g2_decap_8 FILLER_3_450 ();
 sg13g2_decap_4 FILLER_3_457 ();
 sg13g2_fill_2 FILLER_3_461 ();
 sg13g2_decap_4 FILLER_3_468 ();
 sg13g2_fill_1 FILLER_3_472 ();
 sg13g2_decap_8 FILLER_3_498 ();
 sg13g2_decap_8 FILLER_3_505 ();
 sg13g2_decap_8 FILLER_3_512 ();
 sg13g2_decap_8 FILLER_3_519 ();
 sg13g2_decap_8 FILLER_3_526 ();
 sg13g2_decap_8 FILLER_3_533 ();
 sg13g2_decap_8 FILLER_3_540 ();
 sg13g2_decap_8 FILLER_3_547 ();
 sg13g2_decap_8 FILLER_3_554 ();
 sg13g2_decap_8 FILLER_3_561 ();
 sg13g2_decap_8 FILLER_3_568 ();
 sg13g2_decap_8 FILLER_3_575 ();
 sg13g2_decap_8 FILLER_3_582 ();
 sg13g2_decap_8 FILLER_3_589 ();
 sg13g2_decap_8 FILLER_3_596 ();
 sg13g2_decap_4 FILLER_3_603 ();
 sg13g2_fill_1 FILLER_3_607 ();
 sg13g2_decap_8 FILLER_3_674 ();
 sg13g2_fill_2 FILLER_3_681 ();
 sg13g2_fill_1 FILLER_3_709 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_fill_1 FILLER_3_721 ();
 sg13g2_fill_1 FILLER_3_748 ();
 sg13g2_fill_1 FILLER_3_753 ();
 sg13g2_fill_1 FILLER_3_759 ();
 sg13g2_fill_2 FILLER_3_768 ();
 sg13g2_fill_2 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_4 FILLER_3_861 ();
 sg13g2_fill_1 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_874 ();
 sg13g2_decap_4 FILLER_3_881 ();
 sg13g2_fill_1 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_932 ();
 sg13g2_decap_4 FILLER_3_939 ();
 sg13g2_fill_1 FILLER_3_981 ();
 sg13g2_fill_1 FILLER_3_988 ();
 sg13g2_fill_2 FILLER_3_1001 ();
 sg13g2_fill_1 FILLER_3_1003 ();
 sg13g2_fill_2 FILLER_3_1012 ();
 sg13g2_fill_1 FILLER_3_1014 ();
 sg13g2_fill_2 FILLER_3_1053 ();
 sg13g2_fill_2 FILLER_3_1081 ();
 sg13g2_fill_1 FILLER_3_1083 ();
 sg13g2_fill_1 FILLER_3_1092 ();
 sg13g2_decap_4 FILLER_3_1127 ();
 sg13g2_decap_4 FILLER_3_1165 ();
 sg13g2_decap_8 FILLER_3_1173 ();
 sg13g2_fill_1 FILLER_3_1184 ();
 sg13g2_decap_4 FILLER_3_1189 ();
 sg13g2_fill_1 FILLER_3_1193 ();
 sg13g2_decap_4 FILLER_3_1198 ();
 sg13g2_fill_2 FILLER_3_1206 ();
 sg13g2_fill_1 FILLER_3_1208 ();
 sg13g2_decap_4 FILLER_3_1213 ();
 sg13g2_fill_2 FILLER_3_1217 ();
 sg13g2_decap_8 FILLER_3_1275 ();
 sg13g2_fill_2 FILLER_3_1282 ();
 sg13g2_fill_1 FILLER_3_1284 ();
 sg13g2_fill_2 FILLER_3_1371 ();
 sg13g2_fill_2 FILLER_3_1377 ();
 sg13g2_fill_1 FILLER_3_1379 ();
 sg13g2_fill_2 FILLER_3_1386 ();
 sg13g2_fill_1 FILLER_3_1388 ();
 sg13g2_fill_2 FILLER_3_1393 ();
 sg13g2_fill_1 FILLER_3_1399 ();
 sg13g2_decap_8 FILLER_3_1404 ();
 sg13g2_fill_2 FILLER_3_1428 ();
 sg13g2_fill_2 FILLER_3_1446 ();
 sg13g2_fill_1 FILLER_3_1455 ();
 sg13g2_decap_8 FILLER_3_1466 ();
 sg13g2_decap_4 FILLER_3_1473 ();
 sg13g2_decap_8 FILLER_3_1480 ();
 sg13g2_fill_2 FILLER_3_1499 ();
 sg13g2_fill_1 FILLER_3_1506 ();
 sg13g2_fill_2 FILLER_3_1512 ();
 sg13g2_fill_1 FILLER_3_1518 ();
 sg13g2_decap_4 FILLER_3_1524 ();
 sg13g2_fill_2 FILLER_3_1528 ();
 sg13g2_decap_8 FILLER_3_1578 ();
 sg13g2_decap_4 FILLER_3_1585 ();
 sg13g2_fill_2 FILLER_3_1589 ();
 sg13g2_decap_4 FILLER_3_1596 ();
 sg13g2_fill_2 FILLER_3_1604 ();
 sg13g2_fill_1 FILLER_3_1606 ();
 sg13g2_fill_1 FILLER_3_1612 ();
 sg13g2_fill_1 FILLER_3_1639 ();
 sg13g2_fill_1 FILLER_3_1645 ();
 sg13g2_decap_8 FILLER_3_1650 ();
 sg13g2_fill_1 FILLER_3_1714 ();
 sg13g2_decap_4 FILLER_3_1750 ();
 sg13g2_decap_8 FILLER_3_1759 ();
 sg13g2_fill_2 FILLER_3_1771 ();
 sg13g2_decap_4 FILLER_3_1778 ();
 sg13g2_fill_2 FILLER_3_1782 ();
 sg13g2_fill_2 FILLER_3_1797 ();
 sg13g2_fill_1 FILLER_3_1799 ();
 sg13g2_fill_2 FILLER_3_1830 ();
 sg13g2_decap_8 FILLER_3_1863 ();
 sg13g2_fill_1 FILLER_3_1870 ();
 sg13g2_decap_8 FILLER_3_1902 ();
 sg13g2_fill_2 FILLER_3_1909 ();
 sg13g2_fill_1 FILLER_3_1911 ();
 sg13g2_fill_1 FILLER_3_1917 ();
 sg13g2_decap_4 FILLER_3_1928 ();
 sg13g2_fill_2 FILLER_3_1932 ();
 sg13g2_decap_4 FILLER_3_1942 ();
 sg13g2_fill_2 FILLER_3_1946 ();
 sg13g2_fill_1 FILLER_3_1953 ();
 sg13g2_fill_2 FILLER_3_1984 ();
 sg13g2_fill_1 FILLER_3_1986 ();
 sg13g2_fill_2 FILLER_3_2000 ();
 sg13g2_fill_1 FILLER_3_2002 ();
 sg13g2_fill_1 FILLER_3_2006 ();
 sg13g2_fill_2 FILLER_3_2033 ();
 sg13g2_fill_1 FILLER_3_2035 ();
 sg13g2_decap_4 FILLER_3_2054 ();
 sg13g2_fill_2 FILLER_3_2058 ();
 sg13g2_decap_8 FILLER_3_2095 ();
 sg13g2_decap_4 FILLER_3_2102 ();
 sg13g2_fill_2 FILLER_3_2106 ();
 sg13g2_fill_1 FILLER_3_2122 ();
 sg13g2_decap_4 FILLER_3_2128 ();
 sg13g2_fill_2 FILLER_3_2132 ();
 sg13g2_decap_8 FILLER_3_2147 ();
 sg13g2_decap_8 FILLER_3_2154 ();
 sg13g2_decap_8 FILLER_3_2161 ();
 sg13g2_decap_4 FILLER_3_2168 ();
 sg13g2_fill_2 FILLER_3_2172 ();
 sg13g2_decap_4 FILLER_3_2179 ();
 sg13g2_fill_1 FILLER_3_2183 ();
 sg13g2_decap_8 FILLER_3_2205 ();
 sg13g2_decap_8 FILLER_3_2238 ();
 sg13g2_decap_8 FILLER_3_2245 ();
 sg13g2_decap_8 FILLER_3_2252 ();
 sg13g2_fill_2 FILLER_3_2259 ();
 sg13g2_decap_8 FILLER_3_2269 ();
 sg13g2_fill_2 FILLER_3_2276 ();
 sg13g2_fill_1 FILLER_3_2278 ();
 sg13g2_fill_2 FILLER_3_2284 ();
 sg13g2_fill_1 FILLER_3_2286 ();
 sg13g2_decap_8 FILLER_3_2291 ();
 sg13g2_decap_8 FILLER_3_2298 ();
 sg13g2_decap_8 FILLER_3_2305 ();
 sg13g2_fill_2 FILLER_3_2312 ();
 sg13g2_fill_1 FILLER_3_2314 ();
 sg13g2_decap_4 FILLER_3_2320 ();
 sg13g2_fill_2 FILLER_3_2342 ();
 sg13g2_fill_1 FILLER_3_2349 ();
 sg13g2_decap_4 FILLER_3_2355 ();
 sg13g2_fill_2 FILLER_3_2359 ();
 sg13g2_fill_1 FILLER_3_2365 ();
 sg13g2_decap_8 FILLER_3_2371 ();
 sg13g2_decap_8 FILLER_3_2422 ();
 sg13g2_decap_8 FILLER_3_2429 ();
 sg13g2_decap_8 FILLER_3_2436 ();
 sg13g2_decap_8 FILLER_3_2443 ();
 sg13g2_decap_8 FILLER_3_2450 ();
 sg13g2_decap_8 FILLER_3_2457 ();
 sg13g2_decap_8 FILLER_3_2464 ();
 sg13g2_decap_8 FILLER_3_2471 ();
 sg13g2_decap_8 FILLER_3_2478 ();
 sg13g2_decap_8 FILLER_3_2485 ();
 sg13g2_decap_8 FILLER_3_2492 ();
 sg13g2_decap_8 FILLER_3_2499 ();
 sg13g2_decap_8 FILLER_3_2506 ();
 sg13g2_decap_8 FILLER_3_2513 ();
 sg13g2_decap_8 FILLER_3_2520 ();
 sg13g2_decap_8 FILLER_3_2527 ();
 sg13g2_decap_8 FILLER_3_2534 ();
 sg13g2_decap_8 FILLER_3_2541 ();
 sg13g2_decap_8 FILLER_3_2548 ();
 sg13g2_decap_8 FILLER_3_2555 ();
 sg13g2_decap_8 FILLER_3_2562 ();
 sg13g2_decap_8 FILLER_3_2569 ();
 sg13g2_decap_8 FILLER_3_2576 ();
 sg13g2_decap_8 FILLER_3_2583 ();
 sg13g2_decap_8 FILLER_3_2590 ();
 sg13g2_decap_8 FILLER_3_2597 ();
 sg13g2_decap_8 FILLER_3_2604 ();
 sg13g2_decap_8 FILLER_3_2611 ();
 sg13g2_decap_8 FILLER_3_2618 ();
 sg13g2_decap_8 FILLER_3_2625 ();
 sg13g2_decap_8 FILLER_3_2632 ();
 sg13g2_decap_8 FILLER_3_2639 ();
 sg13g2_decap_8 FILLER_3_2646 ();
 sg13g2_decap_8 FILLER_3_2653 ();
 sg13g2_decap_8 FILLER_3_2660 ();
 sg13g2_fill_2 FILLER_3_2667 ();
 sg13g2_fill_1 FILLER_3_2669 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_4 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_51 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_decap_4 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_188 ();
 sg13g2_decap_4 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_4 FILLER_4_232 ();
 sg13g2_decap_4 FILLER_4_246 ();
 sg13g2_fill_1 FILLER_4_250 ();
 sg13g2_fill_2 FILLER_4_272 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_fill_2 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_4 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_fill_1 FILLER_4_390 ();
 sg13g2_fill_1 FILLER_4_395 ();
 sg13g2_fill_2 FILLER_4_422 ();
 sg13g2_decap_8 FILLER_4_433 ();
 sg13g2_decap_4 FILLER_4_440 ();
 sg13g2_fill_2 FILLER_4_444 ();
 sg13g2_fill_1 FILLER_4_496 ();
 sg13g2_decap_8 FILLER_4_523 ();
 sg13g2_decap_8 FILLER_4_530 ();
 sg13g2_decap_8 FILLER_4_537 ();
 sg13g2_decap_8 FILLER_4_544 ();
 sg13g2_decap_8 FILLER_4_551 ();
 sg13g2_decap_8 FILLER_4_558 ();
 sg13g2_decap_4 FILLER_4_565 ();
 sg13g2_fill_2 FILLER_4_569 ();
 sg13g2_decap_8 FILLER_4_584 ();
 sg13g2_decap_8 FILLER_4_591 ();
 sg13g2_decap_8 FILLER_4_598 ();
 sg13g2_decap_4 FILLER_4_605 ();
 sg13g2_fill_2 FILLER_4_639 ();
 sg13g2_decap_4 FILLER_4_649 ();
 sg13g2_fill_1 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_667 ();
 sg13g2_decap_8 FILLER_4_674 ();
 sg13g2_decap_8 FILLER_4_681 ();
 sg13g2_fill_2 FILLER_4_688 ();
 sg13g2_fill_1 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_695 ();
 sg13g2_decap_4 FILLER_4_712 ();
 sg13g2_fill_2 FILLER_4_716 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_4 FILLER_4_735 ();
 sg13g2_fill_2 FILLER_4_739 ();
 sg13g2_fill_2 FILLER_4_745 ();
 sg13g2_fill_1 FILLER_4_747 ();
 sg13g2_fill_1 FILLER_4_773 ();
 sg13g2_fill_2 FILLER_4_783 ();
 sg13g2_fill_1 FILLER_4_794 ();
 sg13g2_fill_2 FILLER_4_799 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_fill_1 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_864 ();
 sg13g2_decap_8 FILLER_4_871 ();
 sg13g2_decap_8 FILLER_4_878 ();
 sg13g2_decap_8 FILLER_4_885 ();
 sg13g2_decap_8 FILLER_4_892 ();
 sg13g2_decap_8 FILLER_4_899 ();
 sg13g2_decap_8 FILLER_4_906 ();
 sg13g2_decap_8 FILLER_4_913 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_decap_4 FILLER_4_927 ();
 sg13g2_fill_1 FILLER_4_931 ();
 sg13g2_fill_1 FILLER_4_940 ();
 sg13g2_decap_8 FILLER_4_971 ();
 sg13g2_decap_4 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_988 ();
 sg13g2_decap_8 FILLER_4_995 ();
 sg13g2_decap_8 FILLER_4_1002 ();
 sg13g2_fill_2 FILLER_4_1009 ();
 sg13g2_fill_1 FILLER_4_1011 ();
 sg13g2_decap_8 FILLER_4_1051 ();
 sg13g2_decap_4 FILLER_4_1058 ();
 sg13g2_fill_2 FILLER_4_1062 ();
 sg13g2_decap_8 FILLER_4_1068 ();
 sg13g2_decap_4 FILLER_4_1079 ();
 sg13g2_fill_2 FILLER_4_1083 ();
 sg13g2_decap_8 FILLER_4_1089 ();
 sg13g2_decap_8 FILLER_4_1096 ();
 sg13g2_decap_8 FILLER_4_1115 ();
 sg13g2_decap_8 FILLER_4_1122 ();
 sg13g2_decap_8 FILLER_4_1129 ();
 sg13g2_decap_4 FILLER_4_1136 ();
 sg13g2_fill_2 FILLER_4_1140 ();
 sg13g2_decap_8 FILLER_4_1150 ();
 sg13g2_decap_4 FILLER_4_1157 ();
 sg13g2_fill_1 FILLER_4_1161 ();
 sg13g2_decap_8 FILLER_4_1192 ();
 sg13g2_decap_8 FILLER_4_1199 ();
 sg13g2_decap_8 FILLER_4_1206 ();
 sg13g2_fill_2 FILLER_4_1217 ();
 sg13g2_fill_2 FILLER_4_1245 ();
 sg13g2_fill_2 FILLER_4_1273 ();
 sg13g2_fill_1 FILLER_4_1275 ();
 sg13g2_decap_8 FILLER_4_1306 ();
 sg13g2_fill_2 FILLER_4_1313 ();
 sg13g2_fill_1 FILLER_4_1315 ();
 sg13g2_decap_4 FILLER_4_1320 ();
 sg13g2_fill_1 FILLER_4_1328 ();
 sg13g2_fill_2 FILLER_4_1346 ();
 sg13g2_fill_1 FILLER_4_1348 ();
 sg13g2_fill_1 FILLER_4_1353 ();
 sg13g2_decap_8 FILLER_4_1359 ();
 sg13g2_decap_8 FILLER_4_1366 ();
 sg13g2_decap_8 FILLER_4_1373 ();
 sg13g2_decap_8 FILLER_4_1380 ();
 sg13g2_decap_8 FILLER_4_1387 ();
 sg13g2_fill_1 FILLER_4_1426 ();
 sg13g2_decap_8 FILLER_4_1459 ();
 sg13g2_decap_8 FILLER_4_1466 ();
 sg13g2_decap_4 FILLER_4_1473 ();
 sg13g2_fill_1 FILLER_4_1486 ();
 sg13g2_fill_2 FILLER_4_1492 ();
 sg13g2_fill_1 FILLER_4_1494 ();
 sg13g2_fill_2 FILLER_4_1508 ();
 sg13g2_fill_1 FILLER_4_1519 ();
 sg13g2_decap_4 FILLER_4_1525 ();
 sg13g2_fill_1 FILLER_4_1529 ();
 sg13g2_fill_2 FILLER_4_1538 ();
 sg13g2_decap_4 FILLER_4_1570 ();
 sg13g2_decap_4 FILLER_4_1579 ();
 sg13g2_decap_8 FILLER_4_1591 ();
 sg13g2_decap_8 FILLER_4_1598 ();
 sg13g2_decap_4 FILLER_4_1605 ();
 sg13g2_decap_4 FILLER_4_1622 ();
 sg13g2_fill_1 FILLER_4_1630 ();
 sg13g2_decap_8 FILLER_4_1637 ();
 sg13g2_decap_8 FILLER_4_1644 ();
 sg13g2_fill_1 FILLER_4_1651 ();
 sg13g2_fill_2 FILLER_4_1665 ();
 sg13g2_fill_1 FILLER_4_1667 ();
 sg13g2_decap_4 FILLER_4_1679 ();
 sg13g2_decap_4 FILLER_4_1733 ();
 sg13g2_decap_8 FILLER_4_1741 ();
 sg13g2_decap_4 FILLER_4_1748 ();
 sg13g2_fill_1 FILLER_4_1752 ();
 sg13g2_fill_2 FILLER_4_1784 ();
 sg13g2_decap_8 FILLER_4_1795 ();
 sg13g2_decap_8 FILLER_4_1802 ();
 sg13g2_decap_8 FILLER_4_1809 ();
 sg13g2_decap_8 FILLER_4_1816 ();
 sg13g2_decap_8 FILLER_4_1823 ();
 sg13g2_decap_8 FILLER_4_1830 ();
 sg13g2_fill_1 FILLER_4_1837 ();
 sg13g2_decap_4 FILLER_4_1843 ();
 sg13g2_fill_2 FILLER_4_1847 ();
 sg13g2_fill_2 FILLER_4_1853 ();
 sg13g2_decap_8 FILLER_4_1859 ();
 sg13g2_decap_4 FILLER_4_1866 ();
 sg13g2_fill_2 FILLER_4_1879 ();
 sg13g2_fill_1 FILLER_4_1881 ();
 sg13g2_decap_4 FILLER_4_1900 ();
 sg13g2_fill_2 FILLER_4_1909 ();
 sg13g2_fill_1 FILLER_4_1911 ();
 sg13g2_fill_2 FILLER_4_1941 ();
 sg13g2_decap_8 FILLER_4_1948 ();
 sg13g2_fill_1 FILLER_4_1955 ();
 sg13g2_decap_8 FILLER_4_1960 ();
 sg13g2_fill_2 FILLER_4_1967 ();
 sg13g2_fill_1 FILLER_4_1995 ();
 sg13g2_fill_2 FILLER_4_1999 ();
 sg13g2_decap_4 FILLER_4_2030 ();
 sg13g2_fill_2 FILLER_4_2039 ();
 sg13g2_decap_8 FILLER_4_2049 ();
 sg13g2_fill_1 FILLER_4_2056 ();
 sg13g2_decap_4 FILLER_4_2062 ();
 sg13g2_fill_2 FILLER_4_2066 ();
 sg13g2_decap_8 FILLER_4_2105 ();
 sg13g2_decap_8 FILLER_4_2112 ();
 sg13g2_fill_1 FILLER_4_2119 ();
 sg13g2_decap_4 FILLER_4_2125 ();
 sg13g2_fill_1 FILLER_4_2129 ();
 sg13g2_fill_2 FILLER_4_2141 ();
 sg13g2_decap_8 FILLER_4_2178 ();
 sg13g2_fill_1 FILLER_4_2185 ();
 sg13g2_fill_1 FILLER_4_2189 ();
 sg13g2_decap_8 FILLER_4_2198 ();
 sg13g2_decap_4 FILLER_4_2205 ();
 sg13g2_fill_1 FILLER_4_2209 ();
 sg13g2_fill_1 FILLER_4_2220 ();
 sg13g2_decap_8 FILLER_4_2225 ();
 sg13g2_fill_1 FILLER_4_2232 ();
 sg13g2_fill_2 FILLER_4_2236 ();
 sg13g2_fill_2 FILLER_4_2243 ();
 sg13g2_decap_8 FILLER_4_2249 ();
 sg13g2_decap_4 FILLER_4_2256 ();
 sg13g2_fill_1 FILLER_4_2260 ();
 sg13g2_decap_8 FILLER_4_2267 ();
 sg13g2_fill_2 FILLER_4_2274 ();
 sg13g2_fill_1 FILLER_4_2276 ();
 sg13g2_decap_8 FILLER_4_2283 ();
 sg13g2_decap_8 FILLER_4_2290 ();
 sg13g2_decap_4 FILLER_4_2297 ();
 sg13g2_decap_8 FILLER_4_2314 ();
 sg13g2_fill_2 FILLER_4_2321 ();
 sg13g2_fill_1 FILLER_4_2323 ();
 sg13g2_decap_4 FILLER_4_2333 ();
 sg13g2_fill_2 FILLER_4_2337 ();
 sg13g2_decap_4 FILLER_4_2343 ();
 sg13g2_fill_1 FILLER_4_2347 ();
 sg13g2_decap_8 FILLER_4_2352 ();
 sg13g2_decap_8 FILLER_4_2359 ();
 sg13g2_decap_8 FILLER_4_2366 ();
 sg13g2_decap_8 FILLER_4_2373 ();
 sg13g2_decap_8 FILLER_4_2380 ();
 sg13g2_decap_8 FILLER_4_2387 ();
 sg13g2_decap_8 FILLER_4_2394 ();
 sg13g2_decap_8 FILLER_4_2401 ();
 sg13g2_decap_8 FILLER_4_2408 ();
 sg13g2_decap_8 FILLER_4_2415 ();
 sg13g2_decap_8 FILLER_4_2422 ();
 sg13g2_decap_8 FILLER_4_2429 ();
 sg13g2_decap_8 FILLER_4_2436 ();
 sg13g2_decap_8 FILLER_4_2443 ();
 sg13g2_decap_8 FILLER_4_2450 ();
 sg13g2_decap_8 FILLER_4_2457 ();
 sg13g2_decap_8 FILLER_4_2464 ();
 sg13g2_decap_8 FILLER_4_2471 ();
 sg13g2_decap_8 FILLER_4_2478 ();
 sg13g2_decap_8 FILLER_4_2485 ();
 sg13g2_decap_8 FILLER_4_2492 ();
 sg13g2_decap_8 FILLER_4_2499 ();
 sg13g2_decap_8 FILLER_4_2506 ();
 sg13g2_decap_8 FILLER_4_2513 ();
 sg13g2_decap_8 FILLER_4_2520 ();
 sg13g2_decap_8 FILLER_4_2527 ();
 sg13g2_decap_8 FILLER_4_2534 ();
 sg13g2_decap_8 FILLER_4_2541 ();
 sg13g2_decap_8 FILLER_4_2548 ();
 sg13g2_decap_8 FILLER_4_2555 ();
 sg13g2_decap_8 FILLER_4_2562 ();
 sg13g2_decap_8 FILLER_4_2569 ();
 sg13g2_decap_8 FILLER_4_2576 ();
 sg13g2_decap_8 FILLER_4_2583 ();
 sg13g2_decap_8 FILLER_4_2590 ();
 sg13g2_decap_8 FILLER_4_2597 ();
 sg13g2_decap_8 FILLER_4_2604 ();
 sg13g2_decap_8 FILLER_4_2611 ();
 sg13g2_decap_8 FILLER_4_2618 ();
 sg13g2_decap_8 FILLER_4_2625 ();
 sg13g2_decap_8 FILLER_4_2632 ();
 sg13g2_decap_8 FILLER_4_2639 ();
 sg13g2_decap_8 FILLER_4_2646 ();
 sg13g2_decap_8 FILLER_4_2653 ();
 sg13g2_decap_8 FILLER_4_2660 ();
 sg13g2_fill_2 FILLER_4_2667 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_23 ();
 sg13g2_decap_4 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_48 ();
 sg13g2_decap_4 FILLER_5_55 ();
 sg13g2_decap_8 FILLER_5_78 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_4 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_113 ();
 sg13g2_fill_1 FILLER_5_120 ();
 sg13g2_fill_2 FILLER_5_127 ();
 sg13g2_decap_8 FILLER_5_159 ();
 sg13g2_decap_8 FILLER_5_166 ();
 sg13g2_decap_8 FILLER_5_173 ();
 sg13g2_decap_4 FILLER_5_180 ();
 sg13g2_fill_2 FILLER_5_212 ();
 sg13g2_fill_2 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_decap_4 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_decap_4 FILLER_5_254 ();
 sg13g2_fill_1 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_367 ();
 sg13g2_fill_2 FILLER_5_378 ();
 sg13g2_decap_4 FILLER_5_385 ();
 sg13g2_fill_1 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_5_435 ();
 sg13g2_decap_8 FILLER_5_442 ();
 sg13g2_fill_2 FILLER_5_449 ();
 sg13g2_fill_1 FILLER_5_451 ();
 sg13g2_decap_4 FILLER_5_456 ();
 sg13g2_decap_4 FILLER_5_498 ();
 sg13g2_fill_2 FILLER_5_502 ();
 sg13g2_decap_8 FILLER_5_530 ();
 sg13g2_decap_8 FILLER_5_537 ();
 sg13g2_decap_8 FILLER_5_544 ();
 sg13g2_decap_8 FILLER_5_551 ();
 sg13g2_decap_8 FILLER_5_562 ();
 sg13g2_fill_2 FILLER_5_569 ();
 sg13g2_fill_1 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_580 ();
 sg13g2_decap_8 FILLER_5_587 ();
 sg13g2_decap_8 FILLER_5_594 ();
 sg13g2_decap_8 FILLER_5_601 ();
 sg13g2_fill_1 FILLER_5_608 ();
 sg13g2_fill_1 FILLER_5_639 ();
 sg13g2_fill_2 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_678 ();
 sg13g2_decap_8 FILLER_5_685 ();
 sg13g2_fill_2 FILLER_5_692 ();
 sg13g2_fill_1 FILLER_5_694 ();
 sg13g2_decap_8 FILLER_5_734 ();
 sg13g2_fill_2 FILLER_5_741 ();
 sg13g2_fill_2 FILLER_5_824 ();
 sg13g2_fill_1 FILLER_5_826 ();
 sg13g2_decap_4 FILLER_5_887 ();
 sg13g2_decap_8 FILLER_5_934 ();
 sg13g2_decap_4 FILLER_5_941 ();
 sg13g2_fill_1 FILLER_5_945 ();
 sg13g2_decap_8 FILLER_5_950 ();
 sg13g2_fill_2 FILLER_5_988 ();
 sg13g2_decap_8 FILLER_5_1046 ();
 sg13g2_decap_8 FILLER_5_1053 ();
 sg13g2_decap_8 FILLER_5_1060 ();
 sg13g2_decap_8 FILLER_5_1067 ();
 sg13g2_decap_8 FILLER_5_1074 ();
 sg13g2_decap_8 FILLER_5_1081 ();
 sg13g2_decap_8 FILLER_5_1088 ();
 sg13g2_decap_8 FILLER_5_1095 ();
 sg13g2_decap_8 FILLER_5_1102 ();
 sg13g2_decap_8 FILLER_5_1109 ();
 sg13g2_decap_8 FILLER_5_1116 ();
 sg13g2_decap_8 FILLER_5_1123 ();
 sg13g2_decap_8 FILLER_5_1130 ();
 sg13g2_decap_8 FILLER_5_1137 ();
 sg13g2_decap_8 FILLER_5_1144 ();
 sg13g2_decap_8 FILLER_5_1151 ();
 sg13g2_decap_8 FILLER_5_1158 ();
 sg13g2_fill_2 FILLER_5_1165 ();
 sg13g2_decap_8 FILLER_5_1201 ();
 sg13g2_decap_8 FILLER_5_1212 ();
 sg13g2_fill_2 FILLER_5_1223 ();
 sg13g2_fill_1 FILLER_5_1225 ();
 sg13g2_fill_2 FILLER_5_1230 ();
 sg13g2_fill_1 FILLER_5_1232 ();
 sg13g2_decap_8 FILLER_5_1237 ();
 sg13g2_fill_2 FILLER_5_1244 ();
 sg13g2_fill_1 FILLER_5_1246 ();
 sg13g2_fill_1 FILLER_5_1255 ();
 sg13g2_fill_1 FILLER_5_1260 ();
 sg13g2_fill_1 FILLER_5_1291 ();
 sg13g2_decap_4 FILLER_5_1296 ();
 sg13g2_fill_2 FILLER_5_1300 ();
 sg13g2_fill_2 FILLER_5_1306 ();
 sg13g2_fill_2 FILLER_5_1334 ();
 sg13g2_fill_1 FILLER_5_1336 ();
 sg13g2_decap_4 FILLER_5_1367 ();
 sg13g2_fill_2 FILLER_5_1375 ();
 sg13g2_fill_1 FILLER_5_1407 ();
 sg13g2_fill_2 FILLER_5_1424 ();
 sg13g2_decap_8 FILLER_5_1486 ();
 sg13g2_fill_2 FILLER_5_1493 ();
 sg13g2_decap_4 FILLER_5_1508 ();
 sg13g2_fill_2 FILLER_5_1525 ();
 sg13g2_decap_4 FILLER_5_1540 ();
 sg13g2_fill_2 FILLER_5_1544 ();
 sg13g2_decap_4 FILLER_5_1551 ();
 sg13g2_fill_2 FILLER_5_1555 ();
 sg13g2_fill_2 FILLER_5_1560 ();
 sg13g2_decap_4 FILLER_5_1568 ();
 sg13g2_decap_8 FILLER_5_1624 ();
 sg13g2_decap_8 FILLER_5_1631 ();
 sg13g2_fill_2 FILLER_5_1638 ();
 sg13g2_fill_2 FILLER_5_1671 ();
 sg13g2_fill_1 FILLER_5_1673 ();
 sg13g2_fill_2 FILLER_5_1695 ();
 sg13g2_fill_1 FILLER_5_1705 ();
 sg13g2_decap_8 FILLER_5_1710 ();
 sg13g2_fill_1 FILLER_5_1717 ();
 sg13g2_decap_8 FILLER_5_1723 ();
 sg13g2_fill_1 FILLER_5_1730 ();
 sg13g2_fill_1 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1744 ();
 sg13g2_decap_8 FILLER_5_1751 ();
 sg13g2_decap_8 FILLER_5_1758 ();
 sg13g2_fill_1 FILLER_5_1765 ();
 sg13g2_decap_8 FILLER_5_1770 ();
 sg13g2_decap_8 FILLER_5_1777 ();
 sg13g2_decap_8 FILLER_5_1784 ();
 sg13g2_decap_4 FILLER_5_1791 ();
 sg13g2_decap_8 FILLER_5_1801 ();
 sg13g2_decap_8 FILLER_5_1808 ();
 sg13g2_decap_8 FILLER_5_1815 ();
 sg13g2_decap_8 FILLER_5_1822 ();
 sg13g2_decap_8 FILLER_5_1829 ();
 sg13g2_fill_1 FILLER_5_1836 ();
 sg13g2_decap_4 FILLER_5_1842 ();
 sg13g2_decap_8 FILLER_5_1860 ();
 sg13g2_fill_1 FILLER_5_1867 ();
 sg13g2_fill_2 FILLER_5_1894 ();
 sg13g2_decap_4 FILLER_5_1901 ();
 sg13g2_decap_8 FILLER_5_1969 ();
 sg13g2_decap_4 FILLER_5_1976 ();
 sg13g2_fill_2 FILLER_5_1980 ();
 sg13g2_fill_1 FILLER_5_1992 ();
 sg13g2_fill_1 FILLER_5_2015 ();
 sg13g2_fill_2 FILLER_5_2021 ();
 sg13g2_fill_1 FILLER_5_2023 ();
 sg13g2_fill_2 FILLER_5_2032 ();
 sg13g2_fill_1 FILLER_5_2038 ();
 sg13g2_decap_8 FILLER_5_2091 ();
 sg13g2_decap_8 FILLER_5_2098 ();
 sg13g2_decap_8 FILLER_5_2105 ();
 sg13g2_decap_8 FILLER_5_2112 ();
 sg13g2_fill_1 FILLER_5_2119 ();
 sg13g2_decap_8 FILLER_5_2146 ();
 sg13g2_decap_4 FILLER_5_2153 ();
 sg13g2_decap_8 FILLER_5_2162 ();
 sg13g2_fill_2 FILLER_5_2169 ();
 sg13g2_decap_4 FILLER_5_2227 ();
 sg13g2_fill_2 FILLER_5_2231 ();
 sg13g2_fill_2 FILLER_5_2239 ();
 sg13g2_fill_2 FILLER_5_2267 ();
 sg13g2_fill_1 FILLER_5_2269 ();
 sg13g2_decap_8 FILLER_5_2278 ();
 sg13g2_fill_2 FILLER_5_2285 ();
 sg13g2_fill_2 FILLER_5_2292 ();
 sg13g2_decap_4 FILLER_5_2320 ();
 sg13g2_fill_2 FILLER_5_2324 ();
 sg13g2_decap_8 FILLER_5_2339 ();
 sg13g2_decap_8 FILLER_5_2346 ();
 sg13g2_decap_4 FILLER_5_2353 ();
 sg13g2_fill_2 FILLER_5_2371 ();
 sg13g2_fill_1 FILLER_5_2373 ();
 sg13g2_decap_8 FILLER_5_2380 ();
 sg13g2_decap_8 FILLER_5_2387 ();
 sg13g2_decap_8 FILLER_5_2407 ();
 sg13g2_decap_8 FILLER_5_2414 ();
 sg13g2_decap_8 FILLER_5_2421 ();
 sg13g2_decap_8 FILLER_5_2441 ();
 sg13g2_decap_8 FILLER_5_2448 ();
 sg13g2_decap_8 FILLER_5_2455 ();
 sg13g2_decap_8 FILLER_5_2462 ();
 sg13g2_decap_8 FILLER_5_2469 ();
 sg13g2_decap_8 FILLER_5_2476 ();
 sg13g2_decap_8 FILLER_5_2483 ();
 sg13g2_decap_8 FILLER_5_2490 ();
 sg13g2_decap_8 FILLER_5_2497 ();
 sg13g2_decap_8 FILLER_5_2504 ();
 sg13g2_decap_8 FILLER_5_2511 ();
 sg13g2_decap_8 FILLER_5_2518 ();
 sg13g2_decap_8 FILLER_5_2525 ();
 sg13g2_decap_8 FILLER_5_2532 ();
 sg13g2_decap_8 FILLER_5_2539 ();
 sg13g2_decap_8 FILLER_5_2546 ();
 sg13g2_decap_8 FILLER_5_2553 ();
 sg13g2_decap_8 FILLER_5_2560 ();
 sg13g2_decap_8 FILLER_5_2567 ();
 sg13g2_decap_8 FILLER_5_2574 ();
 sg13g2_decap_8 FILLER_5_2581 ();
 sg13g2_decap_8 FILLER_5_2588 ();
 sg13g2_decap_8 FILLER_5_2595 ();
 sg13g2_decap_8 FILLER_5_2602 ();
 sg13g2_decap_8 FILLER_5_2609 ();
 sg13g2_decap_8 FILLER_5_2616 ();
 sg13g2_decap_8 FILLER_5_2623 ();
 sg13g2_decap_8 FILLER_5_2630 ();
 sg13g2_decap_8 FILLER_5_2637 ();
 sg13g2_decap_8 FILLER_5_2644 ();
 sg13g2_decap_8 FILLER_5_2651 ();
 sg13g2_decap_8 FILLER_5_2658 ();
 sg13g2_decap_4 FILLER_5_2665 ();
 sg13g2_fill_1 FILLER_5_2669 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_4 ();
 sg13g2_fill_2 FILLER_6_47 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_4 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_182 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_230 ();
 sg13g2_decap_8 FILLER_6_237 ();
 sg13g2_decap_4 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_4 FILLER_6_398 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_fill_2 FILLER_6_448 ();
 sg13g2_fill_2 FILLER_6_454 ();
 sg13g2_fill_1 FILLER_6_480 ();
 sg13g2_fill_1 FILLER_6_494 ();
 sg13g2_decap_4 FILLER_6_499 ();
 sg13g2_fill_2 FILLER_6_503 ();
 sg13g2_fill_1 FILLER_6_535 ();
 sg13g2_fill_1 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_598 ();
 sg13g2_fill_2 FILLER_6_605 ();
 sg13g2_fill_1 FILLER_6_607 ();
 sg13g2_decap_4 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_621 ();
 sg13g2_decap_8 FILLER_6_628 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_decap_8 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_fill_2 FILLER_6_697 ();
 sg13g2_fill_1 FILLER_6_733 ();
 sg13g2_fill_2 FILLER_6_738 ();
 sg13g2_fill_1 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_fill_1 FILLER_6_839 ();
 sg13g2_fill_2 FILLER_6_849 ();
 sg13g2_fill_1 FILLER_6_851 ();
 sg13g2_fill_2 FILLER_6_860 ();
 sg13g2_fill_1 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_898 ();
 sg13g2_decap_4 FILLER_6_905 ();
 sg13g2_fill_2 FILLER_6_909 ();
 sg13g2_decap_8 FILLER_6_915 ();
 sg13g2_fill_2 FILLER_6_922 ();
 sg13g2_fill_1 FILLER_6_924 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_4 FILLER_6_942 ();
 sg13g2_fill_1 FILLER_6_946 ();
 sg13g2_decap_8 FILLER_6_976 ();
 sg13g2_decap_8 FILLER_6_983 ();
 sg13g2_decap_8 FILLER_6_994 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_fill_1 FILLER_6_1008 ();
 sg13g2_decap_4 FILLER_6_1018 ();
 sg13g2_fill_1 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1049 ();
 sg13g2_decap_4 FILLER_6_1056 ();
 sg13g2_fill_1 FILLER_6_1060 ();
 sg13g2_decap_8 FILLER_6_1087 ();
 sg13g2_decap_8 FILLER_6_1094 ();
 sg13g2_fill_2 FILLER_6_1101 ();
 sg13g2_fill_1 FILLER_6_1103 ();
 sg13g2_decap_8 FILLER_6_1140 ();
 sg13g2_decap_8 FILLER_6_1147 ();
 sg13g2_fill_2 FILLER_6_1154 ();
 sg13g2_decap_8 FILLER_6_1162 ();
 sg13g2_decap_8 FILLER_6_1169 ();
 sg13g2_decap_4 FILLER_6_1176 ();
 sg13g2_fill_2 FILLER_6_1180 ();
 sg13g2_decap_8 FILLER_6_1186 ();
 sg13g2_decap_4 FILLER_6_1193 ();
 sg13g2_fill_1 FILLER_6_1197 ();
 sg13g2_decap_8 FILLER_6_1241 ();
 sg13g2_decap_8 FILLER_6_1248 ();
 sg13g2_decap_8 FILLER_6_1255 ();
 sg13g2_decap_8 FILLER_6_1262 ();
 sg13g2_decap_4 FILLER_6_1269 ();
 sg13g2_decap_8 FILLER_6_1281 ();
 sg13g2_decap_8 FILLER_6_1288 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_decap_8 FILLER_6_1302 ();
 sg13g2_decap_8 FILLER_6_1309 ();
 sg13g2_decap_8 FILLER_6_1320 ();
 sg13g2_decap_8 FILLER_6_1327 ();
 sg13g2_decap_8 FILLER_6_1334 ();
 sg13g2_decap_8 FILLER_6_1394 ();
 sg13g2_decap_8 FILLER_6_1401 ();
 sg13g2_decap_8 FILLER_6_1408 ();
 sg13g2_fill_2 FILLER_6_1415 ();
 sg13g2_fill_2 FILLER_6_1420 ();
 sg13g2_fill_1 FILLER_6_1422 ();
 sg13g2_fill_2 FILLER_6_1466 ();
 sg13g2_fill_1 FILLER_6_1468 ();
 sg13g2_fill_1 FILLER_6_1499 ();
 sg13g2_fill_1 FILLER_6_1504 ();
 sg13g2_decap_8 FILLER_6_1509 ();
 sg13g2_decap_8 FILLER_6_1516 ();
 sg13g2_decap_8 FILLER_6_1523 ();
 sg13g2_decap_8 FILLER_6_1530 ();
 sg13g2_fill_2 FILLER_6_1537 ();
 sg13g2_decap_8 FILLER_6_1544 ();
 sg13g2_fill_2 FILLER_6_1551 ();
 sg13g2_fill_1 FILLER_6_1561 ();
 sg13g2_fill_1 FILLER_6_1565 ();
 sg13g2_fill_2 FILLER_6_1596 ();
 sg13g2_fill_1 FILLER_6_1598 ();
 sg13g2_decap_8 FILLER_6_1607 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_fill_1 FILLER_6_1625 ();
 sg13g2_decap_8 FILLER_6_1684 ();
 sg13g2_fill_1 FILLER_6_1696 ();
 sg13g2_decap_8 FILLER_6_1703 ();
 sg13g2_fill_1 FILLER_6_1740 ();
 sg13g2_fill_2 FILLER_6_1748 ();
 sg13g2_fill_1 FILLER_6_1750 ();
 sg13g2_decap_8 FILLER_6_1812 ();
 sg13g2_fill_1 FILLER_6_1819 ();
 sg13g2_fill_1 FILLER_6_1826 ();
 sg13g2_decap_8 FILLER_6_2011 ();
 sg13g2_fill_2 FILLER_6_2018 ();
 sg13g2_fill_1 FILLER_6_2020 ();
 sg13g2_decap_8 FILLER_6_2033 ();
 sg13g2_fill_2 FILLER_6_2040 ();
 sg13g2_fill_1 FILLER_6_2047 ();
 sg13g2_decap_4 FILLER_6_2052 ();
 sg13g2_fill_2 FILLER_6_2056 ();
 sg13g2_fill_1 FILLER_6_2061 ();
 sg13g2_decap_8 FILLER_6_2071 ();
 sg13g2_decap_8 FILLER_6_2078 ();
 sg13g2_decap_8 FILLER_6_2085 ();
 sg13g2_decap_8 FILLER_6_2092 ();
 sg13g2_fill_2 FILLER_6_2099 ();
 sg13g2_fill_1 FILLER_6_2101 ();
 sg13g2_fill_1 FILLER_6_2107 ();
 sg13g2_fill_2 FILLER_6_2158 ();
 sg13g2_fill_1 FILLER_6_2160 ();
 sg13g2_decap_4 FILLER_6_2169 ();
 sg13g2_fill_2 FILLER_6_2187 ();
 sg13g2_decap_8 FILLER_6_2255 ();
 sg13g2_decap_8 FILLER_6_2262 ();
 sg13g2_fill_2 FILLER_6_2290 ();
 sg13g2_fill_1 FILLER_6_2292 ();
 sg13g2_decap_4 FILLER_6_2350 ();
 sg13g2_fill_1 FILLER_6_2354 ();
 sg13g2_fill_2 FILLER_6_2358 ();
 sg13g2_fill_1 FILLER_6_2368 ();
 sg13g2_fill_1 FILLER_6_2425 ();
 sg13g2_decap_8 FILLER_6_2452 ();
 sg13g2_decap_8 FILLER_6_2459 ();
 sg13g2_decap_8 FILLER_6_2466 ();
 sg13g2_decap_8 FILLER_6_2473 ();
 sg13g2_decap_8 FILLER_6_2480 ();
 sg13g2_decap_8 FILLER_6_2487 ();
 sg13g2_decap_8 FILLER_6_2494 ();
 sg13g2_decap_8 FILLER_6_2501 ();
 sg13g2_decap_8 FILLER_6_2508 ();
 sg13g2_decap_8 FILLER_6_2515 ();
 sg13g2_decap_8 FILLER_6_2522 ();
 sg13g2_decap_8 FILLER_6_2529 ();
 sg13g2_decap_8 FILLER_6_2536 ();
 sg13g2_decap_8 FILLER_6_2543 ();
 sg13g2_decap_8 FILLER_6_2550 ();
 sg13g2_decap_8 FILLER_6_2557 ();
 sg13g2_decap_8 FILLER_6_2564 ();
 sg13g2_decap_8 FILLER_6_2571 ();
 sg13g2_decap_8 FILLER_6_2578 ();
 sg13g2_decap_8 FILLER_6_2585 ();
 sg13g2_decap_8 FILLER_6_2592 ();
 sg13g2_decap_8 FILLER_6_2599 ();
 sg13g2_decap_8 FILLER_6_2606 ();
 sg13g2_decap_8 FILLER_6_2613 ();
 sg13g2_decap_8 FILLER_6_2620 ();
 sg13g2_decap_8 FILLER_6_2627 ();
 sg13g2_decap_8 FILLER_6_2634 ();
 sg13g2_decap_8 FILLER_6_2641 ();
 sg13g2_decap_8 FILLER_6_2648 ();
 sg13g2_decap_8 FILLER_6_2655 ();
 sg13g2_decap_8 FILLER_6_2662 ();
 sg13g2_fill_1 FILLER_6_2669 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_50 ();
 sg13g2_decap_8 FILLER_7_86 ();
 sg13g2_decap_8 FILLER_7_93 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_decap_4 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_fill_1 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_4 FILLER_7_238 ();
 sg13g2_fill_1 FILLER_7_242 ();
 sg13g2_fill_2 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_4 FILLER_7_400 ();
 sg13g2_fill_1 FILLER_7_415 ();
 sg13g2_fill_2 FILLER_7_456 ();
 sg13g2_fill_1 FILLER_7_463 ();
 sg13g2_fill_1 FILLER_7_482 ();
 sg13g2_fill_2 FILLER_7_492 ();
 sg13g2_decap_8 FILLER_7_498 ();
 sg13g2_decap_8 FILLER_7_505 ();
 sg13g2_decap_4 FILLER_7_538 ();
 sg13g2_fill_1 FILLER_7_542 ();
 sg13g2_fill_1 FILLER_7_547 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_4 FILLER_7_560 ();
 sg13g2_fill_1 FILLER_7_568 ();
 sg13g2_fill_1 FILLER_7_604 ();
 sg13g2_fill_2 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_645 ();
 sg13g2_decap_4 FILLER_7_652 ();
 sg13g2_decap_8 FILLER_7_664 ();
 sg13g2_decap_8 FILLER_7_671 ();
 sg13g2_decap_8 FILLER_7_678 ();
 sg13g2_fill_1 FILLER_7_685 ();
 sg13g2_fill_2 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_fill_2 FILLER_7_777 ();
 sg13g2_fill_1 FILLER_7_779 ();
 sg13g2_fill_2 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_decap_8 FILLER_7_860 ();
 sg13g2_decap_4 FILLER_7_867 ();
 sg13g2_fill_2 FILLER_7_871 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_4 FILLER_7_887 ();
 sg13g2_fill_2 FILLER_7_891 ();
 sg13g2_decap_8 FILLER_7_897 ();
 sg13g2_decap_8 FILLER_7_904 ();
 sg13g2_decap_4 FILLER_7_911 ();
 sg13g2_fill_2 FILLER_7_915 ();
 sg13g2_fill_2 FILLER_7_923 ();
 sg13g2_fill_2 FILLER_7_976 ();
 sg13g2_fill_2 FILLER_7_981 ();
 sg13g2_fill_1 FILLER_7_983 ();
 sg13g2_fill_1 FILLER_7_1013 ();
 sg13g2_decap_4 FILLER_7_1019 ();
 sg13g2_fill_1 FILLER_7_1023 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_7_1034 ();
 sg13g2_decap_8 FILLER_7_1041 ();
 sg13g2_decap_8 FILLER_7_1048 ();
 sg13g2_decap_4 FILLER_7_1055 ();
 sg13g2_fill_1 FILLER_7_1059 ();
 sg13g2_decap_8 FILLER_7_1065 ();
 sg13g2_decap_4 FILLER_7_1072 ();
 sg13g2_fill_1 FILLER_7_1076 ();
 sg13g2_decap_4 FILLER_7_1103 ();
 sg13g2_fill_1 FILLER_7_1107 ();
 sg13g2_decap_8 FILLER_7_1118 ();
 sg13g2_fill_1 FILLER_7_1125 ();
 sg13g2_decap_4 FILLER_7_1152 ();
 sg13g2_fill_2 FILLER_7_1182 ();
 sg13g2_decap_8 FILLER_7_1190 ();
 sg13g2_decap_4 FILLER_7_1197 ();
 sg13g2_fill_2 FILLER_7_1201 ();
 sg13g2_decap_8 FILLER_7_1229 ();
 sg13g2_decap_8 FILLER_7_1236 ();
 sg13g2_decap_8 FILLER_7_1243 ();
 sg13g2_decap_8 FILLER_7_1250 ();
 sg13g2_fill_1 FILLER_7_1268 ();
 sg13g2_decap_8 FILLER_7_1274 ();
 sg13g2_decap_4 FILLER_7_1281 ();
 sg13g2_fill_1 FILLER_7_1285 ();
 sg13g2_fill_2 FILLER_7_1304 ();
 sg13g2_decap_4 FILLER_7_1332 ();
 sg13g2_fill_1 FILLER_7_1367 ();
 sg13g2_decap_8 FILLER_7_1394 ();
 sg13g2_decap_8 FILLER_7_1401 ();
 sg13g2_decap_8 FILLER_7_1408 ();
 sg13g2_decap_4 FILLER_7_1415 ();
 sg13g2_fill_1 FILLER_7_1419 ();
 sg13g2_decap_8 FILLER_7_1446 ();
 sg13g2_decap_4 FILLER_7_1462 ();
 sg13g2_fill_1 FILLER_7_1466 ();
 sg13g2_fill_1 FILLER_7_1471 ();
 sg13g2_fill_2 FILLER_7_1492 ();
 sg13g2_fill_1 FILLER_7_1494 ();
 sg13g2_decap_8 FILLER_7_1499 ();
 sg13g2_decap_8 FILLER_7_1506 ();
 sg13g2_decap_8 FILLER_7_1513 ();
 sg13g2_decap_8 FILLER_7_1520 ();
 sg13g2_decap_4 FILLER_7_1527 ();
 sg13g2_decap_8 FILLER_7_1566 ();
 sg13g2_fill_2 FILLER_7_1573 ();
 sg13g2_fill_1 FILLER_7_1575 ();
 sg13g2_decap_4 FILLER_7_1581 ();
 sg13g2_fill_1 FILLER_7_1585 ();
 sg13g2_fill_2 FILLER_7_1589 ();
 sg13g2_fill_1 FILLER_7_1591 ();
 sg13g2_fill_2 FILLER_7_1597 ();
 sg13g2_fill_1 FILLER_7_1599 ();
 sg13g2_fill_1 FILLER_7_1606 ();
 sg13g2_fill_2 FILLER_7_1612 ();
 sg13g2_fill_2 FILLER_7_1640 ();
 sg13g2_fill_1 FILLER_7_1656 ();
 sg13g2_fill_2 FILLER_7_1661 ();
 sg13g2_decap_4 FILLER_7_1689 ();
 sg13g2_decap_8 FILLER_7_1719 ();
 sg13g2_decap_8 FILLER_7_1726 ();
 sg13g2_fill_1 FILLER_7_1733 ();
 sg13g2_fill_1 FILLER_7_1739 ();
 sg13g2_fill_2 FILLER_7_1751 ();
 sg13g2_decap_8 FILLER_7_1784 ();
 sg13g2_decap_4 FILLER_7_1791 ();
 sg13g2_fill_2 FILLER_7_1795 ();
 sg13g2_fill_2 FILLER_7_1826 ();
 sg13g2_fill_1 FILLER_7_1828 ();
 sg13g2_fill_1 FILLER_7_1872 ();
 sg13g2_fill_1 FILLER_7_1879 ();
 sg13g2_fill_2 FILLER_7_1908 ();
 sg13g2_fill_1 FILLER_7_1916 ();
 sg13g2_fill_1 FILLER_7_1954 ();
 sg13g2_fill_2 FILLER_7_1977 ();
 sg13g2_fill_1 FILLER_7_1979 ();
 sg13g2_decap_8 FILLER_7_2040 ();
 sg13g2_decap_4 FILLER_7_2047 ();
 sg13g2_fill_1 FILLER_7_2051 ();
 sg13g2_decap_8 FILLER_7_2064 ();
 sg13g2_fill_2 FILLER_7_2071 ();
 sg13g2_fill_1 FILLER_7_2073 ();
 sg13g2_fill_1 FILLER_7_2079 ();
 sg13g2_fill_2 FILLER_7_2106 ();
 sg13g2_fill_1 FILLER_7_2141 ();
 sg13g2_fill_2 FILLER_7_2173 ();
 sg13g2_fill_2 FILLER_7_2181 ();
 sg13g2_decap_4 FILLER_7_2196 ();
 sg13g2_fill_1 FILLER_7_2200 ();
 sg13g2_decap_8 FILLER_7_2205 ();
 sg13g2_decap_8 FILLER_7_2212 ();
 sg13g2_fill_2 FILLER_7_2219 ();
 sg13g2_fill_1 FILLER_7_2221 ();
 sg13g2_decap_4 FILLER_7_2252 ();
 sg13g2_fill_2 FILLER_7_2256 ();
 sg13g2_fill_1 FILLER_7_2301 ();
 sg13g2_fill_1 FILLER_7_2333 ();
 sg13g2_fill_1 FILLER_7_2360 ();
 sg13g2_fill_1 FILLER_7_2367 ();
 sg13g2_fill_2 FILLER_7_2420 ();
 sg13g2_decap_8 FILLER_7_2458 ();
 sg13g2_decap_8 FILLER_7_2465 ();
 sg13g2_decap_8 FILLER_7_2472 ();
 sg13g2_decap_8 FILLER_7_2479 ();
 sg13g2_decap_8 FILLER_7_2486 ();
 sg13g2_decap_8 FILLER_7_2493 ();
 sg13g2_decap_8 FILLER_7_2500 ();
 sg13g2_decap_8 FILLER_7_2507 ();
 sg13g2_decap_8 FILLER_7_2514 ();
 sg13g2_decap_8 FILLER_7_2521 ();
 sg13g2_decap_8 FILLER_7_2528 ();
 sg13g2_decap_8 FILLER_7_2535 ();
 sg13g2_decap_8 FILLER_7_2542 ();
 sg13g2_decap_8 FILLER_7_2549 ();
 sg13g2_decap_8 FILLER_7_2556 ();
 sg13g2_decap_8 FILLER_7_2563 ();
 sg13g2_decap_8 FILLER_7_2570 ();
 sg13g2_decap_8 FILLER_7_2577 ();
 sg13g2_decap_8 FILLER_7_2584 ();
 sg13g2_decap_8 FILLER_7_2591 ();
 sg13g2_decap_8 FILLER_7_2598 ();
 sg13g2_decap_8 FILLER_7_2605 ();
 sg13g2_decap_8 FILLER_7_2612 ();
 sg13g2_decap_8 FILLER_7_2619 ();
 sg13g2_decap_8 FILLER_7_2626 ();
 sg13g2_decap_8 FILLER_7_2633 ();
 sg13g2_decap_8 FILLER_7_2640 ();
 sg13g2_decap_8 FILLER_7_2647 ();
 sg13g2_decap_8 FILLER_7_2654 ();
 sg13g2_decap_8 FILLER_7_2661 ();
 sg13g2_fill_2 FILLER_7_2668 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_11 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_fill_1 FILLER_8_55 ();
 sg13g2_fill_1 FILLER_8_69 ();
 sg13g2_decap_8 FILLER_8_82 ();
 sg13g2_fill_2 FILLER_8_89 ();
 sg13g2_fill_1 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_fill_2 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_142 ();
 sg13g2_decap_4 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_174 ();
 sg13g2_fill_2 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_222 ();
 sg13g2_decap_8 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_236 ();
 sg13g2_decap_8 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_250 ();
 sg13g2_decap_8 FILLER_8_257 ();
 sg13g2_fill_2 FILLER_8_264 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_1 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_decap_4 FILLER_8_364 ();
 sg13g2_fill_2 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_fill_1 FILLER_8_459 ();
 sg13g2_fill_2 FILLER_8_464 ();
 sg13g2_decap_8 FILLER_8_524 ();
 sg13g2_decap_8 FILLER_8_535 ();
 sg13g2_decap_8 FILLER_8_542 ();
 sg13g2_fill_1 FILLER_8_554 ();
 sg13g2_decap_8 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_597 ();
 sg13g2_decap_8 FILLER_8_647 ();
 sg13g2_decap_4 FILLER_8_654 ();
 sg13g2_fill_1 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_663 ();
 sg13g2_decap_4 FILLER_8_670 ();
 sg13g2_fill_1 FILLER_8_674 ();
 sg13g2_fill_2 FILLER_8_679 ();
 sg13g2_fill_1 FILLER_8_681 ();
 sg13g2_fill_1 FILLER_8_708 ();
 sg13g2_fill_1 FILLER_8_719 ();
 sg13g2_decap_8 FILLER_8_755 ();
 sg13g2_decap_4 FILLER_8_762 ();
 sg13g2_fill_1 FILLER_8_766 ();
 sg13g2_fill_1 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_4 FILLER_8_814 ();
 sg13g2_fill_1 FILLER_8_818 ();
 sg13g2_fill_2 FILLER_8_822 ();
 sg13g2_fill_2 FILLER_8_893 ();
 sg13g2_fill_2 FILLER_8_959 ();
 sg13g2_fill_1 FILLER_8_966 ();
 sg13g2_fill_1 FILLER_8_971 ();
 sg13g2_fill_2 FILLER_8_976 ();
 sg13g2_fill_1 FILLER_8_989 ();
 sg13g2_decap_4 FILLER_8_1016 ();
 sg13g2_fill_2 FILLER_8_1020 ();
 sg13g2_fill_1 FILLER_8_1027 ();
 sg13g2_fill_2 FILLER_8_1032 ();
 sg13g2_fill_1 FILLER_8_1060 ();
 sg13g2_fill_2 FILLER_8_1070 ();
 sg13g2_decap_4 FILLER_8_1104 ();
 sg13g2_fill_2 FILLER_8_1108 ();
 sg13g2_decap_8 FILLER_8_1140 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_4 FILLER_8_1246 ();
 sg13g2_fill_2 FILLER_8_1250 ();
 sg13g2_fill_2 FILLER_8_1260 ();
 sg13g2_fill_1 FILLER_8_1262 ();
 sg13g2_fill_2 FILLER_8_1323 ();
 sg13g2_fill_1 FILLER_8_1366 ();
 sg13g2_decap_4 FILLER_8_1403 ();
 sg13g2_fill_1 FILLER_8_1407 ();
 sg13g2_decap_8 FILLER_8_1416 ();
 sg13g2_decap_8 FILLER_8_1423 ();
 sg13g2_fill_1 FILLER_8_1430 ();
 sg13g2_fill_2 FILLER_8_1458 ();
 sg13g2_decap_4 FILLER_8_1469 ();
 sg13g2_fill_2 FILLER_8_1473 ();
 sg13g2_decap_8 FILLER_8_1488 ();
 sg13g2_decap_8 FILLER_8_1495 ();
 sg13g2_decap_8 FILLER_8_1502 ();
 sg13g2_decap_4 FILLER_8_1509 ();
 sg13g2_fill_1 FILLER_8_1513 ();
 sg13g2_decap_4 FILLER_8_1518 ();
 sg13g2_fill_2 FILLER_8_1522 ();
 sg13g2_fill_2 FILLER_8_1550 ();
 sg13g2_fill_2 FILLER_8_1592 ();
 sg13g2_fill_1 FILLER_8_1594 ();
 sg13g2_fill_2 FILLER_8_1616 ();
 sg13g2_fill_1 FILLER_8_1618 ();
 sg13g2_fill_2 FILLER_8_1624 ();
 sg13g2_fill_1 FILLER_8_1626 ();
 sg13g2_fill_2 FILLER_8_1649 ();
 sg13g2_fill_1 FILLER_8_1651 ();
 sg13g2_fill_1 FILLER_8_1657 ();
 sg13g2_decap_8 FILLER_8_1662 ();
 sg13g2_decap_4 FILLER_8_1669 ();
 sg13g2_decap_8 FILLER_8_1676 ();
 sg13g2_decap_4 FILLER_8_1683 ();
 sg13g2_fill_2 FILLER_8_1687 ();
 sg13g2_decap_4 FILLER_8_1698 ();
 sg13g2_decap_8 FILLER_8_1708 ();
 sg13g2_decap_8 FILLER_8_1715 ();
 sg13g2_decap_8 FILLER_8_1722 ();
 sg13g2_fill_2 FILLER_8_1729 ();
 sg13g2_decap_4 FILLER_8_1763 ();
 sg13g2_fill_1 FILLER_8_1767 ();
 sg13g2_fill_2 FILLER_8_1788 ();
 sg13g2_fill_1 FILLER_8_1790 ();
 sg13g2_fill_1 FILLER_8_1803 ();
 sg13g2_decap_8 FILLER_8_1834 ();
 sg13g2_decap_8 FILLER_8_1841 ();
 sg13g2_decap_4 FILLER_8_1848 ();
 sg13g2_fill_2 FILLER_8_1852 ();
 sg13g2_fill_2 FILLER_8_1857 ();
 sg13g2_fill_1 FILLER_8_1859 ();
 sg13g2_fill_1 FILLER_8_1924 ();
 sg13g2_decap_4 FILLER_8_1957 ();
 sg13g2_decap_4 FILLER_8_1965 ();
 sg13g2_fill_1 FILLER_8_1969 ();
 sg13g2_decap_4 FILLER_8_1975 ();
 sg13g2_fill_2 FILLER_8_1979 ();
 sg13g2_fill_1 FILLER_8_1993 ();
 sg13g2_decap_8 FILLER_8_2006 ();
 sg13g2_fill_2 FILLER_8_2013 ();
 sg13g2_fill_2 FILLER_8_2020 ();
 sg13g2_fill_2 FILLER_8_2026 ();
 sg13g2_fill_1 FILLER_8_2054 ();
 sg13g2_fill_1 FILLER_8_2058 ();
 sg13g2_decap_8 FILLER_8_2071 ();
 sg13g2_fill_2 FILLER_8_2078 ();
 sg13g2_fill_1 FILLER_8_2080 ();
 sg13g2_fill_1 FILLER_8_2123 ();
 sg13g2_fill_2 FILLER_8_2141 ();
 sg13g2_decap_8 FILLER_8_2149 ();
 sg13g2_decap_8 FILLER_8_2156 ();
 sg13g2_decap_4 FILLER_8_2169 ();
 sg13g2_fill_2 FILLER_8_2189 ();
 sg13g2_fill_1 FILLER_8_2196 ();
 sg13g2_fill_1 FILLER_8_2223 ();
 sg13g2_fill_1 FILLER_8_2229 ();
 sg13g2_fill_1 FILLER_8_2234 ();
 sg13g2_fill_1 FILLER_8_2239 ();
 sg13g2_fill_1 FILLER_8_2246 ();
 sg13g2_fill_1 FILLER_8_2278 ();
 sg13g2_fill_2 FILLER_8_2294 ();
 sg13g2_fill_1 FILLER_8_2296 ();
 sg13g2_fill_2 FILLER_8_2302 ();
 sg13g2_fill_1 FILLER_8_2304 ();
 sg13g2_decap_8 FILLER_8_2309 ();
 sg13g2_fill_1 FILLER_8_2316 ();
 sg13g2_fill_2 FILLER_8_2326 ();
 sg13g2_decap_8 FILLER_8_2463 ();
 sg13g2_decap_8 FILLER_8_2470 ();
 sg13g2_decap_8 FILLER_8_2477 ();
 sg13g2_decap_8 FILLER_8_2484 ();
 sg13g2_decap_8 FILLER_8_2491 ();
 sg13g2_decap_8 FILLER_8_2498 ();
 sg13g2_decap_8 FILLER_8_2505 ();
 sg13g2_decap_8 FILLER_8_2512 ();
 sg13g2_decap_8 FILLER_8_2519 ();
 sg13g2_decap_8 FILLER_8_2526 ();
 sg13g2_decap_8 FILLER_8_2533 ();
 sg13g2_decap_8 FILLER_8_2540 ();
 sg13g2_decap_8 FILLER_8_2547 ();
 sg13g2_decap_8 FILLER_8_2554 ();
 sg13g2_decap_8 FILLER_8_2561 ();
 sg13g2_decap_8 FILLER_8_2568 ();
 sg13g2_decap_8 FILLER_8_2575 ();
 sg13g2_decap_8 FILLER_8_2582 ();
 sg13g2_decap_8 FILLER_8_2589 ();
 sg13g2_decap_8 FILLER_8_2596 ();
 sg13g2_decap_8 FILLER_8_2603 ();
 sg13g2_decap_8 FILLER_8_2610 ();
 sg13g2_decap_8 FILLER_8_2617 ();
 sg13g2_decap_8 FILLER_8_2624 ();
 sg13g2_decap_8 FILLER_8_2631 ();
 sg13g2_decap_8 FILLER_8_2638 ();
 sg13g2_decap_8 FILLER_8_2645 ();
 sg13g2_decap_8 FILLER_8_2652 ();
 sg13g2_decap_8 FILLER_8_2659 ();
 sg13g2_decap_4 FILLER_8_2666 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_85 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_101 ();
 sg13g2_fill_2 FILLER_9_114 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_4 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_fill_1 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_4 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_221 ();
 sg13g2_decap_4 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_fill_1 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_4 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_fill_1 FILLER_9_414 ();
 sg13g2_fill_2 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_433 ();
 sg13g2_fill_1 FILLER_9_435 ();
 sg13g2_decap_4 FILLER_9_441 ();
 sg13g2_fill_2 FILLER_9_445 ();
 sg13g2_fill_1 FILLER_9_473 ();
 sg13g2_fill_1 FILLER_9_478 ();
 sg13g2_fill_2 FILLER_9_487 ();
 sg13g2_fill_2 FILLER_9_515 ();
 sg13g2_fill_2 FILLER_9_522 ();
 sg13g2_fill_1 FILLER_9_555 ();
 sg13g2_fill_1 FILLER_9_586 ();
 sg13g2_decap_8 FILLER_9_591 ();
 sg13g2_decap_4 FILLER_9_598 ();
 sg13g2_fill_2 FILLER_9_610 ();
 sg13g2_fill_1 FILLER_9_612 ();
 sg13g2_fill_2 FILLER_9_643 ();
 sg13g2_fill_1 FILLER_9_645 ();
 sg13g2_decap_4 FILLER_9_682 ();
 sg13g2_fill_1 FILLER_9_686 ();
 sg13g2_fill_2 FILLER_9_691 ();
 sg13g2_decap_8 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_704 ();
 sg13g2_decap_8 FILLER_9_711 ();
 sg13g2_fill_2 FILLER_9_718 ();
 sg13g2_fill_2 FILLER_9_723 ();
 sg13g2_fill_2 FILLER_9_768 ();
 sg13g2_fill_1 FILLER_9_770 ();
 sg13g2_decap_4 FILLER_9_775 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_4 FILLER_9_791 ();
 sg13g2_fill_2 FILLER_9_795 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_fill_1 FILLER_9_815 ();
 sg13g2_fill_2 FILLER_9_824 ();
 sg13g2_decap_4 FILLER_9_863 ();
 sg13g2_fill_2 FILLER_9_867 ();
 sg13g2_decap_8 FILLER_9_874 ();
 sg13g2_decap_4 FILLER_9_881 ();
 sg13g2_fill_2 FILLER_9_889 ();
 sg13g2_fill_2 FILLER_9_931 ();
 sg13g2_fill_2 FILLER_9_974 ();
 sg13g2_fill_2 FILLER_9_984 ();
 sg13g2_decap_8 FILLER_9_1004 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_fill_1 FILLER_9_1029 ();
 sg13g2_decap_8 FILLER_9_1040 ();
 sg13g2_decap_8 FILLER_9_1047 ();
 sg13g2_decap_8 FILLER_9_1054 ();
 sg13g2_decap_4 FILLER_9_1061 ();
 sg13g2_fill_2 FILLER_9_1065 ();
 sg13g2_decap_4 FILLER_9_1115 ();
 sg13g2_fill_1 FILLER_9_1119 ();
 sg13g2_decap_4 FILLER_9_1129 ();
 sg13g2_decap_8 FILLER_9_1168 ();
 sg13g2_decap_4 FILLER_9_1175 ();
 sg13g2_fill_1 FILLER_9_1179 ();
 sg13g2_fill_1 FILLER_9_1193 ();
 sg13g2_fill_2 FILLER_9_1210 ();
 sg13g2_fill_1 FILLER_9_1212 ();
 sg13g2_fill_2 FILLER_9_1226 ();
 sg13g2_decap_4 FILLER_9_1263 ();
 sg13g2_fill_2 FILLER_9_1267 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_fill_2 FILLER_9_1285 ();
 sg13g2_fill_1 FILLER_9_1287 ();
 sg13g2_decap_8 FILLER_9_1299 ();
 sg13g2_decap_8 FILLER_9_1306 ();
 sg13g2_decap_8 FILLER_9_1313 ();
 sg13g2_decap_8 FILLER_9_1320 ();
 sg13g2_decap_8 FILLER_9_1327 ();
 sg13g2_decap_8 FILLER_9_1334 ();
 sg13g2_decap_8 FILLER_9_1341 ();
 sg13g2_fill_2 FILLER_9_1348 ();
 sg13g2_fill_1 FILLER_9_1378 ();
 sg13g2_fill_1 FILLER_9_1430 ();
 sg13g2_fill_1 FILLER_9_1449 ();
 sg13g2_decap_8 FILLER_9_1489 ();
 sg13g2_decap_8 FILLER_9_1500 ();
 sg13g2_decap_4 FILLER_9_1507 ();
 sg13g2_decap_8 FILLER_9_1545 ();
 sg13g2_fill_2 FILLER_9_1552 ();
 sg13g2_decap_8 FILLER_9_1559 ();
 sg13g2_fill_2 FILLER_9_1566 ();
 sg13g2_decap_8 FILLER_9_1573 ();
 sg13g2_fill_1 FILLER_9_1580 ();
 sg13g2_fill_1 FILLER_9_1585 ();
 sg13g2_fill_1 FILLER_9_1589 ();
 sg13g2_fill_2 FILLER_9_1597 ();
 sg13g2_decap_8 FILLER_9_1654 ();
 sg13g2_fill_2 FILLER_9_1670 ();
 sg13g2_fill_1 FILLER_9_1672 ();
 sg13g2_decap_4 FILLER_9_1679 ();
 sg13g2_fill_1 FILLER_9_1687 ();
 sg13g2_decap_8 FILLER_9_1719 ();
 sg13g2_decap_8 FILLER_9_1726 ();
 sg13g2_decap_8 FILLER_9_1733 ();
 sg13g2_fill_2 FILLER_9_1740 ();
 sg13g2_decap_4 FILLER_9_1747 ();
 sg13g2_fill_1 FILLER_9_1751 ();
 sg13g2_fill_2 FILLER_9_1756 ();
 sg13g2_fill_1 FILLER_9_1758 ();
 sg13g2_fill_1 FILLER_9_1765 ();
 sg13g2_fill_2 FILLER_9_1770 ();
 sg13g2_fill_1 FILLER_9_1772 ();
 sg13g2_fill_2 FILLER_9_1799 ();
 sg13g2_fill_1 FILLER_9_1801 ();
 sg13g2_fill_1 FILLER_9_1823 ();
 sg13g2_decap_4 FILLER_9_1850 ();
 sg13g2_fill_1 FILLER_9_1869 ();
 sg13g2_fill_1 FILLER_9_1951 ();
 sg13g2_decap_8 FILLER_9_1986 ();
 sg13g2_decap_4 FILLER_9_1993 ();
 sg13g2_fill_1 FILLER_9_1997 ();
 sg13g2_fill_2 FILLER_9_2021 ();
 sg13g2_decap_4 FILLER_9_2028 ();
 sg13g2_fill_2 FILLER_9_2040 ();
 sg13g2_decap_4 FILLER_9_2047 ();
 sg13g2_decap_8 FILLER_9_2065 ();
 sg13g2_fill_1 FILLER_9_2072 ();
 sg13g2_fill_1 FILLER_9_2078 ();
 sg13g2_fill_2 FILLER_9_2096 ();
 sg13g2_fill_1 FILLER_9_2098 ();
 sg13g2_fill_2 FILLER_9_2114 ();
 sg13g2_decap_4 FILLER_9_2213 ();
 sg13g2_fill_2 FILLER_9_2217 ();
 sg13g2_decap_8 FILLER_9_2230 ();
 sg13g2_fill_2 FILLER_9_2237 ();
 sg13g2_fill_1 FILLER_9_2262 ();
 sg13g2_decap_4 FILLER_9_2269 ();
 sg13g2_decap_8 FILLER_9_2293 ();
 sg13g2_decap_8 FILLER_9_2300 ();
 sg13g2_decap_8 FILLER_9_2307 ();
 sg13g2_decap_8 FILLER_9_2314 ();
 sg13g2_decap_8 FILLER_9_2321 ();
 sg13g2_fill_1 FILLER_9_2328 ();
 sg13g2_fill_1 FILLER_9_2345 ();
 sg13g2_fill_2 FILLER_9_2358 ();
 sg13g2_fill_2 FILLER_9_2380 ();
 sg13g2_fill_1 FILLER_9_2390 ();
 sg13g2_decap_8 FILLER_9_2486 ();
 sg13g2_decap_8 FILLER_9_2493 ();
 sg13g2_decap_8 FILLER_9_2500 ();
 sg13g2_decap_8 FILLER_9_2507 ();
 sg13g2_decap_8 FILLER_9_2514 ();
 sg13g2_decap_8 FILLER_9_2521 ();
 sg13g2_decap_8 FILLER_9_2528 ();
 sg13g2_decap_8 FILLER_9_2535 ();
 sg13g2_decap_8 FILLER_9_2542 ();
 sg13g2_decap_8 FILLER_9_2549 ();
 sg13g2_decap_8 FILLER_9_2556 ();
 sg13g2_decap_8 FILLER_9_2563 ();
 sg13g2_decap_8 FILLER_9_2570 ();
 sg13g2_decap_8 FILLER_9_2577 ();
 sg13g2_decap_8 FILLER_9_2584 ();
 sg13g2_decap_8 FILLER_9_2591 ();
 sg13g2_decap_8 FILLER_9_2598 ();
 sg13g2_decap_8 FILLER_9_2605 ();
 sg13g2_decap_8 FILLER_9_2612 ();
 sg13g2_decap_8 FILLER_9_2619 ();
 sg13g2_decap_8 FILLER_9_2626 ();
 sg13g2_decap_8 FILLER_9_2633 ();
 sg13g2_decap_8 FILLER_9_2640 ();
 sg13g2_decap_8 FILLER_9_2647 ();
 sg13g2_decap_8 FILLER_9_2654 ();
 sg13g2_decap_8 FILLER_9_2661 ();
 sg13g2_fill_2 FILLER_9_2668 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_17 ();
 sg13g2_fill_1 FILLER_10_24 ();
 sg13g2_decap_8 FILLER_10_33 ();
 sg13g2_decap_8 FILLER_10_40 ();
 sg13g2_decap_8 FILLER_10_47 ();
 sg13g2_decap_4 FILLER_10_54 ();
 sg13g2_fill_2 FILLER_10_58 ();
 sg13g2_decap_8 FILLER_10_64 ();
 sg13g2_decap_8 FILLER_10_71 ();
 sg13g2_decap_8 FILLER_10_78 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_4 FILLER_10_92 ();
 sg13g2_fill_1 FILLER_10_129 ();
 sg13g2_decap_8 FILLER_10_134 ();
 sg13g2_decap_8 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_148 ();
 sg13g2_decap_8 FILLER_10_157 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_178 ();
 sg13g2_decap_8 FILLER_10_185 ();
 sg13g2_decap_8 FILLER_10_192 ();
 sg13g2_decap_8 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_4 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_4 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_298 ();
 sg13g2_decap_4 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_decap_4 FILLER_10_323 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_4 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_4 FILLER_10_385 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_fill_2 FILLER_10_395 ();
 sg13g2_fill_1 FILLER_10_397 ();
 sg13g2_fill_2 FILLER_10_412 ();
 sg13g2_fill_2 FILLER_10_420 ();
 sg13g2_fill_1 FILLER_10_435 ();
 sg13g2_decap_8 FILLER_10_449 ();
 sg13g2_decap_4 FILLER_10_456 ();
 sg13g2_decap_8 FILLER_10_465 ();
 sg13g2_decap_8 FILLER_10_472 ();
 sg13g2_decap_8 FILLER_10_479 ();
 sg13g2_decap_8 FILLER_10_486 ();
 sg13g2_decap_8 FILLER_10_493 ();
 sg13g2_decap_4 FILLER_10_500 ();
 sg13g2_fill_1 FILLER_10_504 ();
 sg13g2_fill_1 FILLER_10_510 ();
 sg13g2_fill_1 FILLER_10_515 ();
 sg13g2_fill_1 FILLER_10_521 ();
 sg13g2_fill_1 FILLER_10_526 ();
 sg13g2_fill_1 FILLER_10_532 ();
 sg13g2_fill_1 FILLER_10_537 ();
 sg13g2_decap_8 FILLER_10_542 ();
 sg13g2_decap_4 FILLER_10_549 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_fill_2 FILLER_10_603 ();
 sg13g2_fill_2 FILLER_10_608 ();
 sg13g2_decap_4 FILLER_10_615 ();
 sg13g2_fill_2 FILLER_10_661 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_4 FILLER_10_674 ();
 sg13g2_decap_4 FILLER_10_687 ();
 sg13g2_decap_8 FILLER_10_717 ();
 sg13g2_decap_4 FILLER_10_733 ();
 sg13g2_fill_2 FILLER_10_737 ();
 sg13g2_fill_2 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_4 FILLER_10_784 ();
 sg13g2_fill_1 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_fill_2 FILLER_10_826 ();
 sg13g2_decap_4 FILLER_10_838 ();
 sg13g2_decap_8 FILLER_10_855 ();
 sg13g2_fill_1 FILLER_10_905 ();
 sg13g2_fill_1 FILLER_10_916 ();
 sg13g2_fill_2 FILLER_10_960 ();
 sg13g2_fill_2 FILLER_10_995 ();
 sg13g2_fill_2 FILLER_10_1003 ();
 sg13g2_decap_4 FILLER_10_1011 ();
 sg13g2_fill_2 FILLER_10_1015 ();
 sg13g2_fill_1 FILLER_10_1049 ();
 sg13g2_fill_1 FILLER_10_1062 ();
 sg13g2_fill_2 FILLER_10_1067 ();
 sg13g2_fill_1 FILLER_10_1077 ();
 sg13g2_decap_8 FILLER_10_1133 ();
 sg13g2_decap_8 FILLER_10_1144 ();
 sg13g2_fill_2 FILLER_10_1151 ();
 sg13g2_fill_1 FILLER_10_1153 ();
 sg13g2_fill_2 FILLER_10_1159 ();
 sg13g2_fill_2 FILLER_10_1165 ();
 sg13g2_fill_1 FILLER_10_1167 ();
 sg13g2_fill_2 FILLER_10_1203 ();
 sg13g2_decap_4 FILLER_10_1217 ();
 sg13g2_fill_1 FILLER_10_1221 ();
 sg13g2_decap_4 FILLER_10_1226 ();
 sg13g2_decap_4 FILLER_10_1242 ();
 sg13g2_decap_8 FILLER_10_1256 ();
 sg13g2_decap_4 FILLER_10_1263 ();
 sg13g2_fill_1 FILLER_10_1267 ();
 sg13g2_fill_1 FILLER_10_1300 ();
 sg13g2_decap_4 FILLER_10_1310 ();
 sg13g2_fill_1 FILLER_10_1314 ();
 sg13g2_fill_1 FILLER_10_1324 ();
 sg13g2_decap_4 FILLER_10_1351 ();
 sg13g2_fill_2 FILLER_10_1366 ();
 sg13g2_decap_4 FILLER_10_1392 ();
 sg13g2_fill_1 FILLER_10_1396 ();
 sg13g2_fill_2 FILLER_10_1432 ();
 sg13g2_decap_4 FILLER_10_1463 ();
 sg13g2_decap_8 FILLER_10_1498 ();
 sg13g2_decap_4 FILLER_10_1509 ();
 sg13g2_decap_4 FILLER_10_1523 ();
 sg13g2_fill_1 FILLER_10_1527 ();
 sg13g2_fill_1 FILLER_10_1537 ();
 sg13g2_decap_4 FILLER_10_1542 ();
 sg13g2_fill_1 FILLER_10_1552 ();
 sg13g2_decap_8 FILLER_10_1579 ();
 sg13g2_fill_1 FILLER_10_1586 ();
 sg13g2_decap_8 FILLER_10_1592 ();
 sg13g2_fill_2 FILLER_10_1614 ();
 sg13g2_fill_1 FILLER_10_1633 ();
 sg13g2_fill_2 FILLER_10_1639 ();
 sg13g2_fill_1 FILLER_10_1645 ();
 sg13g2_decap_8 FILLER_10_1678 ();
 sg13g2_fill_1 FILLER_10_1685 ();
 sg13g2_decap_8 FILLER_10_1724 ();
 sg13g2_decap_8 FILLER_10_1731 ();
 sg13g2_decap_4 FILLER_10_1738 ();
 sg13g2_fill_2 FILLER_10_1742 ();
 sg13g2_fill_2 FILLER_10_1749 ();
 sg13g2_fill_1 FILLER_10_1751 ();
 sg13g2_decap_8 FILLER_10_1795 ();
 sg13g2_decap_8 FILLER_10_1802 ();
 sg13g2_decap_4 FILLER_10_1814 ();
 sg13g2_fill_1 FILLER_10_1818 ();
 sg13g2_fill_1 FILLER_10_1824 ();
 sg13g2_fill_2 FILLER_10_1834 ();
 sg13g2_fill_2 FILLER_10_1840 ();
 sg13g2_fill_1 FILLER_10_1846 ();
 sg13g2_fill_2 FILLER_10_1855 ();
 sg13g2_decap_4 FILLER_10_1866 ();
 sg13g2_fill_2 FILLER_10_1870 ();
 sg13g2_fill_2 FILLER_10_1938 ();
 sg13g2_fill_1 FILLER_10_1940 ();
 sg13g2_decap_4 FILLER_10_1967 ();
 sg13g2_fill_2 FILLER_10_1981 ();
 sg13g2_fill_1 FILLER_10_1983 ();
 sg13g2_decap_4 FILLER_10_2048 ();
 sg13g2_fill_1 FILLER_10_2052 ();
 sg13g2_fill_2 FILLER_10_2057 ();
 sg13g2_decap_4 FILLER_10_2088 ();
 sg13g2_fill_1 FILLER_10_2092 ();
 sg13g2_fill_1 FILLER_10_2133 ();
 sg13g2_fill_1 FILLER_10_2138 ();
 sg13g2_fill_2 FILLER_10_2146 ();
 sg13g2_fill_1 FILLER_10_2153 ();
 sg13g2_fill_2 FILLER_10_2172 ();
 sg13g2_fill_2 FILLER_10_2226 ();
 sg13g2_fill_2 FILLER_10_2257 ();
 sg13g2_fill_1 FILLER_10_2259 ();
 sg13g2_decap_8 FILLER_10_2298 ();
 sg13g2_fill_2 FILLER_10_2305 ();
 sg13g2_fill_1 FILLER_10_2345 ();
 sg13g2_fill_1 FILLER_10_2364 ();
 sg13g2_fill_1 FILLER_10_2369 ();
 sg13g2_fill_1 FILLER_10_2411 ();
 sg13g2_fill_1 FILLER_10_2436 ();
 sg13g2_decap_8 FILLER_10_2486 ();
 sg13g2_decap_8 FILLER_10_2493 ();
 sg13g2_decap_8 FILLER_10_2500 ();
 sg13g2_decap_8 FILLER_10_2507 ();
 sg13g2_decap_8 FILLER_10_2514 ();
 sg13g2_decap_8 FILLER_10_2521 ();
 sg13g2_decap_8 FILLER_10_2528 ();
 sg13g2_decap_8 FILLER_10_2535 ();
 sg13g2_decap_8 FILLER_10_2542 ();
 sg13g2_decap_8 FILLER_10_2549 ();
 sg13g2_decap_8 FILLER_10_2556 ();
 sg13g2_decap_8 FILLER_10_2563 ();
 sg13g2_decap_8 FILLER_10_2570 ();
 sg13g2_decap_8 FILLER_10_2577 ();
 sg13g2_decap_8 FILLER_10_2584 ();
 sg13g2_decap_8 FILLER_10_2591 ();
 sg13g2_decap_8 FILLER_10_2598 ();
 sg13g2_decap_8 FILLER_10_2605 ();
 sg13g2_decap_8 FILLER_10_2612 ();
 sg13g2_decap_8 FILLER_10_2619 ();
 sg13g2_decap_8 FILLER_10_2626 ();
 sg13g2_decap_8 FILLER_10_2633 ();
 sg13g2_decap_8 FILLER_10_2640 ();
 sg13g2_decap_8 FILLER_10_2647 ();
 sg13g2_decap_8 FILLER_10_2654 ();
 sg13g2_decap_8 FILLER_10_2661 ();
 sg13g2_fill_2 FILLER_10_2668 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_1 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_50 ();
 sg13g2_decap_8 FILLER_11_57 ();
 sg13g2_decap_8 FILLER_11_64 ();
 sg13g2_decap_8 FILLER_11_71 ();
 sg13g2_decap_4 FILLER_11_78 ();
 sg13g2_decap_4 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_123 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_fill_2 FILLER_11_179 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_208 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_fill_1 FILLER_11_254 ();
 sg13g2_fill_2 FILLER_11_289 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_4 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_fill_2 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_374 ();
 sg13g2_fill_1 FILLER_11_379 ();
 sg13g2_fill_1 FILLER_11_386 ();
 sg13g2_decap_4 FILLER_11_398 ();
 sg13g2_fill_1 FILLER_11_428 ();
 sg13g2_fill_2 FILLER_11_447 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_4 FILLER_11_476 ();
 sg13g2_fill_2 FILLER_11_480 ();
 sg13g2_decap_4 FILLER_11_486 ();
 sg13g2_decap_4 FILLER_11_520 ();
 sg13g2_fill_1 FILLER_11_534 ();
 sg13g2_fill_1 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_556 ();
 sg13g2_decap_8 FILLER_11_563 ();
 sg13g2_decap_8 FILLER_11_570 ();
 sg13g2_decap_8 FILLER_11_577 ();
 sg13g2_decap_4 FILLER_11_584 ();
 sg13g2_fill_2 FILLER_11_588 ();
 sg13g2_fill_2 FILLER_11_614 ();
 sg13g2_decap_8 FILLER_11_625 ();
 sg13g2_decap_4 FILLER_11_632 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_4 FILLER_11_647 ();
 sg13g2_fill_2 FILLER_11_687 ();
 sg13g2_fill_1 FILLER_11_689 ();
 sg13g2_fill_2 FILLER_11_748 ();
 sg13g2_decap_8 FILLER_11_758 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_fill_2 FILLER_11_780 ();
 sg13g2_fill_1 FILLER_11_814 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_4 FILLER_11_858 ();
 sg13g2_fill_1 FILLER_11_862 ();
 sg13g2_fill_2 FILLER_11_868 ();
 sg13g2_fill_1 FILLER_11_878 ();
 sg13g2_fill_1 FILLER_11_897 ();
 sg13g2_fill_1 FILLER_11_911 ();
 sg13g2_fill_2 FILLER_11_941 ();
 sg13g2_fill_2 FILLER_11_979 ();
 sg13g2_decap_8 FILLER_11_993 ();
 sg13g2_fill_2 FILLER_11_1000 ();
 sg13g2_fill_1 FILLER_11_1008 ();
 sg13g2_fill_2 FILLER_11_1109 ();
 sg13g2_decap_8 FILLER_11_1143 ();
 sg13g2_decap_4 FILLER_11_1150 ();
 sg13g2_fill_1 FILLER_11_1154 ();
 sg13g2_fill_1 FILLER_11_1177 ();
 sg13g2_fill_2 FILLER_11_1183 ();
 sg13g2_fill_1 FILLER_11_1231 ();
 sg13g2_fill_2 FILLER_11_1258 ();
 sg13g2_decap_8 FILLER_11_1266 ();
 sg13g2_decap_4 FILLER_11_1273 ();
 sg13g2_decap_4 FILLER_11_1287 ();
 sg13g2_fill_2 FILLER_11_1291 ();
 sg13g2_decap_8 FILLER_11_1327 ();
 sg13g2_decap_4 FILLER_11_1334 ();
 sg13g2_fill_2 FILLER_11_1338 ();
 sg13g2_fill_1 FILLER_11_1345 ();
 sg13g2_decap_8 FILLER_11_1350 ();
 sg13g2_fill_2 FILLER_11_1377 ();
 sg13g2_fill_2 FILLER_11_1387 ();
 sg13g2_decap_4 FILLER_11_1396 ();
 sg13g2_fill_1 FILLER_11_1400 ();
 sg13g2_fill_1 FILLER_11_1410 ();
 sg13g2_fill_1 FILLER_11_1418 ();
 sg13g2_decap_8 FILLER_11_1440 ();
 sg13g2_decap_4 FILLER_11_1447 ();
 sg13g2_fill_2 FILLER_11_1451 ();
 sg13g2_fill_1 FILLER_11_1482 ();
 sg13g2_fill_1 FILLER_11_1510 ();
 sg13g2_decap_8 FILLER_11_1516 ();
 sg13g2_decap_4 FILLER_11_1523 ();
 sg13g2_fill_1 FILLER_11_1527 ();
 sg13g2_decap_8 FILLER_11_1531 ();
 sg13g2_decap_4 FILLER_11_1538 ();
 sg13g2_fill_2 FILLER_11_1547 ();
 sg13g2_fill_1 FILLER_11_1579 ();
 sg13g2_decap_4 FILLER_11_1585 ();
 sg13g2_fill_1 FILLER_11_1598 ();
 sg13g2_fill_2 FILLER_11_1616 ();
 sg13g2_fill_2 FILLER_11_1631 ();
 sg13g2_fill_2 FILLER_11_1664 ();
 sg13g2_fill_1 FILLER_11_1666 ();
 sg13g2_decap_8 FILLER_11_1673 ();
 sg13g2_decap_8 FILLER_11_1733 ();
 sg13g2_decap_8 FILLER_11_1740 ();
 sg13g2_decap_8 FILLER_11_1747 ();
 sg13g2_decap_4 FILLER_11_1754 ();
 sg13g2_decap_4 FILLER_11_1789 ();
 sg13g2_fill_2 FILLER_11_1828 ();
 sg13g2_fill_1 FILLER_11_1830 ();
 sg13g2_decap_8 FILLER_11_1868 ();
 sg13g2_decap_8 FILLER_11_1933 ();
 sg13g2_fill_2 FILLER_11_1940 ();
 sg13g2_fill_1 FILLER_11_1962 ();
 sg13g2_decap_8 FILLER_11_1966 ();
 sg13g2_decap_4 FILLER_11_1973 ();
 sg13g2_fill_2 FILLER_11_1977 ();
 sg13g2_fill_2 FILLER_11_1983 ();
 sg13g2_fill_2 FILLER_11_1989 ();
 sg13g2_fill_1 FILLER_11_1991 ();
 sg13g2_decap_4 FILLER_11_1997 ();
 sg13g2_fill_1 FILLER_11_2001 ();
 sg13g2_decap_4 FILLER_11_2013 ();
 sg13g2_decap_8 FILLER_11_2021 ();
 sg13g2_decap_8 FILLER_11_2028 ();
 sg13g2_decap_8 FILLER_11_2035 ();
 sg13g2_decap_8 FILLER_11_2042 ();
 sg13g2_decap_4 FILLER_11_2049 ();
 sg13g2_decap_8 FILLER_11_2069 ();
 sg13g2_decap_8 FILLER_11_2076 ();
 sg13g2_decap_8 FILLER_11_2112 ();
 sg13g2_decap_4 FILLER_11_2119 ();
 sg13g2_fill_1 FILLER_11_2123 ();
 sg13g2_decap_4 FILLER_11_2127 ();
 sg13g2_fill_1 FILLER_11_2140 ();
 sg13g2_fill_2 FILLER_11_2147 ();
 sg13g2_fill_1 FILLER_11_2175 ();
 sg13g2_fill_2 FILLER_11_2185 ();
 sg13g2_decap_4 FILLER_11_2193 ();
 sg13g2_decap_8 FILLER_11_2202 ();
 sg13g2_decap_8 FILLER_11_2209 ();
 sg13g2_decap_8 FILLER_11_2216 ();
 sg13g2_fill_2 FILLER_11_2223 ();
 sg13g2_fill_1 FILLER_11_2225 ();
 sg13g2_decap_8 FILLER_11_2230 ();
 sg13g2_decap_4 FILLER_11_2237 ();
 sg13g2_fill_2 FILLER_11_2241 ();
 sg13g2_decap_8 FILLER_11_2247 ();
 sg13g2_fill_1 FILLER_11_2254 ();
 sg13g2_decap_8 FILLER_11_2258 ();
 sg13g2_decap_8 FILLER_11_2265 ();
 sg13g2_decap_4 FILLER_11_2272 ();
 sg13g2_fill_2 FILLER_11_2276 ();
 sg13g2_fill_1 FILLER_11_2282 ();
 sg13g2_fill_2 FILLER_11_2286 ();
 sg13g2_fill_1 FILLER_11_2297 ();
 sg13g2_fill_1 FILLER_11_2305 ();
 sg13g2_decap_4 FILLER_11_2311 ();
 sg13g2_fill_2 FILLER_11_2331 ();
 sg13g2_fill_1 FILLER_11_2339 ();
 sg13g2_fill_1 FILLER_11_2384 ();
 sg13g2_fill_2 FILLER_11_2412 ();
 sg13g2_fill_2 FILLER_11_2462 ();
 sg13g2_fill_2 FILLER_11_2482 ();
 sg13g2_fill_1 FILLER_11_2484 ();
 sg13g2_decap_8 FILLER_11_2489 ();
 sg13g2_decap_8 FILLER_11_2496 ();
 sg13g2_decap_8 FILLER_11_2503 ();
 sg13g2_decap_8 FILLER_11_2510 ();
 sg13g2_decap_8 FILLER_11_2517 ();
 sg13g2_decap_8 FILLER_11_2524 ();
 sg13g2_decap_8 FILLER_11_2531 ();
 sg13g2_decap_8 FILLER_11_2538 ();
 sg13g2_decap_8 FILLER_11_2545 ();
 sg13g2_decap_8 FILLER_11_2552 ();
 sg13g2_decap_8 FILLER_11_2559 ();
 sg13g2_decap_8 FILLER_11_2566 ();
 sg13g2_decap_8 FILLER_11_2573 ();
 sg13g2_decap_8 FILLER_11_2580 ();
 sg13g2_decap_8 FILLER_11_2587 ();
 sg13g2_decap_8 FILLER_11_2594 ();
 sg13g2_decap_8 FILLER_11_2601 ();
 sg13g2_decap_8 FILLER_11_2608 ();
 sg13g2_decap_8 FILLER_11_2615 ();
 sg13g2_decap_8 FILLER_11_2622 ();
 sg13g2_decap_8 FILLER_11_2629 ();
 sg13g2_decap_8 FILLER_11_2636 ();
 sg13g2_decap_8 FILLER_11_2643 ();
 sg13g2_decap_8 FILLER_11_2650 ();
 sg13g2_decap_8 FILLER_11_2657 ();
 sg13g2_decap_4 FILLER_11_2664 ();
 sg13g2_fill_2 FILLER_11_2668 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_50 ();
 sg13g2_decap_8 FILLER_12_57 ();
 sg13g2_decap_8 FILLER_12_64 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_1 FILLER_12_76 ();
 sg13g2_decap_4 FILLER_12_89 ();
 sg13g2_fill_2 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_decap_4 FILLER_12_139 ();
 sg13g2_decap_8 FILLER_12_173 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_fill_2 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_194 ();
 sg13g2_fill_2 FILLER_12_206 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_297 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_decap_4 FILLER_12_316 ();
 sg13g2_decap_4 FILLER_12_325 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_4 FILLER_12_363 ();
 sg13g2_fill_2 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_433 ();
 sg13g2_decap_8 FILLER_12_470 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_fill_2 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_510 ();
 sg13g2_fill_1 FILLER_12_538 ();
 sg13g2_fill_1 FILLER_12_545 ();
 sg13g2_fill_1 FILLER_12_619 ();
 sg13g2_decap_8 FILLER_12_626 ();
 sg13g2_decap_4 FILLER_12_633 ();
 sg13g2_fill_2 FILLER_12_652 ();
 sg13g2_fill_2 FILLER_12_727 ();
 sg13g2_fill_1 FILLER_12_764 ();
 sg13g2_decap_8 FILLER_12_824 ();
 sg13g2_decap_8 FILLER_12_831 ();
 sg13g2_fill_2 FILLER_12_838 ();
 sg13g2_decap_4 FILLER_12_845 ();
 sg13g2_fill_1 FILLER_12_849 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_fill_1 FILLER_12_888 ();
 sg13g2_fill_2 FILLER_12_908 ();
 sg13g2_fill_2 FILLER_12_937 ();
 sg13g2_fill_1 FILLER_12_950 ();
 sg13g2_fill_2 FILLER_12_976 ();
 sg13g2_fill_1 FILLER_12_1009 ();
 sg13g2_fill_2 FILLER_12_1016 ();
 sg13g2_decap_8 FILLER_12_1023 ();
 sg13g2_fill_2 FILLER_12_1034 ();
 sg13g2_fill_1 FILLER_12_1036 ();
 sg13g2_fill_1 FILLER_12_1046 ();
 sg13g2_decap_4 FILLER_12_1052 ();
 sg13g2_fill_2 FILLER_12_1056 ();
 sg13g2_fill_2 FILLER_12_1069 ();
 sg13g2_decap_8 FILLER_12_1075 ();
 sg13g2_fill_1 FILLER_12_1082 ();
 sg13g2_fill_1 FILLER_12_1148 ();
 sg13g2_fill_2 FILLER_12_1155 ();
 sg13g2_fill_1 FILLER_12_1157 ();
 sg13g2_fill_2 FILLER_12_1195 ();
 sg13g2_fill_1 FILLER_12_1230 ();
 sg13g2_decap_8 FILLER_12_1240 ();
 sg13g2_fill_2 FILLER_12_1247 ();
 sg13g2_decap_8 FILLER_12_1259 ();
 sg13g2_decap_4 FILLER_12_1297 ();
 sg13g2_fill_2 FILLER_12_1383 ();
 sg13g2_fill_1 FILLER_12_1443 ();
 sg13g2_fill_2 FILLER_12_1491 ();
 sg13g2_fill_1 FILLER_12_1519 ();
 sg13g2_fill_2 FILLER_12_1581 ();
 sg13g2_fill_2 FILLER_12_1595 ();
 sg13g2_decap_8 FILLER_12_1623 ();
 sg13g2_fill_1 FILLER_12_1630 ();
 sg13g2_fill_1 FILLER_12_1641 ();
 sg13g2_fill_1 FILLER_12_1646 ();
 sg13g2_decap_8 FILLER_12_1651 ();
 sg13g2_fill_2 FILLER_12_1658 ();
 sg13g2_fill_2 FILLER_12_1718 ();
 sg13g2_fill_1 FILLER_12_1720 ();
 sg13g2_decap_8 FILLER_12_1747 ();
 sg13g2_decap_8 FILLER_12_1754 ();
 sg13g2_fill_2 FILLER_12_1761 ();
 sg13g2_fill_1 FILLER_12_1763 ();
 sg13g2_decap_8 FILLER_12_1769 ();
 sg13g2_fill_2 FILLER_12_1776 ();
 sg13g2_decap_8 FILLER_12_1782 ();
 sg13g2_decap_8 FILLER_12_1789 ();
 sg13g2_decap_8 FILLER_12_1796 ();
 sg13g2_decap_8 FILLER_12_1803 ();
 sg13g2_fill_2 FILLER_12_1810 ();
 sg13g2_fill_1 FILLER_12_1817 ();
 sg13g2_fill_2 FILLER_12_1826 ();
 sg13g2_decap_8 FILLER_12_1842 ();
 sg13g2_fill_2 FILLER_12_1861 ();
 sg13g2_fill_1 FILLER_12_1863 ();
 sg13g2_decap_8 FILLER_12_1868 ();
 sg13g2_decap_8 FILLER_12_1875 ();
 sg13g2_fill_2 FILLER_12_1882 ();
 sg13g2_fill_2 FILLER_12_1887 ();
 sg13g2_decap_4 FILLER_12_1894 ();
 sg13g2_fill_2 FILLER_12_1898 ();
 sg13g2_decap_4 FILLER_12_1918 ();
 sg13g2_fill_2 FILLER_12_1922 ();
 sg13g2_decap_4 FILLER_12_1934 ();
 sg13g2_fill_1 FILLER_12_1938 ();
 sg13g2_decap_4 FILLER_12_1956 ();
 sg13g2_fill_2 FILLER_12_1972 ();
 sg13g2_fill_2 FILLER_12_2000 ();
 sg13g2_decap_8 FILLER_12_2028 ();
 sg13g2_decap_8 FILLER_12_2035 ();
 sg13g2_decap_4 FILLER_12_2042 ();
 sg13g2_fill_2 FILLER_12_2081 ();
 sg13g2_decap_8 FILLER_12_2099 ();
 sg13g2_fill_2 FILLER_12_2106 ();
 sg13g2_decap_8 FILLER_12_2113 ();
 sg13g2_decap_8 FILLER_12_2120 ();
 sg13g2_decap_8 FILLER_12_2153 ();
 sg13g2_decap_8 FILLER_12_2164 ();
 sg13g2_decap_8 FILLER_12_2175 ();
 sg13g2_decap_8 FILLER_12_2182 ();
 sg13g2_decap_8 FILLER_12_2189 ();
 sg13g2_decap_4 FILLER_12_2196 ();
 sg13g2_fill_1 FILLER_12_2204 ();
 sg13g2_fill_1 FILLER_12_2231 ();
 sg13g2_fill_1 FILLER_12_2242 ();
 sg13g2_decap_4 FILLER_12_2274 ();
 sg13g2_fill_2 FILLER_12_2278 ();
 sg13g2_fill_2 FILLER_12_2331 ();
 sg13g2_fill_1 FILLER_12_2341 ();
 sg13g2_fill_1 FILLER_12_2455 ();
 sg13g2_decap_8 FILLER_12_2462 ();
 sg13g2_decap_4 FILLER_12_2469 ();
 sg13g2_fill_1 FILLER_12_2473 ();
 sg13g2_fill_2 FILLER_12_2504 ();
 sg13g2_decap_8 FILLER_12_2510 ();
 sg13g2_decap_4 FILLER_12_2517 ();
 sg13g2_fill_2 FILLER_12_2521 ();
 sg13g2_decap_8 FILLER_12_2553 ();
 sg13g2_decap_8 FILLER_12_2560 ();
 sg13g2_decap_8 FILLER_12_2567 ();
 sg13g2_decap_8 FILLER_12_2574 ();
 sg13g2_decap_8 FILLER_12_2581 ();
 sg13g2_decap_8 FILLER_12_2588 ();
 sg13g2_decap_8 FILLER_12_2595 ();
 sg13g2_decap_8 FILLER_12_2602 ();
 sg13g2_decap_8 FILLER_12_2609 ();
 sg13g2_decap_8 FILLER_12_2616 ();
 sg13g2_decap_8 FILLER_12_2623 ();
 sg13g2_decap_8 FILLER_12_2630 ();
 sg13g2_decap_8 FILLER_12_2637 ();
 sg13g2_decap_8 FILLER_12_2644 ();
 sg13g2_decap_8 FILLER_12_2651 ();
 sg13g2_decap_8 FILLER_12_2658 ();
 sg13g2_decap_4 FILLER_12_2665 ();
 sg13g2_fill_1 FILLER_12_2669 ();
 sg13g2_fill_2 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_143 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_2 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_220 ();
 sg13g2_fill_1 FILLER_13_222 ();
 sg13g2_decap_8 FILLER_13_227 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_decap_4 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_decap_4 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_4 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_fill_2 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_13_418 ();
 sg13g2_fill_2 FILLER_13_452 ();
 sg13g2_fill_1 FILLER_13_459 ();
 sg13g2_fill_2 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_492 ();
 sg13g2_decap_8 FILLER_13_499 ();
 sg13g2_fill_2 FILLER_13_519 ();
 sg13g2_fill_1 FILLER_13_529 ();
 sg13g2_fill_2 FILLER_13_535 ();
 sg13g2_fill_1 FILLER_13_537 ();
 sg13g2_fill_2 FILLER_13_573 ();
 sg13g2_fill_2 FILLER_13_606 ();
 sg13g2_fill_1 FILLER_13_693 ();
 sg13g2_fill_2 FILLER_13_701 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_fill_2 FILLER_13_721 ();
 sg13g2_fill_1 FILLER_13_723 ();
 sg13g2_fill_1 FILLER_13_754 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_decap_8 FILLER_13_797 ();
 sg13g2_decap_8 FILLER_13_804 ();
 sg13g2_decap_8 FILLER_13_811 ();
 sg13g2_decap_8 FILLER_13_818 ();
 sg13g2_decap_8 FILLER_13_825 ();
 sg13g2_decap_4 FILLER_13_832 ();
 sg13g2_fill_2 FILLER_13_836 ();
 sg13g2_decap_8 FILLER_13_864 ();
 sg13g2_fill_2 FILLER_13_871 ();
 sg13g2_fill_1 FILLER_13_873 ();
 sg13g2_decap_8 FILLER_13_878 ();
 sg13g2_fill_2 FILLER_13_893 ();
 sg13g2_fill_1 FILLER_13_942 ();
 sg13g2_fill_1 FILLER_13_985 ();
 sg13g2_fill_1 FILLER_13_992 ();
 sg13g2_fill_1 FILLER_13_999 ();
 sg13g2_fill_1 FILLER_13_1010 ();
 sg13g2_decap_8 FILLER_13_1018 ();
 sg13g2_fill_1 FILLER_13_1025 ();
 sg13g2_decap_8 FILLER_13_1031 ();
 sg13g2_fill_2 FILLER_13_1038 ();
 sg13g2_fill_1 FILLER_13_1040 ();
 sg13g2_decap_8 FILLER_13_1057 ();
 sg13g2_decap_4 FILLER_13_1064 ();
 sg13g2_fill_2 FILLER_13_1068 ();
 sg13g2_decap_8 FILLER_13_1073 ();
 sg13g2_fill_2 FILLER_13_1080 ();
 sg13g2_fill_1 FILLER_13_1082 ();
 sg13g2_decap_8 FILLER_13_1091 ();
 sg13g2_decap_8 FILLER_13_1098 ();
 sg13g2_fill_2 FILLER_13_1111 ();
 sg13g2_fill_2 FILLER_13_1121 ();
 sg13g2_fill_1 FILLER_13_1129 ();
 sg13g2_fill_2 FILLER_13_1136 ();
 sg13g2_fill_1 FILLER_13_1138 ();
 sg13g2_decap_4 FILLER_13_1145 ();
 sg13g2_fill_1 FILLER_13_1149 ();
 sg13g2_fill_2 FILLER_13_1156 ();
 sg13g2_decap_8 FILLER_13_1208 ();
 sg13g2_decap_4 FILLER_13_1215 ();
 sg13g2_fill_1 FILLER_13_1219 ();
 sg13g2_decap_8 FILLER_13_1232 ();
 sg13g2_decap_8 FILLER_13_1239 ();
 sg13g2_decap_8 FILLER_13_1246 ();
 sg13g2_decap_8 FILLER_13_1253 ();
 sg13g2_decap_8 FILLER_13_1260 ();
 sg13g2_decap_8 FILLER_13_1267 ();
 sg13g2_decap_8 FILLER_13_1274 ();
 sg13g2_decap_4 FILLER_13_1281 ();
 sg13g2_fill_1 FILLER_13_1296 ();
 sg13g2_fill_2 FILLER_13_1325 ();
 sg13g2_fill_1 FILLER_13_1347 ();
 sg13g2_fill_2 FILLER_13_1360 ();
 sg13g2_fill_2 FILLER_13_1373 ();
 sg13g2_fill_2 FILLER_13_1422 ();
 sg13g2_fill_2 FILLER_13_1431 ();
 sg13g2_decap_8 FILLER_13_1505 ();
 sg13g2_decap_8 FILLER_13_1512 ();
 sg13g2_fill_2 FILLER_13_1519 ();
 sg13g2_fill_1 FILLER_13_1521 ();
 sg13g2_decap_8 FILLER_13_1543 ();
 sg13g2_fill_1 FILLER_13_1550 ();
 sg13g2_fill_2 FILLER_13_1565 ();
 sg13g2_decap_8 FILLER_13_1593 ();
 sg13g2_decap_4 FILLER_13_1600 ();
 sg13g2_fill_2 FILLER_13_1604 ();
 sg13g2_decap_8 FILLER_13_1615 ();
 sg13g2_decap_4 FILLER_13_1622 ();
 sg13g2_fill_2 FILLER_13_1631 ();
 sg13g2_fill_2 FILLER_13_1651 ();
 sg13g2_fill_1 FILLER_13_1653 ();
 sg13g2_decap_8 FILLER_13_1685 ();
 sg13g2_decap_8 FILLER_13_1692 ();
 sg13g2_fill_2 FILLER_13_1699 ();
 sg13g2_fill_1 FILLER_13_1701 ();
 sg13g2_decap_8 FILLER_13_1711 ();
 sg13g2_fill_2 FILLER_13_1718 ();
 sg13g2_fill_1 FILLER_13_1720 ();
 sg13g2_fill_1 FILLER_13_1727 ();
 sg13g2_decap_8 FILLER_13_1732 ();
 sg13g2_fill_2 FILLER_13_1747 ();
 sg13g2_fill_1 FILLER_13_1749 ();
 sg13g2_fill_1 FILLER_13_1784 ();
 sg13g2_decap_8 FILLER_13_1790 ();
 sg13g2_decap_8 FILLER_13_1797 ();
 sg13g2_fill_1 FILLER_13_1804 ();
 sg13g2_fill_2 FILLER_13_1834 ();
 sg13g2_fill_2 FILLER_13_1854 ();
 sg13g2_fill_1 FILLER_13_1856 ();
 sg13g2_decap_4 FILLER_13_1894 ();
 sg13g2_fill_1 FILLER_13_1898 ();
 sg13g2_decap_4 FILLER_13_1904 ();
 sg13g2_decap_8 FILLER_13_1913 ();
 sg13g2_fill_2 FILLER_13_1920 ();
 sg13g2_fill_1 FILLER_13_1958 ();
 sg13g2_fill_2 FILLER_13_2021 ();
 sg13g2_fill_1 FILLER_13_2023 ();
 sg13g2_fill_2 FILLER_13_2028 ();
 sg13g2_fill_1 FILLER_13_2030 ();
 sg13g2_decap_8 FILLER_13_2070 ();
 sg13g2_decap_8 FILLER_13_2077 ();
 sg13g2_fill_2 FILLER_13_2084 ();
 sg13g2_fill_1 FILLER_13_2086 ();
 sg13g2_decap_8 FILLER_13_2122 ();
 sg13g2_decap_8 FILLER_13_2129 ();
 sg13g2_decap_8 FILLER_13_2136 ();
 sg13g2_fill_1 FILLER_13_2143 ();
 sg13g2_fill_1 FILLER_13_2170 ();
 sg13g2_decap_8 FILLER_13_2177 ();
 sg13g2_decap_4 FILLER_13_2184 ();
 sg13g2_decap_4 FILLER_13_2193 ();
 sg13g2_fill_1 FILLER_13_2197 ();
 sg13g2_fill_2 FILLER_13_2203 ();
 sg13g2_fill_1 FILLER_13_2205 ();
 sg13g2_fill_2 FILLER_13_2212 ();
 sg13g2_fill_2 FILLER_13_2217 ();
 sg13g2_decap_4 FILLER_13_2228 ();
 sg13g2_fill_1 FILLER_13_2232 ();
 sg13g2_fill_1 FILLER_13_2239 ();
 sg13g2_fill_1 FILLER_13_2299 ();
 sg13g2_fill_1 FILLER_13_2305 ();
 sg13g2_fill_2 FILLER_13_2323 ();
 sg13g2_fill_1 FILLER_13_2331 ();
 sg13g2_fill_1 FILLER_13_2352 ();
 sg13g2_fill_1 FILLER_13_2387 ();
 sg13g2_decap_4 FILLER_13_2398 ();
 sg13g2_fill_1 FILLER_13_2402 ();
 sg13g2_fill_2 FILLER_13_2422 ();
 sg13g2_fill_1 FILLER_13_2430 ();
 sg13g2_fill_1 FILLER_13_2439 ();
 sg13g2_decap_8 FILLER_13_2448 ();
 sg13g2_decap_8 FILLER_13_2455 ();
 sg13g2_decap_4 FILLER_13_2462 ();
 sg13g2_decap_8 FILLER_13_2470 ();
 sg13g2_fill_1 FILLER_13_2477 ();
 sg13g2_fill_2 FILLER_13_2484 ();
 sg13g2_fill_2 FILLER_13_2496 ();
 sg13g2_fill_1 FILLER_13_2498 ();
 sg13g2_fill_2 FILLER_13_2525 ();
 sg13g2_decap_8 FILLER_13_2553 ();
 sg13g2_decap_8 FILLER_13_2560 ();
 sg13g2_decap_8 FILLER_13_2567 ();
 sg13g2_decap_8 FILLER_13_2574 ();
 sg13g2_decap_8 FILLER_13_2581 ();
 sg13g2_decap_8 FILLER_13_2588 ();
 sg13g2_decap_8 FILLER_13_2595 ();
 sg13g2_decap_8 FILLER_13_2602 ();
 sg13g2_decap_8 FILLER_13_2609 ();
 sg13g2_decap_8 FILLER_13_2616 ();
 sg13g2_decap_8 FILLER_13_2623 ();
 sg13g2_decap_8 FILLER_13_2630 ();
 sg13g2_decap_8 FILLER_13_2637 ();
 sg13g2_decap_8 FILLER_13_2644 ();
 sg13g2_decap_8 FILLER_13_2651 ();
 sg13g2_decap_8 FILLER_13_2658 ();
 sg13g2_decap_4 FILLER_13_2665 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_9 ();
 sg13g2_decap_8 FILLER_14_22 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_4 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_106 ();
 sg13g2_decap_8 FILLER_14_113 ();
 sg13g2_decap_4 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_124 ();
 sg13g2_fill_1 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_14_204 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_2 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_decap_4 FILLER_14_397 ();
 sg13g2_fill_2 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_4 FILLER_14_454 ();
 sg13g2_decap_8 FILLER_14_471 ();
 sg13g2_decap_8 FILLER_14_478 ();
 sg13g2_fill_2 FILLER_14_485 ();
 sg13g2_decap_4 FILLER_14_490 ();
 sg13g2_fill_2 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_527 ();
 sg13g2_decap_4 FILLER_14_570 ();
 sg13g2_decap_4 FILLER_14_587 ();
 sg13g2_fill_1 FILLER_14_591 ();
 sg13g2_fill_2 FILLER_14_651 ();
 sg13g2_fill_1 FILLER_14_697 ();
 sg13g2_fill_1 FILLER_14_708 ();
 sg13g2_decap_4 FILLER_14_713 ();
 sg13g2_fill_2 FILLER_14_717 ();
 sg13g2_decap_8 FILLER_14_723 ();
 sg13g2_decap_4 FILLER_14_730 ();
 sg13g2_fill_1 FILLER_14_734 ();
 sg13g2_fill_2 FILLER_14_743 ();
 sg13g2_fill_1 FILLER_14_745 ();
 sg13g2_fill_1 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_fill_2 FILLER_14_800 ();
 sg13g2_fill_1 FILLER_14_802 ();
 sg13g2_fill_2 FILLER_14_843 ();
 sg13g2_fill_1 FILLER_14_845 ();
 sg13g2_fill_1 FILLER_14_876 ();
 sg13g2_decap_8 FILLER_14_882 ();
 sg13g2_decap_4 FILLER_14_889 ();
 sg13g2_fill_2 FILLER_14_893 ();
 sg13g2_fill_1 FILLER_14_901 ();
 sg13g2_fill_1 FILLER_14_968 ();
 sg13g2_decap_8 FILLER_14_1021 ();
 sg13g2_decap_4 FILLER_14_1028 ();
 sg13g2_fill_1 FILLER_14_1063 ();
 sg13g2_fill_1 FILLER_14_1073 ();
 sg13g2_decap_8 FILLER_14_1081 ();
 sg13g2_decap_4 FILLER_14_1097 ();
 sg13g2_fill_2 FILLER_14_1101 ();
 sg13g2_decap_8 FILLER_14_1123 ();
 sg13g2_fill_2 FILLER_14_1130 ();
 sg13g2_fill_2 FILLER_14_1143 ();
 sg13g2_decap_4 FILLER_14_1159 ();
 sg13g2_fill_2 FILLER_14_1163 ();
 sg13g2_fill_2 FILLER_14_1169 ();
 sg13g2_fill_2 FILLER_14_1182 ();
 sg13g2_fill_2 FILLER_14_1205 ();
 sg13g2_decap_4 FILLER_14_1213 ();
 sg13g2_fill_2 FILLER_14_1217 ();
 sg13g2_fill_1 FILLER_14_1227 ();
 sg13g2_fill_2 FILLER_14_1254 ();
 sg13g2_fill_1 FILLER_14_1256 ();
 sg13g2_decap_4 FILLER_14_1292 ();
 sg13g2_fill_1 FILLER_14_1296 ();
 sg13g2_fill_2 FILLER_14_1362 ();
 sg13g2_fill_1 FILLER_14_1370 ();
 sg13g2_fill_2 FILLER_14_1409 ();
 sg13g2_fill_2 FILLER_14_1416 ();
 sg13g2_fill_1 FILLER_14_1428 ();
 sg13g2_fill_1 FILLER_14_1460 ();
 sg13g2_fill_1 FILLER_14_1488 ();
 sg13g2_fill_2 FILLER_14_1515 ();
 sg13g2_fill_1 FILLER_14_1517 ();
 sg13g2_fill_1 FILLER_14_1544 ();
 sg13g2_fill_1 FILLER_14_1550 ();
 sg13g2_fill_1 FILLER_14_1555 ();
 sg13g2_fill_2 FILLER_14_1560 ();
 sg13g2_decap_8 FILLER_14_1571 ();
 sg13g2_decap_8 FILLER_14_1578 ();
 sg13g2_fill_1 FILLER_14_1585 ();
 sg13g2_fill_1 FILLER_14_1590 ();
 sg13g2_fill_1 FILLER_14_1645 ();
 sg13g2_fill_2 FILLER_14_1677 ();
 sg13g2_fill_2 FILLER_14_1705 ();
 sg13g2_fill_1 FILLER_14_1707 ();
 sg13g2_fill_1 FILLER_14_1714 ();
 sg13g2_fill_1 FILLER_14_1721 ();
 sg13g2_fill_1 FILLER_14_1748 ();
 sg13g2_fill_2 FILLER_14_1753 ();
 sg13g2_fill_1 FILLER_14_1760 ();
 sg13g2_fill_1 FILLER_14_1787 ();
 sg13g2_fill_2 FILLER_14_1829 ();
 sg13g2_decap_4 FILLER_14_1857 ();
 sg13g2_decap_4 FILLER_14_1869 ();
 sg13g2_decap_4 FILLER_14_1879 ();
 sg13g2_fill_2 FILLER_14_2006 ();
 sg13g2_decap_4 FILLER_14_2048 ();
 sg13g2_decap_4 FILLER_14_2056 ();
 sg13g2_decap_8 FILLER_14_2066 ();
 sg13g2_decap_8 FILLER_14_2073 ();
 sg13g2_fill_2 FILLER_14_2080 ();
 sg13g2_fill_1 FILLER_14_2082 ();
 sg13g2_decap_8 FILLER_14_2093 ();
 sg13g2_decap_8 FILLER_14_2130 ();
 sg13g2_decap_4 FILLER_14_2137 ();
 sg13g2_decap_4 FILLER_14_2150 ();
 sg13g2_fill_2 FILLER_14_2154 ();
 sg13g2_decap_4 FILLER_14_2178 ();
 sg13g2_fill_1 FILLER_14_2182 ();
 sg13g2_fill_2 FILLER_14_2267 ();
 sg13g2_fill_2 FILLER_14_2300 ();
 sg13g2_fill_1 FILLER_14_2352 ();
 sg13g2_fill_1 FILLER_14_2385 ();
 sg13g2_fill_2 FILLER_14_2394 ();
 sg13g2_decap_8 FILLER_14_2404 ();
 sg13g2_decap_8 FILLER_14_2411 ();
 sg13g2_decap_8 FILLER_14_2418 ();
 sg13g2_fill_1 FILLER_14_2455 ();
 sg13g2_fill_2 FILLER_14_2486 ();
 sg13g2_fill_1 FILLER_14_2488 ();
 sg13g2_decap_4 FILLER_14_2506 ();
 sg13g2_fill_1 FILLER_14_2510 ();
 sg13g2_decap_8 FILLER_14_2517 ();
 sg13g2_fill_1 FILLER_14_2524 ();
 sg13g2_decap_8 FILLER_14_2547 ();
 sg13g2_decap_8 FILLER_14_2554 ();
 sg13g2_decap_8 FILLER_14_2561 ();
 sg13g2_decap_8 FILLER_14_2568 ();
 sg13g2_decap_8 FILLER_14_2575 ();
 sg13g2_decap_8 FILLER_14_2582 ();
 sg13g2_decap_8 FILLER_14_2589 ();
 sg13g2_decap_8 FILLER_14_2596 ();
 sg13g2_decap_8 FILLER_14_2603 ();
 sg13g2_decap_8 FILLER_14_2610 ();
 sg13g2_decap_8 FILLER_14_2617 ();
 sg13g2_decap_8 FILLER_14_2624 ();
 sg13g2_decap_8 FILLER_14_2631 ();
 sg13g2_decap_8 FILLER_14_2638 ();
 sg13g2_decap_8 FILLER_14_2645 ();
 sg13g2_decap_8 FILLER_14_2652 ();
 sg13g2_decap_8 FILLER_14_2659 ();
 sg13g2_decap_4 FILLER_14_2666 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_33 ();
 sg13g2_decap_4 FILLER_15_40 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_decap_8 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_76 ();
 sg13g2_fill_2 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_4 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_246 ();
 sg13g2_decap_4 FILLER_15_261 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_1 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_433 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_fill_2 FILLER_15_459 ();
 sg13g2_fill_1 FILLER_15_461 ();
 sg13g2_decap_8 FILLER_15_499 ();
 sg13g2_fill_1 FILLER_15_510 ();
 sg13g2_fill_2 FILLER_15_515 ();
 sg13g2_fill_1 FILLER_15_517 ();
 sg13g2_decap_4 FILLER_15_571 ();
 sg13g2_fill_2 FILLER_15_575 ();
 sg13g2_fill_2 FILLER_15_616 ();
 sg13g2_fill_1 FILLER_15_618 ();
 sg13g2_fill_1 FILLER_15_658 ();
 sg13g2_fill_2 FILLER_15_668 ();
 sg13g2_fill_1 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_684 ();
 sg13g2_decap_8 FILLER_15_691 ();
 sg13g2_decap_8 FILLER_15_698 ();
 sg13g2_decap_4 FILLER_15_705 ();
 sg13g2_fill_2 FILLER_15_709 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_decap_8 FILLER_15_731 ();
 sg13g2_fill_1 FILLER_15_738 ();
 sg13g2_fill_2 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_fill_2 FILLER_15_798 ();
 sg13g2_fill_1 FILLER_15_830 ();
 sg13g2_fill_2 FILLER_15_839 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_decap_4 FILLER_15_879 ();
 sg13g2_decap_4 FILLER_15_887 ();
 sg13g2_fill_1 FILLER_15_917 ();
 sg13g2_fill_2 FILLER_15_926 ();
 sg13g2_fill_2 FILLER_15_934 ();
 sg13g2_fill_1 FILLER_15_976 ();
 sg13g2_fill_1 FILLER_15_1010 ();
 sg13g2_decap_8 FILLER_15_1016 ();
 sg13g2_decap_8 FILLER_15_1023 ();
 sg13g2_fill_2 FILLER_15_1030 ();
 sg13g2_fill_1 FILLER_15_1032 ();
 sg13g2_decap_4 FILLER_15_1038 ();
 sg13g2_fill_2 FILLER_15_1042 ();
 sg13g2_fill_1 FILLER_15_1052 ();
 sg13g2_fill_1 FILLER_15_1059 ();
 sg13g2_fill_1 FILLER_15_1095 ();
 sg13g2_fill_1 FILLER_15_1102 ();
 sg13g2_decap_4 FILLER_15_1108 ();
 sg13g2_fill_1 FILLER_15_1118 ();
 sg13g2_decap_4 FILLER_15_1124 ();
 sg13g2_fill_2 FILLER_15_1128 ();
 sg13g2_decap_8 FILLER_15_1150 ();
 sg13g2_fill_2 FILLER_15_1157 ();
 sg13g2_fill_1 FILLER_15_1159 ();
 sg13g2_fill_1 FILLER_15_1186 ();
 sg13g2_fill_2 FILLER_15_1195 ();
 sg13g2_decap_4 FILLER_15_1206 ();
 sg13g2_fill_2 FILLER_15_1210 ();
 sg13g2_decap_8 FILLER_15_1218 ();
 sg13g2_fill_1 FILLER_15_1225 ();
 sg13g2_decap_8 FILLER_15_1241 ();
 sg13g2_decap_4 FILLER_15_1258 ();
 sg13g2_decap_8 FILLER_15_1271 ();
 sg13g2_fill_2 FILLER_15_1278 ();
 sg13g2_fill_1 FILLER_15_1280 ();
 sg13g2_fill_1 FILLER_15_1292 ();
 sg13g2_fill_1 FILLER_15_1299 ();
 sg13g2_fill_1 FILLER_15_1305 ();
 sg13g2_fill_1 FILLER_15_1310 ();
 sg13g2_fill_2 FILLER_15_1336 ();
 sg13g2_decap_8 FILLER_15_1347 ();
 sg13g2_decap_4 FILLER_15_1354 ();
 sg13g2_fill_1 FILLER_15_1369 ();
 sg13g2_fill_2 FILLER_15_1448 ();
 sg13g2_fill_1 FILLER_15_1481 ();
 sg13g2_decap_8 FILLER_15_1495 ();
 sg13g2_fill_2 FILLER_15_1502 ();
 sg13g2_fill_2 FILLER_15_1539 ();
 sg13g2_fill_1 FILLER_15_1541 ();
 sg13g2_fill_1 FILLER_15_1578 ();
 sg13g2_decap_8 FILLER_15_1585 ();
 sg13g2_decap_8 FILLER_15_1592 ();
 sg13g2_decap_8 FILLER_15_1599 ();
 sg13g2_fill_1 FILLER_15_1606 ();
 sg13g2_fill_2 FILLER_15_1633 ();
 sg13g2_fill_1 FILLER_15_1635 ();
 sg13g2_decap_8 FILLER_15_1645 ();
 sg13g2_decap_8 FILLER_15_1652 ();
 sg13g2_decap_4 FILLER_15_1659 ();
 sg13g2_decap_8 FILLER_15_1666 ();
 sg13g2_decap_8 FILLER_15_1673 ();
 sg13g2_fill_2 FILLER_15_1680 ();
 sg13g2_fill_1 FILLER_15_1682 ();
 sg13g2_fill_2 FILLER_15_1688 ();
 sg13g2_fill_2 FILLER_15_1712 ();
 sg13g2_decap_8 FILLER_15_1720 ();
 sg13g2_fill_2 FILLER_15_1727 ();
 sg13g2_fill_1 FILLER_15_1735 ();
 sg13g2_fill_1 FILLER_15_1741 ();
 sg13g2_fill_2 FILLER_15_1817 ();
 sg13g2_fill_2 FILLER_15_1825 ();
 sg13g2_fill_2 FILLER_15_1831 ();
 sg13g2_decap_4 FILLER_15_1855 ();
 sg13g2_fill_1 FILLER_15_1859 ();
 sg13g2_decap_8 FILLER_15_1886 ();
 sg13g2_decap_8 FILLER_15_1893 ();
 sg13g2_decap_8 FILLER_15_1900 ();
 sg13g2_decap_8 FILLER_15_1907 ();
 sg13g2_decap_8 FILLER_15_1914 ();
 sg13g2_fill_1 FILLER_15_1929 ();
 sg13g2_fill_2 FILLER_15_1963 ();
 sg13g2_fill_1 FILLER_15_1970 ();
 sg13g2_fill_2 FILLER_15_1977 ();
 sg13g2_fill_1 FILLER_15_1984 ();
 sg13g2_fill_2 FILLER_15_2034 ();
 sg13g2_fill_1 FILLER_15_2036 ();
 sg13g2_decap_8 FILLER_15_2049 ();
 sg13g2_fill_2 FILLER_15_2092 ();
 sg13g2_decap_4 FILLER_15_2140 ();
 sg13g2_fill_2 FILLER_15_2151 ();
 sg13g2_fill_1 FILLER_15_2163 ();
 sg13g2_fill_2 FILLER_15_2167 ();
 sg13g2_fill_2 FILLER_15_2199 ();
 sg13g2_fill_2 FILLER_15_2232 ();
 sg13g2_fill_2 FILLER_15_2260 ();
 sg13g2_fill_2 FILLER_15_2278 ();
 sg13g2_decap_4 FILLER_15_2290 ();
 sg13g2_fill_1 FILLER_15_2294 ();
 sg13g2_fill_2 FILLER_15_2311 ();
 sg13g2_fill_2 FILLER_15_2375 ();
 sg13g2_decap_8 FILLER_15_2408 ();
 sg13g2_decap_8 FILLER_15_2415 ();
 sg13g2_fill_2 FILLER_15_2422 ();
 sg13g2_decap_8 FILLER_15_2428 ();
 sg13g2_decap_8 FILLER_15_2435 ();
 sg13g2_decap_8 FILLER_15_2448 ();
 sg13g2_fill_1 FILLER_15_2455 ();
 sg13g2_fill_2 FILLER_15_2486 ();
 sg13g2_fill_1 FILLER_15_2488 ();
 sg13g2_fill_1 FILLER_15_2519 ();
 sg13g2_decap_8 FILLER_15_2524 ();
 sg13g2_decap_8 FILLER_15_2531 ();
 sg13g2_decap_8 FILLER_15_2538 ();
 sg13g2_decap_8 FILLER_15_2545 ();
 sg13g2_decap_8 FILLER_15_2552 ();
 sg13g2_decap_8 FILLER_15_2559 ();
 sg13g2_decap_8 FILLER_15_2566 ();
 sg13g2_decap_8 FILLER_15_2573 ();
 sg13g2_decap_8 FILLER_15_2580 ();
 sg13g2_decap_8 FILLER_15_2587 ();
 sg13g2_decap_8 FILLER_15_2594 ();
 sg13g2_decap_8 FILLER_15_2601 ();
 sg13g2_decap_8 FILLER_15_2608 ();
 sg13g2_decap_8 FILLER_15_2615 ();
 sg13g2_decap_8 FILLER_15_2622 ();
 sg13g2_decap_8 FILLER_15_2629 ();
 sg13g2_decap_8 FILLER_15_2636 ();
 sg13g2_decap_8 FILLER_15_2643 ();
 sg13g2_decap_8 FILLER_15_2650 ();
 sg13g2_decap_8 FILLER_15_2657 ();
 sg13g2_decap_4 FILLER_15_2664 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_17 ();
 sg13g2_fill_1 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_2 FILLER_16_46 ();
 sg13g2_fill_1 FILLER_16_78 ();
 sg13g2_decap_8 FILLER_16_83 ();
 sg13g2_decap_8 FILLER_16_90 ();
 sg13g2_decap_8 FILLER_16_97 ();
 sg13g2_decap_8 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_fill_2 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_131 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_decap_4 FILLER_16_174 ();
 sg13g2_decap_4 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_decap_4 FILLER_16_327 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_decap_4 FILLER_16_337 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_1 FILLER_16_395 ();
 sg13g2_fill_2 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_403 ();
 sg13g2_decap_4 FILLER_16_409 ();
 sg13g2_fill_2 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_fill_2 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_468 ();
 sg13g2_decap_8 FILLER_16_475 ();
 sg13g2_decap_8 FILLER_16_482 ();
 sg13g2_decap_8 FILLER_16_489 ();
 sg13g2_decap_8 FILLER_16_496 ();
 sg13g2_decap_4 FILLER_16_503 ();
 sg13g2_fill_1 FILLER_16_507 ();
 sg13g2_decap_4 FILLER_16_547 ();
 sg13g2_fill_2 FILLER_16_551 ();
 sg13g2_decap_8 FILLER_16_579 ();
 sg13g2_decap_8 FILLER_16_586 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_fill_2 FILLER_16_600 ();
 sg13g2_fill_1 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_fill_2 FILLER_16_623 ();
 sg13g2_fill_1 FILLER_16_625 ();
 sg13g2_fill_2 FILLER_16_654 ();
 sg13g2_decap_8 FILLER_16_673 ();
 sg13g2_decap_8 FILLER_16_680 ();
 sg13g2_decap_8 FILLER_16_687 ();
 sg13g2_decap_8 FILLER_16_694 ();
 sg13g2_fill_2 FILLER_16_701 ();
 sg13g2_fill_2 FILLER_16_734 ();
 sg13g2_fill_1 FILLER_16_757 ();
 sg13g2_decap_4 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_4 FILLER_16_840 ();
 sg13g2_fill_1 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_857 ();
 sg13g2_fill_2 FILLER_16_868 ();
 sg13g2_fill_1 FILLER_16_905 ();
 sg13g2_fill_2 FILLER_16_944 ();
 sg13g2_fill_2 FILLER_16_954 ();
 sg13g2_fill_2 FILLER_16_961 ();
 sg13g2_fill_1 FILLER_16_989 ();
 sg13g2_fill_1 FILLER_16_995 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_fill_1 FILLER_16_1029 ();
 sg13g2_decap_8 FILLER_16_1061 ();
 sg13g2_fill_2 FILLER_16_1068 ();
 sg13g2_decap_4 FILLER_16_1076 ();
 sg13g2_fill_1 FILLER_16_1125 ();
 sg13g2_fill_2 FILLER_16_1148 ();
 sg13g2_fill_2 FILLER_16_1154 ();
 sg13g2_fill_1 FILLER_16_1156 ();
 sg13g2_decap_8 FILLER_16_1161 ();
 sg13g2_decap_4 FILLER_16_1168 ();
 sg13g2_fill_1 FILLER_16_1172 ();
 sg13g2_fill_1 FILLER_16_1183 ();
 sg13g2_fill_2 FILLER_16_1189 ();
 sg13g2_fill_2 FILLER_16_1203 ();
 sg13g2_decap_8 FILLER_16_1210 ();
 sg13g2_fill_2 FILLER_16_1217 ();
 sg13g2_decap_4 FILLER_16_1233 ();
 sg13g2_fill_2 FILLER_16_1242 ();
 sg13g2_fill_1 FILLER_16_1257 ();
 sg13g2_decap_8 FILLER_16_1268 ();
 sg13g2_decap_4 FILLER_16_1275 ();
 sg13g2_fill_1 FILLER_16_1279 ();
 sg13g2_fill_1 FILLER_16_1285 ();
 sg13g2_fill_1 FILLER_16_1290 ();
 sg13g2_fill_1 FILLER_16_1320 ();
 sg13g2_decap_4 FILLER_16_1358 ();
 sg13g2_fill_2 FILLER_16_1362 ();
 sg13g2_fill_1 FILLER_16_1387 ();
 sg13g2_fill_1 FILLER_16_1404 ();
 sg13g2_fill_2 FILLER_16_1424 ();
 sg13g2_fill_1 FILLER_16_1460 ();
 sg13g2_decap_8 FILLER_16_1466 ();
 sg13g2_decap_4 FILLER_16_1473 ();
 sg13g2_decap_8 FILLER_16_1480 ();
 sg13g2_decap_8 FILLER_16_1487 ();
 sg13g2_decap_8 FILLER_16_1494 ();
 sg13g2_decap_8 FILLER_16_1501 ();
 sg13g2_decap_8 FILLER_16_1508 ();
 sg13g2_fill_1 FILLER_16_1515 ();
 sg13g2_fill_1 FILLER_16_1521 ();
 sg13g2_fill_2 FILLER_16_1526 ();
 sg13g2_decap_4 FILLER_16_1532 ();
 sg13g2_fill_2 FILLER_16_1536 ();
 sg13g2_fill_2 FILLER_16_1569 ();
 sg13g2_fill_1 FILLER_16_1628 ();
 sg13g2_decap_4 FILLER_16_1637 ();
 sg13g2_fill_1 FILLER_16_1641 ();
 sg13g2_decap_8 FILLER_16_1671 ();
 sg13g2_decap_8 FILLER_16_1678 ();
 sg13g2_decap_8 FILLER_16_1685 ();
 sg13g2_decap_8 FILLER_16_1692 ();
 sg13g2_decap_8 FILLER_16_1699 ();
 sg13g2_fill_1 FILLER_16_1706 ();
 sg13g2_decap_4 FILLER_16_1718 ();
 sg13g2_fill_2 FILLER_16_1722 ();
 sg13g2_decap_4 FILLER_16_1750 ();
 sg13g2_fill_1 FILLER_16_1754 ();
 sg13g2_decap_8 FILLER_16_1764 ();
 sg13g2_decap_8 FILLER_16_1771 ();
 sg13g2_fill_2 FILLER_16_1778 ();
 sg13g2_fill_2 FILLER_16_1795 ();
 sg13g2_decap_8 FILLER_16_1802 ();
 sg13g2_fill_2 FILLER_16_1809 ();
 sg13g2_decap_8 FILLER_16_1824 ();
 sg13g2_fill_1 FILLER_16_1831 ();
 sg13g2_fill_1 FILLER_16_1837 ();
 sg13g2_fill_2 FILLER_16_1869 ();
 sg13g2_decap_8 FILLER_16_1875 ();
 sg13g2_decap_8 FILLER_16_1882 ();
 sg13g2_decap_8 FILLER_16_1889 ();
 sg13g2_fill_2 FILLER_16_1950 ();
 sg13g2_fill_1 FILLER_16_1952 ();
 sg13g2_fill_2 FILLER_16_1979 ();
 sg13g2_fill_1 FILLER_16_2003 ();
 sg13g2_decap_8 FILLER_16_2007 ();
 sg13g2_decap_8 FILLER_16_2014 ();
 sg13g2_fill_1 FILLER_16_2021 ();
 sg13g2_decap_8 FILLER_16_2048 ();
 sg13g2_decap_8 FILLER_16_2055 ();
 sg13g2_fill_1 FILLER_16_2062 ();
 sg13g2_decap_4 FILLER_16_2071 ();
 sg13g2_fill_1 FILLER_16_2085 ();
 sg13g2_decap_8 FILLER_16_2106 ();
 sg13g2_fill_1 FILLER_16_2121 ();
 sg13g2_decap_4 FILLER_16_2198 ();
 sg13g2_fill_2 FILLER_16_2202 ();
 sg13g2_fill_2 FILLER_16_2212 ();
 sg13g2_decap_8 FILLER_16_2232 ();
 sg13g2_decap_4 FILLER_16_2248 ();
 sg13g2_fill_2 FILLER_16_2252 ();
 sg13g2_decap_4 FILLER_16_2260 ();
 sg13g2_fill_2 FILLER_16_2319 ();
 sg13g2_fill_1 FILLER_16_2333 ();
 sg13g2_fill_1 FILLER_16_2368 ();
 sg13g2_fill_2 FILLER_16_2385 ();
 sg13g2_fill_2 FILLER_16_2426 ();
 sg13g2_decap_4 FILLER_16_2454 ();
 sg13g2_fill_1 FILLER_16_2458 ();
 sg13g2_fill_2 FILLER_16_2463 ();
 sg13g2_fill_2 FILLER_16_2475 ();
 sg13g2_fill_1 FILLER_16_2477 ();
 sg13g2_decap_8 FILLER_16_2544 ();
 sg13g2_decap_8 FILLER_16_2551 ();
 sg13g2_decap_8 FILLER_16_2558 ();
 sg13g2_decap_8 FILLER_16_2565 ();
 sg13g2_decap_8 FILLER_16_2572 ();
 sg13g2_decap_8 FILLER_16_2579 ();
 sg13g2_decap_8 FILLER_16_2586 ();
 sg13g2_decap_8 FILLER_16_2593 ();
 sg13g2_decap_8 FILLER_16_2600 ();
 sg13g2_decap_8 FILLER_16_2607 ();
 sg13g2_decap_8 FILLER_16_2614 ();
 sg13g2_decap_8 FILLER_16_2621 ();
 sg13g2_decap_8 FILLER_16_2628 ();
 sg13g2_decap_8 FILLER_16_2635 ();
 sg13g2_decap_8 FILLER_16_2642 ();
 sg13g2_decap_8 FILLER_16_2649 ();
 sg13g2_decap_8 FILLER_16_2656 ();
 sg13g2_decap_8 FILLER_16_2663 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_31 ();
 sg13g2_decap_8 FILLER_17_38 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_decap_8 FILLER_17_80 ();
 sg13g2_decap_8 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_decap_8 FILLER_17_104 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_125 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_decap_4 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_decap_4 FILLER_17_247 ();
 sg13g2_decap_4 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_4 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_17_411 ();
 sg13g2_fill_1 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_431 ();
 sg13g2_fill_2 FILLER_17_459 ();
 sg13g2_fill_1 FILLER_17_487 ();
 sg13g2_fill_2 FILLER_17_514 ();
 sg13g2_fill_1 FILLER_17_537 ();
 sg13g2_fill_1 FILLER_17_547 ();
 sg13g2_fill_2 FILLER_17_552 ();
 sg13g2_fill_1 FILLER_17_559 ();
 sg13g2_fill_1 FILLER_17_565 ();
 sg13g2_decap_4 FILLER_17_592 ();
 sg13g2_fill_1 FILLER_17_596 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_fill_2 FILLER_17_689 ();
 sg13g2_fill_1 FILLER_17_696 ();
 sg13g2_fill_1 FILLER_17_707 ();
 sg13g2_fill_1 FILLER_17_712 ();
 sg13g2_fill_1 FILLER_17_753 ();
 sg13g2_fill_2 FILLER_17_762 ();
 sg13g2_fill_1 FILLER_17_764 ();
 sg13g2_decap_8 FILLER_17_773 ();
 sg13g2_fill_1 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_794 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_4 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_fill_2 FILLER_17_836 ();
 sg13g2_fill_1 FILLER_17_838 ();
 sg13g2_decap_8 FILLER_17_874 ();
 sg13g2_decap_8 FILLER_17_881 ();
 sg13g2_decap_8 FILLER_17_888 ();
 sg13g2_decap_4 FILLER_17_895 ();
 sg13g2_decap_8 FILLER_17_908 ();
 sg13g2_decap_8 FILLER_17_915 ();
 sg13g2_decap_8 FILLER_17_922 ();
 sg13g2_fill_1 FILLER_17_929 ();
 sg13g2_fill_1 FILLER_17_934 ();
 sg13g2_fill_1 FILLER_17_943 ();
 sg13g2_fill_2 FILLER_17_948 ();
 sg13g2_decap_4 FILLER_17_967 ();
 sg13g2_fill_1 FILLER_17_971 ();
 sg13g2_fill_1 FILLER_17_979 ();
 sg13g2_fill_2 FILLER_17_989 ();
 sg13g2_decap_8 FILLER_17_997 ();
 sg13g2_fill_1 FILLER_17_1004 ();
 sg13g2_decap_8 FILLER_17_1010 ();
 sg13g2_decap_8 FILLER_17_1017 ();
 sg13g2_decap_4 FILLER_17_1024 ();
 sg13g2_fill_2 FILLER_17_1028 ();
 sg13g2_decap_4 FILLER_17_1035 ();
 sg13g2_fill_2 FILLER_17_1039 ();
 sg13g2_decap_8 FILLER_17_1067 ();
 sg13g2_decap_4 FILLER_17_1074 ();
 sg13g2_fill_1 FILLER_17_1078 ();
 sg13g2_fill_1 FILLER_17_1084 ();
 sg13g2_fill_2 FILLER_17_1089 ();
 sg13g2_fill_1 FILLER_17_1091 ();
 sg13g2_fill_2 FILLER_17_1127 ();
 sg13g2_fill_2 FILLER_17_1141 ();
 sg13g2_fill_1 FILLER_17_1174 ();
 sg13g2_fill_2 FILLER_17_1184 ();
 sg13g2_decap_8 FILLER_17_1226 ();
 sg13g2_fill_1 FILLER_17_1233 ();
 sg13g2_fill_2 FILLER_17_1274 ();
 sg13g2_fill_2 FILLER_17_1302 ();
 sg13g2_fill_1 FILLER_17_1304 ();
 sg13g2_fill_2 FILLER_17_1336 ();
 sg13g2_fill_1 FILLER_17_1338 ();
 sg13g2_decap_8 FILLER_17_1343 ();
 sg13g2_decap_8 FILLER_17_1350 ();
 sg13g2_fill_2 FILLER_17_1357 ();
 sg13g2_decap_4 FILLER_17_1369 ();
 sg13g2_fill_1 FILLER_17_1373 ();
 sg13g2_fill_2 FILLER_17_1408 ();
 sg13g2_fill_1 FILLER_17_1416 ();
 sg13g2_fill_2 FILLER_17_1426 ();
 sg13g2_fill_2 FILLER_17_1464 ();
 sg13g2_decap_8 FILLER_17_1474 ();
 sg13g2_decap_8 FILLER_17_1481 ();
 sg13g2_decap_8 FILLER_17_1488 ();
 sg13g2_decap_8 FILLER_17_1495 ();
 sg13g2_decap_8 FILLER_17_1502 ();
 sg13g2_decap_4 FILLER_17_1509 ();
 sg13g2_decap_4 FILLER_17_1517 ();
 sg13g2_fill_1 FILLER_17_1521 ();
 sg13g2_decap_4 FILLER_17_1553 ();
 sg13g2_fill_1 FILLER_17_1583 ();
 sg13g2_fill_2 FILLER_17_1596 ();
 sg13g2_fill_1 FILLER_17_1607 ();
 sg13g2_fill_2 FILLER_17_1613 ();
 sg13g2_decap_8 FILLER_17_1619 ();
 sg13g2_fill_2 FILLER_17_1626 ();
 sg13g2_fill_1 FILLER_17_1628 ();
 sg13g2_fill_1 FILLER_17_1635 ();
 sg13g2_fill_2 FILLER_17_1650 ();
 sg13g2_fill_1 FILLER_17_1661 ();
 sg13g2_decap_8 FILLER_17_1667 ();
 sg13g2_decap_4 FILLER_17_1674 ();
 sg13g2_fill_2 FILLER_17_1692 ();
 sg13g2_decap_8 FILLER_17_1720 ();
 sg13g2_decap_8 FILLER_17_1727 ();
 sg13g2_decap_4 FILLER_17_1734 ();
 sg13g2_decap_8 FILLER_17_1747 ();
 sg13g2_decap_8 FILLER_17_1754 ();
 sg13g2_decap_8 FILLER_17_1761 ();
 sg13g2_decap_8 FILLER_17_1768 ();
 sg13g2_decap_4 FILLER_17_1775 ();
 sg13g2_fill_2 FILLER_17_1784 ();
 sg13g2_fill_1 FILLER_17_1789 ();
 sg13g2_fill_1 FILLER_17_1798 ();
 sg13g2_decap_8 FILLER_17_1834 ();
 sg13g2_decap_8 FILLER_17_1854 ();
 sg13g2_fill_2 FILLER_17_1861 ();
 sg13g2_decap_8 FILLER_17_1889 ();
 sg13g2_decap_8 FILLER_17_1896 ();
 sg13g2_decap_8 FILLER_17_1903 ();
 sg13g2_fill_1 FILLER_17_1910 ();
 sg13g2_decap_4 FILLER_17_1916 ();
 sg13g2_fill_1 FILLER_17_1920 ();
 sg13g2_fill_2 FILLER_17_1925 ();
 sg13g2_decap_4 FILLER_17_1933 ();
 sg13g2_fill_2 FILLER_17_1937 ();
 sg13g2_decap_8 FILLER_17_1942 ();
 sg13g2_decap_4 FILLER_17_1949 ();
 sg13g2_fill_2 FILLER_17_1953 ();
 sg13g2_decap_4 FILLER_17_1960 ();
 sg13g2_fill_1 FILLER_17_1964 ();
 sg13g2_decap_8 FILLER_17_1969 ();
 sg13g2_decap_8 FILLER_17_1976 ();
 sg13g2_fill_2 FILLER_17_1983 ();
 sg13g2_fill_1 FILLER_17_1998 ();
 sg13g2_fill_1 FILLER_17_2003 ();
 sg13g2_decap_4 FILLER_17_2010 ();
 sg13g2_decap_8 FILLER_17_2044 ();
 sg13g2_decap_8 FILLER_17_2051 ();
 sg13g2_decap_4 FILLER_17_2058 ();
 sg13g2_fill_2 FILLER_17_2062 ();
 sg13g2_decap_8 FILLER_17_2099 ();
 sg13g2_decap_8 FILLER_17_2106 ();
 sg13g2_decap_8 FILLER_17_2113 ();
 sg13g2_decap_4 FILLER_17_2125 ();
 sg13g2_fill_2 FILLER_17_2129 ();
 sg13g2_fill_1 FILLER_17_2135 ();
 sg13g2_fill_1 FILLER_17_2162 ();
 sg13g2_fill_1 FILLER_17_2182 ();
 sg13g2_fill_1 FILLER_17_2193 ();
 sg13g2_decap_8 FILLER_17_2250 ();
 sg13g2_decap_8 FILLER_17_2257 ();
 sg13g2_decap_8 FILLER_17_2264 ();
 sg13g2_decap_8 FILLER_17_2271 ();
 sg13g2_decap_8 FILLER_17_2278 ();
 sg13g2_decap_8 FILLER_17_2285 ();
 sg13g2_decap_8 FILLER_17_2292 ();
 sg13g2_decap_4 FILLER_17_2304 ();
 sg13g2_fill_1 FILLER_17_2347 ();
 sg13g2_fill_1 FILLER_17_2357 ();
 sg13g2_decap_4 FILLER_17_2418 ();
 sg13g2_fill_1 FILLER_17_2422 ();
 sg13g2_decap_8 FILLER_17_2453 ();
 sg13g2_decap_8 FILLER_17_2460 ();
 sg13g2_decap_4 FILLER_17_2467 ();
 sg13g2_fill_1 FILLER_17_2471 ();
 sg13g2_fill_2 FILLER_17_2482 ();
 sg13g2_fill_1 FILLER_17_2488 ();
 sg13g2_decap_8 FILLER_17_2506 ();
 sg13g2_decap_8 FILLER_17_2543 ();
 sg13g2_decap_8 FILLER_17_2550 ();
 sg13g2_decap_8 FILLER_17_2557 ();
 sg13g2_decap_8 FILLER_17_2564 ();
 sg13g2_decap_8 FILLER_17_2571 ();
 sg13g2_decap_8 FILLER_17_2578 ();
 sg13g2_decap_8 FILLER_17_2585 ();
 sg13g2_decap_8 FILLER_17_2592 ();
 sg13g2_decap_8 FILLER_17_2599 ();
 sg13g2_decap_8 FILLER_17_2606 ();
 sg13g2_decap_8 FILLER_17_2613 ();
 sg13g2_decap_8 FILLER_17_2620 ();
 sg13g2_decap_8 FILLER_17_2627 ();
 sg13g2_decap_8 FILLER_17_2634 ();
 sg13g2_decap_8 FILLER_17_2641 ();
 sg13g2_decap_8 FILLER_17_2648 ();
 sg13g2_decap_8 FILLER_17_2655 ();
 sg13g2_decap_8 FILLER_17_2662 ();
 sg13g2_fill_1 FILLER_17_2669 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_decap_4 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_111 ();
 sg13g2_decap_4 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_4 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_decap_4 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_decap_4 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_4 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_decap_4 FILLER_18_413 ();
 sg13g2_decap_4 FILLER_18_423 ();
 sg13g2_fill_2 FILLER_18_437 ();
 sg13g2_fill_1 FILLER_18_439 ();
 sg13g2_fill_2 FILLER_18_444 ();
 sg13g2_fill_1 FILLER_18_446 ();
 sg13g2_fill_1 FILLER_18_457 ();
 sg13g2_decap_8 FILLER_18_492 ();
 sg13g2_fill_1 FILLER_18_499 ();
 sg13g2_fill_1 FILLER_18_539 ();
 sg13g2_fill_1 FILLER_18_543 ();
 sg13g2_fill_2 FILLER_18_557 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_fill_1 FILLER_18_581 ();
 sg13g2_fill_2 FILLER_18_611 ();
 sg13g2_fill_1 FILLER_18_613 ();
 sg13g2_fill_1 FILLER_18_644 ();
 sg13g2_fill_2 FILLER_18_661 ();
 sg13g2_fill_1 FILLER_18_692 ();
 sg13g2_fill_1 FILLER_18_727 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_fill_1 FILLER_18_739 ();
 sg13g2_decap_4 FILLER_18_758 ();
 sg13g2_fill_1 FILLER_18_762 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_fill_1 FILLER_18_775 ();
 sg13g2_fill_2 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_fill_2 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_fill_1 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_948 ();
 sg13g2_decap_4 FILLER_18_955 ();
 sg13g2_decap_8 FILLER_18_963 ();
 sg13g2_fill_2 FILLER_18_970 ();
 sg13g2_decap_8 FILLER_18_981 ();
 sg13g2_decap_8 FILLER_18_988 ();
 sg13g2_fill_1 FILLER_18_995 ();
 sg13g2_fill_2 FILLER_18_1027 ();
 sg13g2_fill_1 FILLER_18_1029 ();
 sg13g2_fill_2 FILLER_18_1034 ();
 sg13g2_fill_1 FILLER_18_1036 ();
 sg13g2_decap_4 FILLER_18_1042 ();
 sg13g2_decap_8 FILLER_18_1054 ();
 sg13g2_decap_8 FILLER_18_1061 ();
 sg13g2_decap_8 FILLER_18_1068 ();
 sg13g2_decap_8 FILLER_18_1075 ();
 sg13g2_fill_1 FILLER_18_1082 ();
 sg13g2_fill_2 FILLER_18_1089 ();
 sg13g2_decap_8 FILLER_18_1099 ();
 sg13g2_decap_4 FILLER_18_1106 ();
 sg13g2_fill_1 FILLER_18_1110 ();
 sg13g2_fill_2 FILLER_18_1143 ();
 sg13g2_fill_1 FILLER_18_1160 ();
 sg13g2_fill_2 FILLER_18_1187 ();
 sg13g2_fill_2 FILLER_18_1218 ();
 sg13g2_fill_2 FILLER_18_1225 ();
 sg13g2_fill_1 FILLER_18_1227 ();
 sg13g2_decap_8 FILLER_18_1237 ();
 sg13g2_fill_2 FILLER_18_1244 ();
 sg13g2_decap_4 FILLER_18_1252 ();
 sg13g2_fill_1 FILLER_18_1256 ();
 sg13g2_decap_4 FILLER_18_1263 ();
 sg13g2_decap_8 FILLER_18_1275 ();
 sg13g2_decap_4 FILLER_18_1282 ();
 sg13g2_decap_8 FILLER_18_1304 ();
 sg13g2_decap_8 FILLER_18_1311 ();
 sg13g2_fill_1 FILLER_18_1323 ();
 sg13g2_decap_4 FILLER_18_1374 ();
 sg13g2_fill_1 FILLER_18_1378 ();
 sg13g2_fill_2 FILLER_18_1395 ();
 sg13g2_fill_2 FILLER_18_1428 ();
 sg13g2_decap_4 FILLER_18_1471 ();
 sg13g2_fill_2 FILLER_18_1505 ();
 sg13g2_fill_1 FILLER_18_1507 ();
 sg13g2_fill_1 FILLER_18_1513 ();
 sg13g2_decap_8 FILLER_18_1527 ();
 sg13g2_decap_8 FILLER_18_1563 ();
 sg13g2_fill_2 FILLER_18_1570 ();
 sg13g2_decap_8 FILLER_18_1616 ();
 sg13g2_fill_2 FILLER_18_1623 ();
 sg13g2_fill_1 FILLER_18_1625 ();
 sg13g2_fill_2 FILLER_18_1665 ();
 sg13g2_decap_8 FILLER_18_1719 ();
 sg13g2_decap_4 FILLER_18_1726 ();
 sg13g2_fill_2 FILLER_18_1730 ();
 sg13g2_fill_2 FILLER_18_1781 ();
 sg13g2_fill_2 FILLER_18_1794 ();
 sg13g2_fill_2 FILLER_18_1822 ();
 sg13g2_fill_1 FILLER_18_1824 ();
 sg13g2_fill_1 FILLER_18_1830 ();
 sg13g2_fill_2 FILLER_18_1857 ();
 sg13g2_fill_1 FILLER_18_1859 ();
 sg13g2_decap_8 FILLER_18_1866 ();
 sg13g2_decap_8 FILLER_18_1873 ();
 sg13g2_fill_2 FILLER_18_1880 ();
 sg13g2_fill_1 FILLER_18_1891 ();
 sg13g2_decap_4 FILLER_18_1918 ();
 sg13g2_fill_2 FILLER_18_1928 ();
 sg13g2_decap_8 FILLER_18_1938 ();
 sg13g2_fill_1 FILLER_18_1945 ();
 sg13g2_fill_1 FILLER_18_1954 ();
 sg13g2_fill_2 FILLER_18_1963 ();
 sg13g2_fill_1 FILLER_18_1974 ();
 sg13g2_fill_1 FILLER_18_2001 ();
 sg13g2_fill_2 FILLER_18_2036 ();
 sg13g2_fill_1 FILLER_18_2038 ();
 sg13g2_decap_8 FILLER_18_2043 ();
 sg13g2_decap_4 FILLER_18_2050 ();
 sg13g2_fill_2 FILLER_18_2054 ();
 sg13g2_decap_8 FILLER_18_2061 ();
 sg13g2_decap_8 FILLER_18_2103 ();
 sg13g2_fill_1 FILLER_18_2110 ();
 sg13g2_decap_4 FILLER_18_2116 ();
 sg13g2_fill_1 FILLER_18_2120 ();
 sg13g2_decap_8 FILLER_18_2183 ();
 sg13g2_fill_2 FILLER_18_2196 ();
 sg13g2_fill_1 FILLER_18_2261 ();
 sg13g2_fill_1 FILLER_18_2268 ();
 sg13g2_decap_4 FILLER_18_2273 ();
 sg13g2_fill_1 FILLER_18_2277 ();
 sg13g2_fill_2 FILLER_18_2304 ();
 sg13g2_decap_8 FILLER_18_2310 ();
 sg13g2_fill_1 FILLER_18_2317 ();
 sg13g2_fill_1 FILLER_18_2370 ();
 sg13g2_fill_1 FILLER_18_2374 ();
 sg13g2_fill_1 FILLER_18_2383 ();
 sg13g2_decap_8 FILLER_18_2406 ();
 sg13g2_decap_8 FILLER_18_2413 ();
 sg13g2_decap_8 FILLER_18_2420 ();
 sg13g2_decap_4 FILLER_18_2427 ();
 sg13g2_fill_2 FILLER_18_2431 ();
 sg13g2_fill_1 FILLER_18_2437 ();
 sg13g2_decap_8 FILLER_18_2442 ();
 sg13g2_decap_8 FILLER_18_2449 ();
 sg13g2_decap_8 FILLER_18_2456 ();
 sg13g2_fill_2 FILLER_18_2463 ();
 sg13g2_fill_1 FILLER_18_2465 ();
 sg13g2_fill_2 FILLER_18_2472 ();
 sg13g2_fill_1 FILLER_18_2482 ();
 sg13g2_fill_1 FILLER_18_2509 ();
 sg13g2_decap_8 FILLER_18_2514 ();
 sg13g2_fill_2 FILLER_18_2521 ();
 sg13g2_fill_1 FILLER_18_2523 ();
 sg13g2_decap_8 FILLER_18_2528 ();
 sg13g2_decap_8 FILLER_18_2535 ();
 sg13g2_decap_8 FILLER_18_2542 ();
 sg13g2_decap_8 FILLER_18_2549 ();
 sg13g2_decap_8 FILLER_18_2556 ();
 sg13g2_decap_8 FILLER_18_2563 ();
 sg13g2_decap_8 FILLER_18_2570 ();
 sg13g2_decap_8 FILLER_18_2577 ();
 sg13g2_decap_8 FILLER_18_2584 ();
 sg13g2_decap_8 FILLER_18_2591 ();
 sg13g2_decap_8 FILLER_18_2598 ();
 sg13g2_decap_8 FILLER_18_2605 ();
 sg13g2_decap_8 FILLER_18_2612 ();
 sg13g2_decap_8 FILLER_18_2619 ();
 sg13g2_decap_8 FILLER_18_2626 ();
 sg13g2_decap_8 FILLER_18_2633 ();
 sg13g2_decap_8 FILLER_18_2640 ();
 sg13g2_decap_8 FILLER_18_2647 ();
 sg13g2_decap_8 FILLER_18_2654 ();
 sg13g2_decap_8 FILLER_18_2661 ();
 sg13g2_fill_2 FILLER_18_2668 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_69 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_171 ();
 sg13g2_decap_4 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_4 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_290 ();
 sg13g2_decap_4 FILLER_19_297 ();
 sg13g2_decap_4 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_decap_4 FILLER_19_324 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_1 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_376 ();
 sg13g2_decap_4 FILLER_19_386 ();
 sg13g2_fill_2 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_436 ();
 sg13g2_fill_2 FILLER_19_440 ();
 sg13g2_fill_2 FILLER_19_475 ();
 sg13g2_fill_1 FILLER_19_477 ();
 sg13g2_decap_8 FILLER_19_482 ();
 sg13g2_decap_8 FILLER_19_576 ();
 sg13g2_decap_8 FILLER_19_583 ();
 sg13g2_decap_4 FILLER_19_590 ();
 sg13g2_fill_1 FILLER_19_613 ();
 sg13g2_fill_1 FILLER_19_619 ();
 sg13g2_fill_1 FILLER_19_640 ();
 sg13g2_fill_2 FILLER_19_657 ();
 sg13g2_fill_2 FILLER_19_685 ();
 sg13g2_fill_1 FILLER_19_687 ();
 sg13g2_fill_2 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_730 ();
 sg13g2_decap_8 FILLER_19_737 ();
 sg13g2_decap_8 FILLER_19_744 ();
 sg13g2_decap_8 FILLER_19_751 ();
 sg13g2_decap_8 FILLER_19_758 ();
 sg13g2_decap_8 FILLER_19_765 ();
 sg13g2_fill_2 FILLER_19_772 ();
 sg13g2_fill_1 FILLER_19_774 ();
 sg13g2_fill_1 FILLER_19_837 ();
 sg13g2_fill_1 FILLER_19_864 ();
 sg13g2_fill_1 FILLER_19_871 ();
 sg13g2_fill_1 FILLER_19_882 ();
 sg13g2_fill_1 FILLER_19_887 ();
 sg13g2_fill_1 FILLER_19_894 ();
 sg13g2_decap_4 FILLER_19_957 ();
 sg13g2_fill_1 FILLER_19_961 ();
 sg13g2_decap_4 FILLER_19_1030 ();
 sg13g2_decap_8 FILLER_19_1040 ();
 sg13g2_fill_2 FILLER_19_1047 ();
 sg13g2_decap_8 FILLER_19_1054 ();
 sg13g2_decap_4 FILLER_19_1061 ();
 sg13g2_decap_8 FILLER_19_1069 ();
 sg13g2_decap_8 FILLER_19_1076 ();
 sg13g2_decap_4 FILLER_19_1083 ();
 sg13g2_fill_2 FILLER_19_1087 ();
 sg13g2_decap_4 FILLER_19_1093 ();
 sg13g2_fill_1 FILLER_19_1097 ();
 sg13g2_decap_4 FILLER_19_1113 ();
 sg13g2_fill_2 FILLER_19_1126 ();
 sg13g2_fill_1 FILLER_19_1128 ();
 sg13g2_fill_1 FILLER_19_1143 ();
 sg13g2_fill_1 FILLER_19_1187 ();
 sg13g2_fill_2 FILLER_19_1205 ();
 sg13g2_fill_1 FILLER_19_1223 ();
 sg13g2_fill_2 FILLER_19_1261 ();
 sg13g2_fill_1 FILLER_19_1263 ();
 sg13g2_decap_8 FILLER_19_1269 ();
 sg13g2_fill_2 FILLER_19_1276 ();
 sg13g2_fill_1 FILLER_19_1278 ();
 sg13g2_decap_8 FILLER_19_1284 ();
 sg13g2_decap_8 FILLER_19_1291 ();
 sg13g2_decap_8 FILLER_19_1298 ();
 sg13g2_decap_8 FILLER_19_1305 ();
 sg13g2_decap_8 FILLER_19_1312 ();
 sg13g2_fill_1 FILLER_19_1319 ();
 sg13g2_fill_1 FILLER_19_1351 ();
 sg13g2_fill_2 FILLER_19_1370 ();
 sg13g2_fill_1 FILLER_19_1372 ();
 sg13g2_fill_2 FILLER_19_1378 ();
 sg13g2_fill_2 FILLER_19_1430 ();
 sg13g2_fill_2 FILLER_19_1439 ();
 sg13g2_decap_4 FILLER_19_1472 ();
 sg13g2_fill_1 FILLER_19_1476 ();
 sg13g2_fill_1 FILLER_19_1507 ();
 sg13g2_fill_1 FILLER_19_1512 ();
 sg13g2_fill_1 FILLER_19_1518 ();
 sg13g2_decap_8 FILLER_19_1545 ();
 sg13g2_fill_1 FILLER_19_1552 ();
 sg13g2_decap_8 FILLER_19_1569 ();
 sg13g2_decap_8 FILLER_19_1576 ();
 sg13g2_decap_8 FILLER_19_1589 ();
 sg13g2_fill_2 FILLER_19_1596 ();
 sg13g2_decap_4 FILLER_19_1611 ();
 sg13g2_fill_1 FILLER_19_1615 ();
 sg13g2_fill_1 FILLER_19_1642 ();
 sg13g2_fill_1 FILLER_19_1690 ();
 sg13g2_fill_2 FILLER_19_1696 ();
 sg13g2_decap_4 FILLER_19_1703 ();
 sg13g2_fill_1 FILLER_19_1707 ();
 sg13g2_fill_2 FILLER_19_1721 ();
 sg13g2_fill_2 FILLER_19_1749 ();
 sg13g2_decap_4 FILLER_19_1755 ();
 sg13g2_fill_1 FILLER_19_1759 ();
 sg13g2_fill_2 FILLER_19_1790 ();
 sg13g2_fill_2 FILLER_19_1797 ();
 sg13g2_fill_1 FILLER_19_1799 ();
 sg13g2_decap_4 FILLER_19_1831 ();
 sg13g2_fill_2 FILLER_19_1848 ();
 sg13g2_fill_2 FILLER_19_1876 ();
 sg13g2_fill_2 FILLER_19_1883 ();
 sg13g2_fill_2 FILLER_19_1900 ();
 sg13g2_fill_1 FILLER_19_1902 ();
 sg13g2_fill_2 FILLER_19_1908 ();
 sg13g2_fill_1 FILLER_19_1910 ();
 sg13g2_decap_4 FILLER_19_1916 ();
 sg13g2_fill_2 FILLER_19_1924 ();
 sg13g2_fill_1 FILLER_19_1930 ();
 sg13g2_decap_8 FILLER_19_1937 ();
 sg13g2_decap_8 FILLER_19_1944 ();
 sg13g2_decap_4 FILLER_19_1951 ();
 sg13g2_decap_8 FILLER_19_1960 ();
 sg13g2_fill_2 FILLER_19_1967 ();
 sg13g2_decap_8 FILLER_19_1973 ();
 sg13g2_decap_8 FILLER_19_1980 ();
 sg13g2_decap_8 FILLER_19_1987 ();
 sg13g2_decap_8 FILLER_19_1994 ();
 sg13g2_decap_4 FILLER_19_2001 ();
 sg13g2_fill_1 FILLER_19_2005 ();
 sg13g2_fill_2 FILLER_19_2026 ();
 sg13g2_decap_8 FILLER_19_2032 ();
 sg13g2_decap_8 FILLER_19_2039 ();
 sg13g2_decap_4 FILLER_19_2046 ();
 sg13g2_fill_1 FILLER_19_2050 ();
 sg13g2_fill_2 FILLER_19_2085 ();
 sg13g2_decap_4 FILLER_19_2091 ();
 sg13g2_decap_4 FILLER_19_2121 ();
 sg13g2_fill_2 FILLER_19_2125 ();
 sg13g2_fill_2 FILLER_19_2142 ();
 sg13g2_fill_1 FILLER_19_2144 ();
 sg13g2_fill_1 FILLER_19_2148 ();
 sg13g2_fill_2 FILLER_19_2155 ();
 sg13g2_fill_1 FILLER_19_2157 ();
 sg13g2_fill_1 FILLER_19_2162 ();
 sg13g2_decap_8 FILLER_19_2169 ();
 sg13g2_decap_8 FILLER_19_2176 ();
 sg13g2_fill_1 FILLER_19_2183 ();
 sg13g2_fill_2 FILLER_19_2199 ();
 sg13g2_fill_2 FILLER_19_2237 ();
 sg13g2_fill_2 FILLER_19_2265 ();
 sg13g2_fill_1 FILLER_19_2298 ();
 sg13g2_fill_2 FILLER_19_2350 ();
 sg13g2_decap_8 FILLER_19_2386 ();
 sg13g2_decap_4 FILLER_19_2393 ();
 sg13g2_fill_1 FILLER_19_2397 ();
 sg13g2_decap_8 FILLER_19_2424 ();
 sg13g2_fill_2 FILLER_19_2431 ();
 sg13g2_fill_1 FILLER_19_2433 ();
 sg13g2_decap_8 FILLER_19_2438 ();
 sg13g2_decap_8 FILLER_19_2445 ();
 sg13g2_decap_8 FILLER_19_2452 ();
 sg13g2_fill_2 FILLER_19_2459 ();
 sg13g2_decap_8 FILLER_19_2465 ();
 sg13g2_fill_2 FILLER_19_2478 ();
 sg13g2_decap_4 FILLER_19_2509 ();
 sg13g2_decap_8 FILLER_19_2539 ();
 sg13g2_decap_8 FILLER_19_2546 ();
 sg13g2_decap_8 FILLER_19_2553 ();
 sg13g2_decap_8 FILLER_19_2560 ();
 sg13g2_decap_8 FILLER_19_2567 ();
 sg13g2_decap_8 FILLER_19_2574 ();
 sg13g2_decap_8 FILLER_19_2581 ();
 sg13g2_decap_8 FILLER_19_2588 ();
 sg13g2_decap_8 FILLER_19_2595 ();
 sg13g2_decap_8 FILLER_19_2602 ();
 sg13g2_decap_8 FILLER_19_2609 ();
 sg13g2_decap_8 FILLER_19_2616 ();
 sg13g2_decap_8 FILLER_19_2623 ();
 sg13g2_decap_8 FILLER_19_2630 ();
 sg13g2_decap_8 FILLER_19_2637 ();
 sg13g2_decap_8 FILLER_19_2644 ();
 sg13g2_decap_8 FILLER_19_2651 ();
 sg13g2_decap_8 FILLER_19_2658 ();
 sg13g2_decap_4 FILLER_19_2665 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_4 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_decap_4 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_4 FILLER_20_351 ();
 sg13g2_decap_4 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_fill_1 FILLER_20_401 ();
 sg13g2_decap_4 FILLER_20_412 ();
 sg13g2_fill_2 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_450 ();
 sg13g2_decap_4 FILLER_20_457 ();
 sg13g2_fill_2 FILLER_20_467 ();
 sg13g2_fill_1 FILLER_20_469 ();
 sg13g2_fill_2 FILLER_20_474 ();
 sg13g2_fill_1 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_fill_2 FILLER_20_524 ();
 sg13g2_fill_2 FILLER_20_532 ();
 sg13g2_decap_4 FILLER_20_578 ();
 sg13g2_fill_2 FILLER_20_582 ();
 sg13g2_decap_4 FILLER_20_589 ();
 sg13g2_fill_2 FILLER_20_593 ();
 sg13g2_fill_1 FILLER_20_601 ();
 sg13g2_decap_8 FILLER_20_608 ();
 sg13g2_fill_1 FILLER_20_615 ();
 sg13g2_fill_1 FILLER_20_625 ();
 sg13g2_decap_8 FILLER_20_634 ();
 sg13g2_fill_1 FILLER_20_641 ();
 sg13g2_decap_8 FILLER_20_647 ();
 sg13g2_fill_1 FILLER_20_654 ();
 sg13g2_fill_1 FILLER_20_660 ();
 sg13g2_fill_2 FILLER_20_666 ();
 sg13g2_decap_8 FILLER_20_673 ();
 sg13g2_fill_2 FILLER_20_680 ();
 sg13g2_decap_4 FILLER_20_687 ();
 sg13g2_decap_8 FILLER_20_725 ();
 sg13g2_decap_8 FILLER_20_732 ();
 sg13g2_fill_2 FILLER_20_769 ();
 sg13g2_fill_1 FILLER_20_771 ();
 sg13g2_fill_1 FILLER_20_828 ();
 sg13g2_fill_1 FILLER_20_839 ();
 sg13g2_fill_1 FILLER_20_844 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_fill_2 FILLER_20_892 ();
 sg13g2_fill_1 FILLER_20_894 ();
 sg13g2_fill_2 FILLER_20_919 ();
 sg13g2_fill_1 FILLER_20_925 ();
 sg13g2_fill_1 FILLER_20_939 ();
 sg13g2_decap_8 FILLER_20_944 ();
 sg13g2_fill_2 FILLER_20_951 ();
 sg13g2_decap_8 FILLER_20_958 ();
 sg13g2_fill_2 FILLER_20_965 ();
 sg13g2_fill_2 FILLER_20_999 ();
 sg13g2_fill_1 FILLER_20_1001 ();
 sg13g2_decap_4 FILLER_20_1042 ();
 sg13g2_fill_1 FILLER_20_1046 ();
 sg13g2_fill_2 FILLER_20_1053 ();
 sg13g2_decap_8 FILLER_20_1061 ();
 sg13g2_fill_1 FILLER_20_1068 ();
 sg13g2_decap_4 FILLER_20_1078 ();
 sg13g2_fill_2 FILLER_20_1102 ();
 sg13g2_decap_8 FILLER_20_1130 ();
 sg13g2_decap_8 FILLER_20_1137 ();
 sg13g2_decap_8 FILLER_20_1144 ();
 sg13g2_decap_4 FILLER_20_1151 ();
 sg13g2_fill_2 FILLER_20_1160 ();
 sg13g2_fill_1 FILLER_20_1162 ();
 sg13g2_decap_8 FILLER_20_1172 ();
 sg13g2_decap_8 FILLER_20_1179 ();
 sg13g2_fill_1 FILLER_20_1186 ();
 sg13g2_fill_1 FILLER_20_1195 ();
 sg13g2_fill_1 FILLER_20_1231 ();
 sg13g2_decap_8 FILLER_20_1237 ();
 sg13g2_fill_1 FILLER_20_1244 ();
 sg13g2_decap_8 FILLER_20_1275 ();
 sg13g2_decap_4 FILLER_20_1282 ();
 sg13g2_fill_2 FILLER_20_1286 ();
 sg13g2_fill_1 FILLER_20_1297 ();
 sg13g2_decap_8 FILLER_20_1314 ();
 sg13g2_decap_4 FILLER_20_1321 ();
 sg13g2_fill_1 FILLER_20_1325 ();
 sg13g2_fill_2 FILLER_20_1331 ();
 sg13g2_fill_1 FILLER_20_1333 ();
 sg13g2_fill_1 FILLER_20_1338 ();
 sg13g2_fill_1 FILLER_20_1343 ();
 sg13g2_decap_4 FILLER_20_1354 ();
 sg13g2_fill_2 FILLER_20_1371 ();
 sg13g2_decap_8 FILLER_20_1444 ();
 sg13g2_decap_8 FILLER_20_1451 ();
 sg13g2_decap_8 FILLER_20_1458 ();
 sg13g2_fill_2 FILLER_20_1465 ();
 sg13g2_fill_1 FILLER_20_1467 ();
 sg13g2_decap_4 FILLER_20_1473 ();
 sg13g2_fill_2 FILLER_20_1477 ();
 sg13g2_decap_8 FILLER_20_1492 ();
 sg13g2_decap_8 FILLER_20_1504 ();
 sg13g2_decap_8 FILLER_20_1511 ();
 sg13g2_fill_2 FILLER_20_1518 ();
 sg13g2_fill_1 FILLER_20_1520 ();
 sg13g2_fill_1 FILLER_20_1562 ();
 sg13g2_fill_2 FILLER_20_1616 ();
 sg13g2_fill_2 FILLER_20_1653 ();
 sg13g2_decap_8 FILLER_20_1681 ();
 sg13g2_decap_4 FILLER_20_1688 ();
 sg13g2_fill_2 FILLER_20_1692 ();
 sg13g2_decap_8 FILLER_20_1707 ();
 sg13g2_fill_1 FILLER_20_1714 ();
 sg13g2_fill_2 FILLER_20_1741 ();
 sg13g2_fill_1 FILLER_20_1743 ();
 sg13g2_decap_4 FILLER_20_1748 ();
 sg13g2_fill_1 FILLER_20_1752 ();
 sg13g2_fill_2 FILLER_20_1772 ();
 sg13g2_decap_8 FILLER_20_1778 ();
 sg13g2_decap_8 FILLER_20_1785 ();
 sg13g2_decap_4 FILLER_20_1792 ();
 sg13g2_fill_2 FILLER_20_1796 ();
 sg13g2_decap_8 FILLER_20_1803 ();
 sg13g2_fill_2 FILLER_20_1810 ();
 sg13g2_decap_8 FILLER_20_1822 ();
 sg13g2_fill_2 FILLER_20_1829 ();
 sg13g2_fill_1 FILLER_20_1852 ();
 sg13g2_fill_1 FILLER_20_1859 ();
 sg13g2_fill_2 FILLER_20_1866 ();
 sg13g2_fill_1 FILLER_20_1873 ();
 sg13g2_fill_1 FILLER_20_1878 ();
 sg13g2_fill_1 FILLER_20_1885 ();
 sg13g2_fill_1 FILLER_20_1891 ();
 sg13g2_fill_2 FILLER_20_1956 ();
 sg13g2_fill_1 FILLER_20_1963 ();
 sg13g2_fill_2 FILLER_20_1968 ();
 sg13g2_fill_1 FILLER_20_1970 ();
 sg13g2_fill_2 FILLER_20_1975 ();
 sg13g2_fill_2 FILLER_20_1987 ();
 sg13g2_fill_1 FILLER_20_1989 ();
 sg13g2_decap_8 FILLER_20_1993 ();
 sg13g2_decap_8 FILLER_20_2000 ();
 sg13g2_fill_1 FILLER_20_2012 ();
 sg13g2_decap_8 FILLER_20_2026 ();
 sg13g2_decap_8 FILLER_20_2033 ();
 sg13g2_decap_8 FILLER_20_2040 ();
 sg13g2_decap_8 FILLER_20_2047 ();
 sg13g2_decap_8 FILLER_20_2059 ();
 sg13g2_decap_8 FILLER_20_2066 ();
 sg13g2_decap_8 FILLER_20_2073 ();
 sg13g2_decap_4 FILLER_20_2080 ();
 sg13g2_fill_2 FILLER_20_2084 ();
 sg13g2_fill_1 FILLER_20_2104 ();
 sg13g2_fill_2 FILLER_20_2109 ();
 sg13g2_decap_8 FILLER_20_2174 ();
 sg13g2_decap_4 FILLER_20_2181 ();
 sg13g2_fill_1 FILLER_20_2185 ();
 sg13g2_fill_1 FILLER_20_2225 ();
 sg13g2_fill_1 FILLER_20_2265 ();
 sg13g2_fill_1 FILLER_20_2292 ();
 sg13g2_decap_8 FILLER_20_2315 ();
 sg13g2_fill_1 FILLER_20_2328 ();
 sg13g2_decap_4 FILLER_20_2367 ();
 sg13g2_fill_2 FILLER_20_2371 ();
 sg13g2_decap_8 FILLER_20_2376 ();
 sg13g2_decap_8 FILLER_20_2383 ();
 sg13g2_decap_4 FILLER_20_2390 ();
 sg13g2_decap_8 FILLER_20_2420 ();
 sg13g2_decap_8 FILLER_20_2427 ();
 sg13g2_decap_4 FILLER_20_2434 ();
 sg13g2_fill_2 FILLER_20_2438 ();
 sg13g2_decap_8 FILLER_20_2444 ();
 sg13g2_decap_4 FILLER_20_2485 ();
 sg13g2_fill_1 FILLER_20_2494 ();
 sg13g2_decap_4 FILLER_20_2499 ();
 sg13g2_decap_8 FILLER_20_2516 ();
 sg13g2_decap_8 FILLER_20_2523 ();
 sg13g2_decap_8 FILLER_20_2530 ();
 sg13g2_decap_8 FILLER_20_2537 ();
 sg13g2_decap_8 FILLER_20_2544 ();
 sg13g2_decap_8 FILLER_20_2551 ();
 sg13g2_decap_8 FILLER_20_2558 ();
 sg13g2_decap_8 FILLER_20_2565 ();
 sg13g2_decap_8 FILLER_20_2572 ();
 sg13g2_decap_8 FILLER_20_2579 ();
 sg13g2_decap_8 FILLER_20_2586 ();
 sg13g2_decap_8 FILLER_20_2593 ();
 sg13g2_decap_8 FILLER_20_2600 ();
 sg13g2_decap_8 FILLER_20_2607 ();
 sg13g2_decap_8 FILLER_20_2614 ();
 sg13g2_decap_8 FILLER_20_2621 ();
 sg13g2_decap_8 FILLER_20_2628 ();
 sg13g2_decap_8 FILLER_20_2635 ();
 sg13g2_decap_8 FILLER_20_2642 ();
 sg13g2_decap_8 FILLER_20_2649 ();
 sg13g2_decap_8 FILLER_20_2656 ();
 sg13g2_decap_8 FILLER_20_2663 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_decap_4 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_371 ();
 sg13g2_decap_4 FILLER_21_385 ();
 sg13g2_decap_4 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_fill_2 FILLER_21_417 ();
 sg13g2_fill_1 FILLER_21_419 ();
 sg13g2_fill_2 FILLER_21_439 ();
 sg13g2_fill_1 FILLER_21_441 ();
 sg13g2_fill_1 FILLER_21_452 ();
 sg13g2_decap_8 FILLER_21_456 ();
 sg13g2_fill_2 FILLER_21_463 ();
 sg13g2_fill_2 FILLER_21_468 ();
 sg13g2_fill_1 FILLER_21_470 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_fill_2 FILLER_21_511 ();
 sg13g2_fill_1 FILLER_21_513 ();
 sg13g2_fill_1 FILLER_21_546 ();
 sg13g2_fill_2 FILLER_21_559 ();
 sg13g2_decap_4 FILLER_21_570 ();
 sg13g2_fill_2 FILLER_21_574 ();
 sg13g2_fill_1 FILLER_21_597 ();
 sg13g2_fill_2 FILLER_21_610 ();
 sg13g2_decap_8 FILLER_21_621 ();
 sg13g2_fill_1 FILLER_21_643 ();
 sg13g2_fill_2 FILLER_21_657 ();
 sg13g2_decap_8 FILLER_21_662 ();
 sg13g2_decap_8 FILLER_21_669 ();
 sg13g2_decap_8 FILLER_21_676 ();
 sg13g2_decap_8 FILLER_21_683 ();
 sg13g2_fill_1 FILLER_21_695 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_4 FILLER_21_762 ();
 sg13g2_fill_1 FILLER_21_766 ();
 sg13g2_fill_2 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_825 ();
 sg13g2_decap_4 FILLER_21_832 ();
 sg13g2_fill_1 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_841 ();
 sg13g2_decap_8 FILLER_21_848 ();
 sg13g2_decap_8 FILLER_21_859 ();
 sg13g2_decap_8 FILLER_21_866 ();
 sg13g2_fill_1 FILLER_21_873 ();
 sg13g2_decap_4 FILLER_21_878 ();
 sg13g2_fill_1 FILLER_21_933 ();
 sg13g2_fill_1 FILLER_21_964 ();
 sg13g2_fill_2 FILLER_21_970 ();
 sg13g2_decap_4 FILLER_21_981 ();
 sg13g2_fill_1 FILLER_21_985 ();
 sg13g2_fill_2 FILLER_21_994 ();
 sg13g2_decap_8 FILLER_21_1001 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_fill_2 FILLER_21_1015 ();
 sg13g2_fill_1 FILLER_21_1017 ();
 sg13g2_decap_8 FILLER_21_1029 ();
 sg13g2_decap_4 FILLER_21_1036 ();
 sg13g2_fill_2 FILLER_21_1040 ();
 sg13g2_fill_2 FILLER_21_1056 ();
 sg13g2_fill_1 FILLER_21_1068 ();
 sg13g2_decap_8 FILLER_21_1110 ();
 sg13g2_decap_4 FILLER_21_1117 ();
 sg13g2_fill_1 FILLER_21_1121 ();
 sg13g2_decap_8 FILLER_21_1128 ();
 sg13g2_decap_8 FILLER_21_1135 ();
 sg13g2_decap_4 FILLER_21_1142 ();
 sg13g2_fill_1 FILLER_21_1146 ();
 sg13g2_decap_4 FILLER_21_1184 ();
 sg13g2_fill_2 FILLER_21_1188 ();
 sg13g2_decap_8 FILLER_21_1200 ();
 sg13g2_decap_8 FILLER_21_1207 ();
 sg13g2_fill_2 FILLER_21_1214 ();
 sg13g2_fill_1 FILLER_21_1216 ();
 sg13g2_decap_8 FILLER_21_1236 ();
 sg13g2_decap_8 FILLER_21_1243 ();
 sg13g2_fill_2 FILLER_21_1250 ();
 sg13g2_decap_4 FILLER_21_1257 ();
 sg13g2_decap_8 FILLER_21_1267 ();
 sg13g2_fill_2 FILLER_21_1274 ();
 sg13g2_fill_2 FILLER_21_1280 ();
 sg13g2_fill_1 FILLER_21_1282 ();
 sg13g2_decap_4 FILLER_21_1300 ();
 sg13g2_fill_1 FILLER_21_1304 ();
 sg13g2_fill_2 FILLER_21_1308 ();
 sg13g2_decap_8 FILLER_21_1317 ();
 sg13g2_decap_4 FILLER_21_1324 ();
 sg13g2_fill_2 FILLER_21_1328 ();
 sg13g2_fill_1 FILLER_21_1335 ();
 sg13g2_decap_8 FILLER_21_1340 ();
 sg13g2_decap_4 FILLER_21_1347 ();
 sg13g2_fill_2 FILLER_21_1351 ();
 sg13g2_fill_2 FILLER_21_1377 ();
 sg13g2_fill_1 FILLER_21_1384 ();
 sg13g2_fill_2 FILLER_21_1390 ();
 sg13g2_fill_1 FILLER_21_1396 ();
 sg13g2_fill_1 FILLER_21_1405 ();
 sg13g2_fill_1 FILLER_21_1411 ();
 sg13g2_fill_2 FILLER_21_1416 ();
 sg13g2_decap_8 FILLER_21_1422 ();
 sg13g2_decap_4 FILLER_21_1429 ();
 sg13g2_fill_1 FILLER_21_1433 ();
 sg13g2_fill_1 FILLER_21_1446 ();
 sg13g2_decap_4 FILLER_21_1455 ();
 sg13g2_fill_2 FILLER_21_1485 ();
 sg13g2_fill_1 FILLER_21_1487 ();
 sg13g2_decap_8 FILLER_21_1523 ();
 sg13g2_fill_1 FILLER_21_1530 ();
 sg13g2_decap_4 FILLER_21_1541 ();
 sg13g2_fill_2 FILLER_21_1557 ();
 sg13g2_fill_1 FILLER_21_1559 ();
 sg13g2_decap_4 FILLER_21_1566 ();
 sg13g2_fill_2 FILLER_21_1596 ();
 sg13g2_fill_1 FILLER_21_1626 ();
 sg13g2_decap_8 FILLER_21_1636 ();
 sg13g2_decap_4 FILLER_21_1643 ();
 sg13g2_decap_4 FILLER_21_1650 ();
 sg13g2_fill_1 FILLER_21_1654 ();
 sg13g2_fill_2 FILLER_21_1664 ();
 sg13g2_fill_1 FILLER_21_1666 ();
 sg13g2_decap_8 FILLER_21_1677 ();
 sg13g2_decap_8 FILLER_21_1684 ();
 sg13g2_decap_8 FILLER_21_1691 ();
 sg13g2_decap_8 FILLER_21_1698 ();
 sg13g2_decap_4 FILLER_21_1705 ();
 sg13g2_fill_2 FILLER_21_1709 ();
 sg13g2_fill_2 FILLER_21_1721 ();
 sg13g2_fill_1 FILLER_21_1727 ();
 sg13g2_decap_8 FILLER_21_1732 ();
 sg13g2_decap_4 FILLER_21_1739 ();
 sg13g2_fill_1 FILLER_21_1743 ();
 sg13g2_decap_4 FILLER_21_1750 ();
 sg13g2_decap_8 FILLER_21_1760 ();
 sg13g2_decap_8 FILLER_21_1767 ();
 sg13g2_decap_8 FILLER_21_1774 ();
 sg13g2_decap_8 FILLER_21_1781 ();
 sg13g2_decap_4 FILLER_21_1788 ();
 sg13g2_fill_1 FILLER_21_1792 ();
 sg13g2_fill_2 FILLER_21_1798 ();
 sg13g2_decap_8 FILLER_21_1810 ();
 sg13g2_decap_8 FILLER_21_1817 ();
 sg13g2_fill_2 FILLER_21_1824 ();
 sg13g2_fill_1 FILLER_21_1826 ();
 sg13g2_fill_1 FILLER_21_1832 ();
 sg13g2_fill_1 FILLER_21_1859 ();
 sg13g2_fill_2 FILLER_21_1916 ();
 sg13g2_fill_1 FILLER_21_1918 ();
 sg13g2_fill_1 FILLER_21_1928 ();
 sg13g2_decap_4 FILLER_21_1938 ();
 sg13g2_fill_2 FILLER_21_1947 ();
 sg13g2_fill_1 FILLER_21_1949 ();
 sg13g2_decap_8 FILLER_21_1981 ();
 sg13g2_fill_2 FILLER_21_1988 ();
 sg13g2_fill_2 FILLER_21_1995 ();
 sg13g2_fill_1 FILLER_21_1997 ();
 sg13g2_fill_2 FILLER_21_2024 ();
 sg13g2_fill_1 FILLER_21_2026 ();
 sg13g2_fill_2 FILLER_21_2053 ();
 sg13g2_fill_2 FILLER_21_2081 ();
 sg13g2_fill_1 FILLER_21_2083 ();
 sg13g2_decap_8 FILLER_21_2096 ();
 sg13g2_decap_8 FILLER_21_2111 ();
 sg13g2_fill_2 FILLER_21_2118 ();
 sg13g2_decap_4 FILLER_21_2134 ();
 sg13g2_fill_2 FILLER_21_2151 ();
 sg13g2_fill_2 FILLER_21_2208 ();
 sg13g2_fill_1 FILLER_21_2230 ();
 sg13g2_fill_1 FILLER_21_2237 ();
 sg13g2_fill_1 FILLER_21_2264 ();
 sg13g2_fill_1 FILLER_21_2270 ();
 sg13g2_decap_8 FILLER_21_2281 ();
 sg13g2_decap_4 FILLER_21_2288 ();
 sg13g2_fill_1 FILLER_21_2297 ();
 sg13g2_decap_8 FILLER_21_2311 ();
 sg13g2_decap_4 FILLER_21_2318 ();
 sg13g2_decap_8 FILLER_21_2339 ();
 sg13g2_fill_2 FILLER_21_2346 ();
 sg13g2_fill_1 FILLER_21_2348 ();
 sg13g2_decap_8 FILLER_21_2378 ();
 sg13g2_fill_2 FILLER_21_2389 ();
 sg13g2_decap_8 FILLER_21_2404 ();
 sg13g2_decap_8 FILLER_21_2411 ();
 sg13g2_decap_8 FILLER_21_2418 ();
 sg13g2_decap_4 FILLER_21_2425 ();
 sg13g2_fill_1 FILLER_21_2429 ();
 sg13g2_decap_8 FILLER_21_2470 ();
 sg13g2_decap_8 FILLER_21_2477 ();
 sg13g2_decap_8 FILLER_21_2484 ();
 sg13g2_fill_2 FILLER_21_2491 ();
 sg13g2_fill_1 FILLER_21_2493 ();
 sg13g2_decap_8 FILLER_21_2532 ();
 sg13g2_decap_8 FILLER_21_2539 ();
 sg13g2_decap_8 FILLER_21_2546 ();
 sg13g2_decap_8 FILLER_21_2553 ();
 sg13g2_decap_8 FILLER_21_2560 ();
 sg13g2_decap_8 FILLER_21_2567 ();
 sg13g2_decap_8 FILLER_21_2574 ();
 sg13g2_decap_8 FILLER_21_2581 ();
 sg13g2_decap_8 FILLER_21_2588 ();
 sg13g2_decap_8 FILLER_21_2595 ();
 sg13g2_decap_8 FILLER_21_2602 ();
 sg13g2_decap_8 FILLER_21_2609 ();
 sg13g2_decap_8 FILLER_21_2616 ();
 sg13g2_decap_8 FILLER_21_2623 ();
 sg13g2_decap_8 FILLER_21_2630 ();
 sg13g2_decap_8 FILLER_21_2637 ();
 sg13g2_decap_8 FILLER_21_2644 ();
 sg13g2_decap_8 FILLER_21_2651 ();
 sg13g2_decap_8 FILLER_21_2658 ();
 sg13g2_decap_4 FILLER_21_2665 ();
 sg13g2_fill_1 FILLER_21_2669 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_4 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_78 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_114 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_129 ();
 sg13g2_decap_8 FILLER_22_136 ();
 sg13g2_decap_8 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_decap_4 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_272 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_4 FILLER_22_369 ();
 sg13g2_fill_2 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_4 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_1 FILLER_22_406 ();
 sg13g2_decap_4 FILLER_22_412 ();
 sg13g2_fill_2 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_433 ();
 sg13g2_decap_4 FILLER_22_441 ();
 sg13g2_fill_2 FILLER_22_451 ();
 sg13g2_fill_1 FILLER_22_453 ();
 sg13g2_decap_8 FILLER_22_491 ();
 sg13g2_decap_4 FILLER_22_498 ();
 sg13g2_fill_2 FILLER_22_502 ();
 sg13g2_decap_8 FILLER_22_509 ();
 sg13g2_decap_4 FILLER_22_516 ();
 sg13g2_fill_2 FILLER_22_529 ();
 sg13g2_decap_4 FILLER_22_561 ();
 sg13g2_fill_2 FILLER_22_599 ();
 sg13g2_fill_2 FILLER_22_633 ();
 sg13g2_fill_1 FILLER_22_635 ();
 sg13g2_decap_8 FILLER_22_649 ();
 sg13g2_fill_2 FILLER_22_656 ();
 sg13g2_fill_1 FILLER_22_663 ();
 sg13g2_fill_1 FILLER_22_744 ();
 sg13g2_fill_2 FILLER_22_754 ();
 sg13g2_fill_1 FILLER_22_756 ();
 sg13g2_fill_1 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_790 ();
 sg13g2_decap_8 FILLER_22_797 ();
 sg13g2_decap_4 FILLER_22_804 ();
 sg13g2_fill_1 FILLER_22_808 ();
 sg13g2_decap_8 FILLER_22_813 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_fill_2 FILLER_22_852 ();
 sg13g2_decap_8 FILLER_22_858 ();
 sg13g2_decap_4 FILLER_22_865 ();
 sg13g2_fill_2 FILLER_22_869 ();
 sg13g2_decap_8 FILLER_22_876 ();
 sg13g2_fill_1 FILLER_22_883 ();
 sg13g2_decap_8 FILLER_22_888 ();
 sg13g2_fill_2 FILLER_22_895 ();
 sg13g2_fill_2 FILLER_22_923 ();
 sg13g2_fill_2 FILLER_22_933 ();
 sg13g2_fill_1 FILLER_22_935 ();
 sg13g2_fill_2 FILLER_22_944 ();
 sg13g2_fill_1 FILLER_22_946 ();
 sg13g2_fill_2 FILLER_22_973 ();
 sg13g2_decap_4 FILLER_22_980 ();
 sg13g2_decap_4 FILLER_22_989 ();
 sg13g2_fill_1 FILLER_22_997 ();
 sg13g2_fill_2 FILLER_22_1032 ();
 sg13g2_fill_1 FILLER_22_1034 ();
 sg13g2_decap_4 FILLER_22_1067 ();
 sg13g2_fill_1 FILLER_22_1071 ();
 sg13g2_decap_8 FILLER_22_1084 ();
 sg13g2_fill_2 FILLER_22_1091 ();
 sg13g2_fill_2 FILLER_22_1101 ();
 sg13g2_fill_1 FILLER_22_1103 ();
 sg13g2_fill_1 FILLER_22_1112 ();
 sg13g2_fill_1 FILLER_22_1139 ();
 sg13g2_fill_1 FILLER_22_1148 ();
 sg13g2_fill_2 FILLER_22_1163 ();
 sg13g2_fill_1 FILLER_22_1183 ();
 sg13g2_fill_2 FILLER_22_1223 ();
 sg13g2_fill_1 FILLER_22_1228 ();
 sg13g2_decap_4 FILLER_22_1271 ();
 sg13g2_fill_1 FILLER_22_1275 ();
 sg13g2_fill_1 FILLER_22_1282 ();
 sg13g2_decap_8 FILLER_22_1347 ();
 sg13g2_decap_4 FILLER_22_1354 ();
 sg13g2_fill_2 FILLER_22_1370 ();
 sg13g2_fill_1 FILLER_22_1372 ();
 sg13g2_fill_1 FILLER_22_1377 ();
 sg13g2_fill_2 FILLER_22_1404 ();
 sg13g2_fill_1 FILLER_22_1406 ();
 sg13g2_decap_8 FILLER_22_1410 ();
 sg13g2_fill_2 FILLER_22_1421 ();
 sg13g2_decap_4 FILLER_22_1463 ();
 sg13g2_fill_2 FILLER_22_1467 ();
 sg13g2_decap_8 FILLER_22_1473 ();
 sg13g2_decap_8 FILLER_22_1480 ();
 sg13g2_fill_2 FILLER_22_1487 ();
 sg13g2_decap_8 FILLER_22_1494 ();
 sg13g2_fill_1 FILLER_22_1501 ();
 sg13g2_decap_8 FILLER_22_1512 ();
 sg13g2_decap_4 FILLER_22_1519 ();
 sg13g2_fill_1 FILLER_22_1523 ();
 sg13g2_fill_2 FILLER_22_1546 ();
 sg13g2_decap_4 FILLER_22_1580 ();
 sg13g2_fill_2 FILLER_22_1584 ();
 sg13g2_fill_2 FILLER_22_1595 ();
 sg13g2_fill_1 FILLER_22_1597 ();
 sg13g2_fill_1 FILLER_22_1607 ();
 sg13g2_decap_8 FILLER_22_1614 ();
 sg13g2_decap_8 FILLER_22_1621 ();
 sg13g2_decap_4 FILLER_22_1628 ();
 sg13g2_fill_1 FILLER_22_1632 ();
 sg13g2_decap_4 FILLER_22_1664 ();
 sg13g2_fill_1 FILLER_22_1668 ();
 sg13g2_decap_8 FILLER_22_1683 ();
 sg13g2_decap_8 FILLER_22_1694 ();
 sg13g2_decap_4 FILLER_22_1701 ();
 sg13g2_decap_8 FILLER_22_1734 ();
 sg13g2_fill_2 FILLER_22_1745 ();
 sg13g2_decap_8 FILLER_22_1773 ();
 sg13g2_fill_2 FILLER_22_1780 ();
 sg13g2_fill_1 FILLER_22_1788 ();
 sg13g2_fill_2 FILLER_22_1815 ();
 sg13g2_fill_1 FILLER_22_1817 ();
 sg13g2_fill_1 FILLER_22_1853 ();
 sg13g2_fill_2 FILLER_22_1858 ();
 sg13g2_decap_4 FILLER_22_1865 ();
 sg13g2_fill_1 FILLER_22_1873 ();
 sg13g2_fill_2 FILLER_22_1880 ();
 sg13g2_fill_2 FILLER_22_1887 ();
 sg13g2_decap_8 FILLER_22_1894 ();
 sg13g2_decap_8 FILLER_22_1901 ();
 sg13g2_decap_8 FILLER_22_1942 ();
 sg13g2_decap_4 FILLER_22_1949 ();
 sg13g2_fill_2 FILLER_22_1953 ();
 sg13g2_fill_1 FILLER_22_1981 ();
 sg13g2_fill_2 FILLER_22_2008 ();
 sg13g2_fill_1 FILLER_22_2010 ();
 sg13g2_fill_2 FILLER_22_2040 ();
 sg13g2_fill_2 FILLER_22_2046 ();
 sg13g2_fill_1 FILLER_22_2048 ();
 sg13g2_fill_2 FILLER_22_2054 ();
 sg13g2_decap_4 FILLER_22_2071 ();
 sg13g2_decap_8 FILLER_22_2096 ();
 sg13g2_decap_8 FILLER_22_2107 ();
 sg13g2_fill_2 FILLER_22_2148 ();
 sg13g2_fill_1 FILLER_22_2150 ();
 sg13g2_decap_4 FILLER_22_2155 ();
 sg13g2_fill_2 FILLER_22_2159 ();
 sg13g2_fill_1 FILLER_22_2192 ();
 sg13g2_fill_1 FILLER_22_2232 ();
 sg13g2_decap_8 FILLER_22_2270 ();
 sg13g2_decap_8 FILLER_22_2277 ();
 sg13g2_fill_2 FILLER_22_2284 ();
 sg13g2_fill_1 FILLER_22_2286 ();
 sg13g2_decap_8 FILLER_22_2300 ();
 sg13g2_decap_8 FILLER_22_2307 ();
 sg13g2_decap_8 FILLER_22_2314 ();
 sg13g2_decap_4 FILLER_22_2321 ();
 sg13g2_fill_2 FILLER_22_2333 ();
 sg13g2_fill_1 FILLER_22_2335 ();
 sg13g2_decap_4 FILLER_22_2353 ();
 sg13g2_fill_2 FILLER_22_2365 ();
 sg13g2_decap_8 FILLER_22_2398 ();
 sg13g2_decap_8 FILLER_22_2405 ();
 sg13g2_decap_8 FILLER_22_2412 ();
 sg13g2_decap_8 FILLER_22_2419 ();
 sg13g2_decap_4 FILLER_22_2456 ();
 sg13g2_decap_8 FILLER_22_2486 ();
 sg13g2_fill_2 FILLER_22_2493 ();
 sg13g2_decap_8 FILLER_22_2499 ();
 sg13g2_decap_4 FILLER_22_2506 ();
 sg13g2_fill_2 FILLER_22_2510 ();
 sg13g2_decap_4 FILLER_22_2516 ();
 sg13g2_decap_8 FILLER_22_2524 ();
 sg13g2_decap_8 FILLER_22_2531 ();
 sg13g2_decap_8 FILLER_22_2538 ();
 sg13g2_decap_8 FILLER_22_2545 ();
 sg13g2_decap_8 FILLER_22_2552 ();
 sg13g2_decap_8 FILLER_22_2559 ();
 sg13g2_decap_8 FILLER_22_2566 ();
 sg13g2_decap_8 FILLER_22_2573 ();
 sg13g2_decap_8 FILLER_22_2580 ();
 sg13g2_decap_8 FILLER_22_2587 ();
 sg13g2_decap_8 FILLER_22_2594 ();
 sg13g2_decap_8 FILLER_22_2601 ();
 sg13g2_decap_8 FILLER_22_2608 ();
 sg13g2_decap_8 FILLER_22_2615 ();
 sg13g2_decap_8 FILLER_22_2622 ();
 sg13g2_decap_8 FILLER_22_2629 ();
 sg13g2_decap_8 FILLER_22_2636 ();
 sg13g2_decap_8 FILLER_22_2643 ();
 sg13g2_decap_8 FILLER_22_2650 ();
 sg13g2_decap_8 FILLER_22_2657 ();
 sg13g2_decap_4 FILLER_22_2664 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_115 ();
 sg13g2_decap_4 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_134 ();
 sg13g2_fill_2 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_decap_8 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_fill_2 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_458 ();
 sg13g2_fill_1 FILLER_23_465 ();
 sg13g2_fill_2 FILLER_23_496 ();
 sg13g2_fill_1 FILLER_23_511 ();
 sg13g2_decap_4 FILLER_23_542 ();
 sg13g2_decap_8 FILLER_23_577 ();
 sg13g2_fill_1 FILLER_23_600 ();
 sg13g2_fill_2 FILLER_23_614 ();
 sg13g2_fill_1 FILLER_23_621 ();
 sg13g2_fill_2 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_694 ();
 sg13g2_fill_2 FILLER_23_701 ();
 sg13g2_fill_1 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_fill_1 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_745 ();
 sg13g2_fill_1 FILLER_23_752 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_fill_1 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_786 ();
 sg13g2_decap_8 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_800 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_831 ();
 sg13g2_fill_2 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_870 ();
 sg13g2_decap_8 FILLER_23_877 ();
 sg13g2_decap_8 FILLER_23_884 ();
 sg13g2_fill_2 FILLER_23_891 ();
 sg13g2_fill_2 FILLER_23_906 ();
 sg13g2_fill_1 FILLER_23_908 ();
 sg13g2_fill_2 FILLER_23_921 ();
 sg13g2_fill_1 FILLER_23_961 ();
 sg13g2_fill_2 FILLER_23_988 ();
 sg13g2_decap_8 FILLER_23_1002 ();
 sg13g2_decap_8 FILLER_23_1009 ();
 sg13g2_decap_8 FILLER_23_1016 ();
 sg13g2_fill_2 FILLER_23_1023 ();
 sg13g2_fill_2 FILLER_23_1030 ();
 sg13g2_fill_1 FILLER_23_1074 ();
 sg13g2_decap_4 FILLER_23_1106 ();
 sg13g2_fill_1 FILLER_23_1110 ();
 sg13g2_fill_1 FILLER_23_1115 ();
 sg13g2_decap_4 FILLER_23_1167 ();
 sg13g2_fill_1 FILLER_23_1179 ();
 sg13g2_decap_4 FILLER_23_1196 ();
 sg13g2_fill_2 FILLER_23_1250 ();
 sg13g2_fill_1 FILLER_23_1292 ();
 sg13g2_fill_2 FILLER_23_1311 ();
 sg13g2_fill_2 FILLER_23_1316 ();
 sg13g2_decap_4 FILLER_23_1344 ();
 sg13g2_fill_2 FILLER_23_1348 ();
 sg13g2_fill_2 FILLER_23_1361 ();
 sg13g2_fill_1 FILLER_23_1367 ();
 sg13g2_fill_1 FILLER_23_1377 ();
 sg13g2_fill_1 FILLER_23_1405 ();
 sg13g2_fill_1 FILLER_23_1411 ();
 sg13g2_decap_8 FILLER_23_1421 ();
 sg13g2_decap_8 FILLER_23_1428 ();
 sg13g2_decap_8 FILLER_23_1435 ();
 sg13g2_fill_2 FILLER_23_1442 ();
 sg13g2_fill_1 FILLER_23_1444 ();
 sg13g2_decap_8 FILLER_23_1476 ();
 sg13g2_decap_4 FILLER_23_1483 ();
 sg13g2_fill_1 FILLER_23_1487 ();
 sg13g2_decap_8 FILLER_23_1497 ();
 sg13g2_decap_8 FILLER_23_1560 ();
 sg13g2_decap_8 FILLER_23_1567 ();
 sg13g2_decap_8 FILLER_23_1574 ();
 sg13g2_fill_2 FILLER_23_1589 ();
 sg13g2_decap_4 FILLER_23_1617 ();
 sg13g2_decap_8 FILLER_23_1624 ();
 sg13g2_decap_8 FILLER_23_1631 ();
 sg13g2_decap_4 FILLER_23_1638 ();
 sg13g2_fill_1 FILLER_23_1642 ();
 sg13g2_fill_2 FILLER_23_1669 ();
 sg13g2_fill_1 FILLER_23_1697 ();
 sg13g2_fill_1 FILLER_23_1710 ();
 sg13g2_decap_4 FILLER_23_1737 ();
 sg13g2_fill_1 FILLER_23_1778 ();
 sg13g2_decap_8 FILLER_23_1819 ();
 sg13g2_fill_2 FILLER_23_1826 ();
 sg13g2_fill_1 FILLER_23_1828 ();
 sg13g2_decap_8 FILLER_23_1833 ();
 sg13g2_decap_8 FILLER_23_1840 ();
 sg13g2_decap_8 FILLER_23_1847 ();
 sg13g2_decap_8 FILLER_23_1939 ();
 sg13g2_decap_8 FILLER_23_1946 ();
 sg13g2_fill_1 FILLER_23_1953 ();
 sg13g2_decap_8 FILLER_23_1958 ();
 sg13g2_decap_8 FILLER_23_1965 ();
 sg13g2_decap_8 FILLER_23_1972 ();
 sg13g2_fill_2 FILLER_23_1979 ();
 sg13g2_fill_2 FILLER_23_1990 ();
 sg13g2_fill_1 FILLER_23_1992 ();
 sg13g2_decap_4 FILLER_23_2082 ();
 sg13g2_fill_1 FILLER_23_2086 ();
 sg13g2_decap_8 FILLER_23_2116 ();
 sg13g2_fill_2 FILLER_23_2123 ();
 sg13g2_fill_1 FILLER_23_2125 ();
 sg13g2_fill_1 FILLER_23_2130 ();
 sg13g2_decap_8 FILLER_23_2139 ();
 sg13g2_decap_8 FILLER_23_2146 ();
 sg13g2_fill_1 FILLER_23_2153 ();
 sg13g2_decap_8 FILLER_23_2167 ();
 sg13g2_decap_8 FILLER_23_2174 ();
 sg13g2_decap_8 FILLER_23_2181 ();
 sg13g2_fill_2 FILLER_23_2188 ();
 sg13g2_fill_2 FILLER_23_2196 ();
 sg13g2_fill_2 FILLER_23_2263 ();
 sg13g2_decap_4 FILLER_23_2300 ();
 sg13g2_fill_1 FILLER_23_2304 ();
 sg13g2_decap_8 FILLER_23_2310 ();
 sg13g2_decap_4 FILLER_23_2317 ();
 sg13g2_fill_2 FILLER_23_2321 ();
 sg13g2_decap_8 FILLER_23_2364 ();
 sg13g2_fill_1 FILLER_23_2371 ();
 sg13g2_decap_8 FILLER_23_2381 ();
 sg13g2_decap_4 FILLER_23_2388 ();
 sg13g2_fill_1 FILLER_23_2392 ();
 sg13g2_decap_8 FILLER_23_2405 ();
 sg13g2_decap_8 FILLER_23_2412 ();
 sg13g2_fill_2 FILLER_23_2419 ();
 sg13g2_fill_1 FILLER_23_2474 ();
 sg13g2_decap_8 FILLER_23_2501 ();
 sg13g2_decap_8 FILLER_23_2508 ();
 sg13g2_decap_8 FILLER_23_2515 ();
 sg13g2_decap_8 FILLER_23_2522 ();
 sg13g2_decap_8 FILLER_23_2529 ();
 sg13g2_decap_8 FILLER_23_2536 ();
 sg13g2_decap_8 FILLER_23_2543 ();
 sg13g2_decap_8 FILLER_23_2550 ();
 sg13g2_decap_8 FILLER_23_2557 ();
 sg13g2_decap_8 FILLER_23_2564 ();
 sg13g2_decap_8 FILLER_23_2571 ();
 sg13g2_decap_8 FILLER_23_2578 ();
 sg13g2_decap_8 FILLER_23_2585 ();
 sg13g2_decap_8 FILLER_23_2592 ();
 sg13g2_decap_8 FILLER_23_2599 ();
 sg13g2_decap_8 FILLER_23_2606 ();
 sg13g2_decap_8 FILLER_23_2613 ();
 sg13g2_decap_8 FILLER_23_2620 ();
 sg13g2_decap_8 FILLER_23_2627 ();
 sg13g2_decap_8 FILLER_23_2634 ();
 sg13g2_decap_8 FILLER_23_2641 ();
 sg13g2_decap_8 FILLER_23_2648 ();
 sg13g2_decap_8 FILLER_23_2655 ();
 sg13g2_decap_8 FILLER_23_2662 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_117 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_fill_2 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_decap_4 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_8 FILLER_24_405 ();
 sg13g2_fill_2 FILLER_24_412 ();
 sg13g2_decap_4 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_428 ();
 sg13g2_fill_2 FILLER_24_436 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_444 ();
 sg13g2_decap_4 FILLER_24_451 ();
 sg13g2_fill_1 FILLER_24_455 ();
 sg13g2_fill_2 FILLER_24_470 ();
 sg13g2_decap_4 FILLER_24_498 ();
 sg13g2_fill_2 FILLER_24_502 ();
 sg13g2_decap_4 FILLER_24_540 ();
 sg13g2_fill_1 FILLER_24_544 ();
 sg13g2_decap_8 FILLER_24_554 ();
 sg13g2_decap_8 FILLER_24_561 ();
 sg13g2_decap_8 FILLER_24_568 ();
 sg13g2_decap_8 FILLER_24_575 ();
 sg13g2_fill_1 FILLER_24_582 ();
 sg13g2_fill_1 FILLER_24_602 ();
 sg13g2_fill_2 FILLER_24_612 ();
 sg13g2_decap_4 FILLER_24_618 ();
 sg13g2_decap_8 FILLER_24_631 ();
 sg13g2_fill_1 FILLER_24_638 ();
 sg13g2_decap_4 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_652 ();
 sg13g2_decap_8 FILLER_24_659 ();
 sg13g2_fill_1 FILLER_24_678 ();
 sg13g2_decap_8 FILLER_24_688 ();
 sg13g2_fill_2 FILLER_24_695 ();
 sg13g2_fill_1 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_724 ();
 sg13g2_decap_8 FILLER_24_731 ();
 sg13g2_decap_4 FILLER_24_738 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_fill_2 FILLER_24_753 ();
 sg13g2_decap_4 FILLER_24_795 ();
 sg13g2_fill_1 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_fill_2 FILLER_24_817 ();
 sg13g2_fill_1 FILLER_24_819 ();
 sg13g2_fill_1 FILLER_24_850 ();
 sg13g2_decap_8 FILLER_24_859 ();
 sg13g2_decap_4 FILLER_24_866 ();
 sg13g2_fill_1 FILLER_24_870 ();
 sg13g2_fill_1 FILLER_24_914 ();
 sg13g2_fill_2 FILLER_24_941 ();
 sg13g2_fill_1 FILLER_24_943 ();
 sg13g2_fill_2 FILLER_24_952 ();
 sg13g2_fill_1 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1009 ();
 sg13g2_decap_4 FILLER_24_1016 ();
 sg13g2_fill_2 FILLER_24_1020 ();
 sg13g2_decap_4 FILLER_24_1085 ();
 sg13g2_decap_8 FILLER_24_1098 ();
 sg13g2_decap_4 FILLER_24_1105 ();
 sg13g2_fill_2 FILLER_24_1109 ();
 sg13g2_fill_1 FILLER_24_1116 ();
 sg13g2_decap_4 FILLER_24_1136 ();
 sg13g2_fill_2 FILLER_24_1140 ();
 sg13g2_fill_1 FILLER_24_1146 ();
 sg13g2_decap_4 FILLER_24_1156 ();
 sg13g2_fill_1 FILLER_24_1160 ();
 sg13g2_decap_4 FILLER_24_1166 ();
 sg13g2_fill_2 FILLER_24_1174 ();
 sg13g2_fill_1 FILLER_24_1176 ();
 sg13g2_fill_2 FILLER_24_1200 ();
 sg13g2_fill_2 FILLER_24_1210 ();
 sg13g2_fill_1 FILLER_24_1242 ();
 sg13g2_decap_8 FILLER_24_1269 ();
 sg13g2_decap_8 FILLER_24_1281 ();
 sg13g2_decap_4 FILLER_24_1288 ();
 sg13g2_fill_2 FILLER_24_1292 ();
 sg13g2_fill_1 FILLER_24_1304 ();
 sg13g2_fill_2 FILLER_24_1318 ();
 sg13g2_fill_1 FILLER_24_1320 ();
 sg13g2_decap_4 FILLER_24_1325 ();
 sg13g2_fill_2 FILLER_24_1350 ();
 sg13g2_decap_4 FILLER_24_1386 ();
 sg13g2_fill_2 FILLER_24_1390 ();
 sg13g2_decap_4 FILLER_24_1407 ();
 sg13g2_decap_8 FILLER_24_1443 ();
 sg13g2_decap_4 FILLER_24_1450 ();
 sg13g2_fill_1 FILLER_24_1454 ();
 sg13g2_decap_8 FILLER_24_1468 ();
 sg13g2_fill_1 FILLER_24_1475 ();
 sg13g2_fill_2 FILLER_24_1485 ();
 sg13g2_decap_8 FILLER_24_1513 ();
 sg13g2_decap_4 FILLER_24_1520 ();
 sg13g2_fill_2 FILLER_24_1524 ();
 sg13g2_decap_8 FILLER_24_1535 ();
 sg13g2_decap_8 FILLER_24_1542 ();
 sg13g2_decap_8 FILLER_24_1549 ();
 sg13g2_decap_8 FILLER_24_1556 ();
 sg13g2_decap_8 FILLER_24_1563 ();
 sg13g2_decap_4 FILLER_24_1575 ();
 sg13g2_fill_1 FILLER_24_1627 ();
 sg13g2_decap_8 FILLER_24_1636 ();
 sg13g2_decap_8 FILLER_24_1648 ();
 sg13g2_decap_8 FILLER_24_1655 ();
 sg13g2_fill_1 FILLER_24_1706 ();
 sg13g2_decap_4 FILLER_24_1746 ();
 sg13g2_fill_1 FILLER_24_1750 ();
 sg13g2_fill_1 FILLER_24_1762 ();
 sg13g2_fill_2 FILLER_24_1772 ();
 sg13g2_fill_1 FILLER_24_1774 ();
 sg13g2_decap_8 FILLER_24_1779 ();
 sg13g2_decap_4 FILLER_24_1786 ();
 sg13g2_fill_2 FILLER_24_1790 ();
 sg13g2_decap_4 FILLER_24_1797 ();
 sg13g2_fill_2 FILLER_24_1801 ();
 sg13g2_decap_8 FILLER_24_1807 ();
 sg13g2_decap_8 FILLER_24_1814 ();
 sg13g2_decap_8 FILLER_24_1821 ();
 sg13g2_decap_8 FILLER_24_1828 ();
 sg13g2_decap_8 FILLER_24_1835 ();
 sg13g2_decap_8 FILLER_24_1842 ();
 sg13g2_decap_8 FILLER_24_1849 ();
 sg13g2_decap_4 FILLER_24_1856 ();
 sg13g2_fill_2 FILLER_24_1860 ();
 sg13g2_decap_8 FILLER_24_1866 ();
 sg13g2_fill_2 FILLER_24_1890 ();
 sg13g2_fill_1 FILLER_24_1892 ();
 sg13g2_decap_8 FILLER_24_1897 ();
 sg13g2_fill_2 FILLER_24_1904 ();
 sg13g2_fill_1 FILLER_24_1906 ();
 sg13g2_decap_8 FILLER_24_1933 ();
 sg13g2_decap_8 FILLER_24_1940 ();
 sg13g2_fill_2 FILLER_24_1947 ();
 sg13g2_fill_1 FILLER_24_1949 ();
 sg13g2_fill_2 FILLER_24_1954 ();
 sg13g2_fill_1 FILLER_24_1956 ();
 sg13g2_decap_8 FILLER_24_1973 ();
 sg13g2_fill_1 FILLER_24_1980 ();
 sg13g2_fill_1 FILLER_24_1999 ();
 sg13g2_fill_1 FILLER_24_2006 ();
 sg13g2_fill_2 FILLER_24_2016 ();
 sg13g2_fill_2 FILLER_24_2022 ();
 sg13g2_fill_1 FILLER_24_2028 ();
 sg13g2_decap_4 FILLER_24_2034 ();
 sg13g2_fill_2 FILLER_24_2038 ();
 sg13g2_fill_2 FILLER_24_2045 ();
 sg13g2_fill_1 FILLER_24_2047 ();
 sg13g2_fill_2 FILLER_24_2057 ();
 sg13g2_fill_1 FILLER_24_2059 ();
 sg13g2_decap_4 FILLER_24_2069 ();
 sg13g2_decap_8 FILLER_24_2103 ();
 sg13g2_decap_8 FILLER_24_2110 ();
 sg13g2_decap_8 FILLER_24_2117 ();
 sg13g2_fill_2 FILLER_24_2124 ();
 sg13g2_fill_1 FILLER_24_2136 ();
 sg13g2_fill_2 FILLER_24_2141 ();
 sg13g2_fill_1 FILLER_24_2147 ();
 sg13g2_decap_8 FILLER_24_2153 ();
 sg13g2_decap_4 FILLER_24_2160 ();
 sg13g2_fill_2 FILLER_24_2164 ();
 sg13g2_fill_1 FILLER_24_2171 ();
 sg13g2_fill_1 FILLER_24_2203 ();
 sg13g2_fill_2 FILLER_24_2231 ();
 sg13g2_decap_8 FILLER_24_2257 ();
 sg13g2_decap_8 FILLER_24_2264 ();
 sg13g2_decap_8 FILLER_24_2271 ();
 sg13g2_fill_1 FILLER_24_2278 ();
 sg13g2_fill_2 FILLER_24_2340 ();
 sg13g2_fill_1 FILLER_24_2348 ();
 sg13g2_fill_2 FILLER_24_2353 ();
 sg13g2_fill_1 FILLER_24_2355 ();
 sg13g2_fill_2 FILLER_24_2362 ();
 sg13g2_fill_2 FILLER_24_2372 ();
 sg13g2_decap_8 FILLER_24_2426 ();
 sg13g2_decap_4 FILLER_24_2433 ();
 sg13g2_fill_1 FILLER_24_2437 ();
 sg13g2_fill_2 FILLER_24_2442 ();
 sg13g2_fill_1 FILLER_24_2444 ();
 sg13g2_fill_2 FILLER_24_2463 ();
 sg13g2_fill_1 FILLER_24_2487 ();
 sg13g2_decap_8 FILLER_24_2492 ();
 sg13g2_decap_8 FILLER_24_2499 ();
 sg13g2_decap_8 FILLER_24_2506 ();
 sg13g2_decap_4 FILLER_24_2513 ();
 sg13g2_fill_2 FILLER_24_2517 ();
 sg13g2_decap_8 FILLER_24_2523 ();
 sg13g2_decap_8 FILLER_24_2530 ();
 sg13g2_decap_8 FILLER_24_2537 ();
 sg13g2_decap_8 FILLER_24_2544 ();
 sg13g2_decap_8 FILLER_24_2551 ();
 sg13g2_decap_8 FILLER_24_2558 ();
 sg13g2_decap_8 FILLER_24_2565 ();
 sg13g2_decap_8 FILLER_24_2572 ();
 sg13g2_decap_8 FILLER_24_2579 ();
 sg13g2_decap_8 FILLER_24_2586 ();
 sg13g2_decap_8 FILLER_24_2593 ();
 sg13g2_decap_8 FILLER_24_2600 ();
 sg13g2_decap_8 FILLER_24_2607 ();
 sg13g2_decap_8 FILLER_24_2614 ();
 sg13g2_decap_8 FILLER_24_2621 ();
 sg13g2_decap_8 FILLER_24_2628 ();
 sg13g2_decap_8 FILLER_24_2635 ();
 sg13g2_decap_8 FILLER_24_2642 ();
 sg13g2_decap_8 FILLER_24_2649 ();
 sg13g2_decap_8 FILLER_24_2656 ();
 sg13g2_decap_8 FILLER_24_2663 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_61 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_decap_4 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_decap_4 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_4 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_25_447 ();
 sg13g2_decap_4 FILLER_25_454 ();
 sg13g2_fill_2 FILLER_25_458 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_4 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_fill_1 FILLER_25_553 ();
 sg13g2_fill_1 FILLER_25_569 ();
 sg13g2_fill_1 FILLER_25_606 ();
 sg13g2_fill_1 FILLER_25_620 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_fill_1 FILLER_25_729 ();
 sg13g2_decap_4 FILLER_25_756 ();
 sg13g2_fill_1 FILLER_25_772 ();
 sg13g2_fill_1 FILLER_25_799 ();
 sg13g2_fill_1 FILLER_25_831 ();
 sg13g2_fill_1 FILLER_25_836 ();
 sg13g2_decap_8 FILLER_25_872 ();
 sg13g2_decap_8 FILLER_25_879 ();
 sg13g2_decap_8 FILLER_25_886 ();
 sg13g2_decap_8 FILLER_25_893 ();
 sg13g2_decap_4 FILLER_25_900 ();
 sg13g2_fill_1 FILLER_25_904 ();
 sg13g2_decap_4 FILLER_25_911 ();
 sg13g2_fill_1 FILLER_25_920 ();
 sg13g2_fill_1 FILLER_25_925 ();
 sg13g2_fill_1 FILLER_25_932 ();
 sg13g2_decap_8 FILLER_25_938 ();
 sg13g2_fill_2 FILLER_25_945 ();
 sg13g2_fill_1 FILLER_25_947 ();
 sg13g2_fill_2 FILLER_25_961 ();
 sg13g2_fill_2 FILLER_25_972 ();
 sg13g2_fill_2 FILLER_25_977 ();
 sg13g2_fill_1 FILLER_25_979 ();
 sg13g2_fill_2 FILLER_25_985 ();
 sg13g2_fill_1 FILLER_25_987 ();
 sg13g2_decap_4 FILLER_25_996 ();
 sg13g2_fill_1 FILLER_25_1000 ();
 sg13g2_decap_4 FILLER_25_1007 ();
 sg13g2_fill_1 FILLER_25_1011 ();
 sg13g2_decap_4 FILLER_25_1018 ();
 sg13g2_fill_1 FILLER_25_1022 ();
 sg13g2_decap_8 FILLER_25_1027 ();
 sg13g2_fill_1 FILLER_25_1034 ();
 sg13g2_fill_2 FILLER_25_1045 ();
 sg13g2_fill_1 FILLER_25_1056 ();
 sg13g2_fill_1 FILLER_25_1083 ();
 sg13g2_fill_1 FILLER_25_1110 ();
 sg13g2_fill_2 FILLER_25_1121 ();
 sg13g2_fill_2 FILLER_25_1129 ();
 sg13g2_fill_1 FILLER_25_1137 ();
 sg13g2_fill_1 FILLER_25_1194 ();
 sg13g2_fill_1 FILLER_25_1204 ();
 sg13g2_fill_2 FILLER_25_1231 ();
 sg13g2_decap_4 FILLER_25_1253 ();
 sg13g2_decap_4 FILLER_25_1263 ();
 sg13g2_fill_2 FILLER_25_1267 ();
 sg13g2_decap_8 FILLER_25_1274 ();
 sg13g2_decap_8 FILLER_25_1281 ();
 sg13g2_decap_8 FILLER_25_1288 ();
 sg13g2_fill_1 FILLER_25_1295 ();
 sg13g2_fill_1 FILLER_25_1304 ();
 sg13g2_fill_1 FILLER_25_1337 ();
 sg13g2_fill_2 FILLER_25_1343 ();
 sg13g2_fill_1 FILLER_25_1345 ();
 sg13g2_fill_2 FILLER_25_1359 ();
 sg13g2_fill_1 FILLER_25_1387 ();
 sg13g2_decap_4 FILLER_25_1393 ();
 sg13g2_fill_2 FILLER_25_1444 ();
 sg13g2_fill_2 FILLER_25_1475 ();
 sg13g2_fill_1 FILLER_25_1503 ();
 sg13g2_decap_8 FILLER_25_1514 ();
 sg13g2_decap_8 FILLER_25_1521 ();
 sg13g2_decap_8 FILLER_25_1528 ();
 sg13g2_decap_8 FILLER_25_1535 ();
 sg13g2_decap_8 FILLER_25_1542 ();
 sg13g2_decap_8 FILLER_25_1549 ();
 sg13g2_decap_8 FILLER_25_1556 ();
 sg13g2_decap_8 FILLER_25_1563 ();
 sg13g2_decap_8 FILLER_25_1570 ();
 sg13g2_decap_8 FILLER_25_1577 ();
 sg13g2_fill_2 FILLER_25_1584 ();
 sg13g2_fill_2 FILLER_25_1613 ();
 sg13g2_fill_1 FILLER_25_1644 ();
 sg13g2_fill_1 FILLER_25_1698 ();
 sg13g2_fill_2 FILLER_25_1705 ();
 sg13g2_fill_2 FILLER_25_1712 ();
 sg13g2_fill_2 FILLER_25_1723 ();
 sg13g2_fill_1 FILLER_25_1729 ();
 sg13g2_decap_8 FILLER_25_1736 ();
 sg13g2_decap_8 FILLER_25_1743 ();
 sg13g2_decap_8 FILLER_25_1750 ();
 sg13g2_decap_8 FILLER_25_1783 ();
 sg13g2_decap_4 FILLER_25_1790 ();
 sg13g2_decap_8 FILLER_25_1798 ();
 sg13g2_decap_8 FILLER_25_1805 ();
 sg13g2_decap_4 FILLER_25_1812 ();
 sg13g2_fill_2 FILLER_25_1816 ();
 sg13g2_decap_4 FILLER_25_1874 ();
 sg13g2_fill_2 FILLER_25_1878 ();
 sg13g2_fill_2 FILLER_25_1911 ();
 sg13g2_fill_1 FILLER_25_1913 ();
 sg13g2_fill_1 FILLER_25_1920 ();
 sg13g2_decap_8 FILLER_25_1925 ();
 sg13g2_decap_8 FILLER_25_1932 ();
 sg13g2_decap_4 FILLER_25_1939 ();
 sg13g2_fill_1 FILLER_25_1943 ();
 sg13g2_decap_8 FILLER_25_1980 ();
 sg13g2_decap_4 FILLER_25_1987 ();
 sg13g2_fill_2 FILLER_25_1991 ();
 sg13g2_fill_2 FILLER_25_2012 ();
 sg13g2_decap_8 FILLER_25_2018 ();
 sg13g2_decap_4 FILLER_25_2025 ();
 sg13g2_fill_1 FILLER_25_2029 ();
 sg13g2_fill_2 FILLER_25_2066 ();
 sg13g2_decap_8 FILLER_25_2078 ();
 sg13g2_decap_8 FILLER_25_2111 ();
 sg13g2_decap_8 FILLER_25_2118 ();
 sg13g2_fill_1 FILLER_25_2125 ();
 sg13g2_fill_2 FILLER_25_2130 ();
 sg13g2_decap_8 FILLER_25_2193 ();
 sg13g2_decap_4 FILLER_25_2200 ();
 sg13g2_fill_1 FILLER_25_2204 ();
 sg13g2_fill_1 FILLER_25_2223 ();
 sg13g2_fill_2 FILLER_25_2230 ();
 sg13g2_fill_1 FILLER_25_2275 ();
 sg13g2_decap_4 FILLER_25_2302 ();
 sg13g2_fill_1 FILLER_25_2306 ();
 sg13g2_fill_2 FILLER_25_2385 ();
 sg13g2_fill_1 FILLER_25_2387 ();
 sg13g2_decap_8 FILLER_25_2423 ();
 sg13g2_decap_4 FILLER_25_2430 ();
 sg13g2_fill_2 FILLER_25_2434 ();
 sg13g2_fill_2 FILLER_25_2471 ();
 sg13g2_fill_1 FILLER_25_2473 ();
 sg13g2_decap_8 FILLER_25_2479 ();
 sg13g2_fill_1 FILLER_25_2486 ();
 sg13g2_decap_8 FILLER_25_2497 ();
 sg13g2_fill_1 FILLER_25_2504 ();
 sg13g2_decap_8 FILLER_25_2543 ();
 sg13g2_decap_8 FILLER_25_2550 ();
 sg13g2_decap_8 FILLER_25_2557 ();
 sg13g2_decap_8 FILLER_25_2564 ();
 sg13g2_decap_8 FILLER_25_2571 ();
 sg13g2_decap_8 FILLER_25_2578 ();
 sg13g2_decap_8 FILLER_25_2585 ();
 sg13g2_decap_8 FILLER_25_2592 ();
 sg13g2_decap_8 FILLER_25_2599 ();
 sg13g2_decap_8 FILLER_25_2606 ();
 sg13g2_decap_8 FILLER_25_2613 ();
 sg13g2_decap_8 FILLER_25_2620 ();
 sg13g2_decap_8 FILLER_25_2627 ();
 sg13g2_decap_8 FILLER_25_2634 ();
 sg13g2_decap_8 FILLER_25_2641 ();
 sg13g2_decap_8 FILLER_25_2648 ();
 sg13g2_decap_8 FILLER_25_2655 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_fill_1 FILLER_25_2669 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_15 ();
 sg13g2_decap_8 FILLER_26_22 ();
 sg13g2_fill_2 FILLER_26_29 ();
 sg13g2_fill_1 FILLER_26_31 ();
 sg13g2_fill_2 FILLER_26_36 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_decap_4 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_decap_4 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_237 ();
 sg13g2_fill_2 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_4 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_4 FILLER_26_382 ();
 sg13g2_fill_2 FILLER_26_386 ();
 sg13g2_decap_4 FILLER_26_396 ();
 sg13g2_fill_1 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_4 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_451 ();
 sg13g2_decap_8 FILLER_26_458 ();
 sg13g2_fill_1 FILLER_26_465 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_4 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_516 ();
 sg13g2_decap_8 FILLER_26_523 ();
 sg13g2_decap_8 FILLER_26_530 ();
 sg13g2_fill_1 FILLER_26_537 ();
 sg13g2_decap_8 FILLER_26_543 ();
 sg13g2_fill_1 FILLER_26_565 ();
 sg13g2_fill_2 FILLER_26_601 ();
 sg13g2_fill_1 FILLER_26_617 ();
 sg13g2_decap_8 FILLER_26_622 ();
 sg13g2_fill_2 FILLER_26_629 ();
 sg13g2_fill_1 FILLER_26_631 ();
 sg13g2_decap_8 FILLER_26_653 ();
 sg13g2_fill_2 FILLER_26_660 ();
 sg13g2_decap_8 FILLER_26_667 ();
 sg13g2_fill_2 FILLER_26_674 ();
 sg13g2_fill_1 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_697 ();
 sg13g2_fill_1 FILLER_26_716 ();
 sg13g2_fill_1 FILLER_26_726 ();
 sg13g2_fill_1 FILLER_26_759 ();
 sg13g2_decap_4 FILLER_26_786 ();
 sg13g2_decap_4 FILLER_26_796 ();
 sg13g2_fill_1 FILLER_26_800 ();
 sg13g2_decap_4 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_867 ();
 sg13g2_decap_8 FILLER_26_874 ();
 sg13g2_decap_8 FILLER_26_881 ();
 sg13g2_fill_2 FILLER_26_888 ();
 sg13g2_fill_1 FILLER_26_907 ();
 sg13g2_fill_2 FILLER_26_912 ();
 sg13g2_decap_8 FILLER_26_944 ();
 sg13g2_decap_4 FILLER_26_951 ();
 sg13g2_fill_1 FILLER_26_955 ();
 sg13g2_fill_2 FILLER_26_972 ();
 sg13g2_decap_4 FILLER_26_996 ();
 sg13g2_fill_1 FILLER_26_1000 ();
 sg13g2_fill_1 FILLER_26_1022 ();
 sg13g2_fill_2 FILLER_26_1055 ();
 sg13g2_fill_2 FILLER_26_1065 ();
 sg13g2_fill_2 FILLER_26_1091 ();
 sg13g2_fill_1 FILLER_26_1093 ();
 sg13g2_fill_2 FILLER_26_1120 ();
 sg13g2_decap_8 FILLER_26_1149 ();
 sg13g2_fill_2 FILLER_26_1156 ();
 sg13g2_fill_1 FILLER_26_1158 ();
 sg13g2_fill_2 FILLER_26_1163 ();
 sg13g2_decap_8 FILLER_26_1170 ();
 sg13g2_fill_1 FILLER_26_1177 ();
 sg13g2_decap_8 FILLER_26_1191 ();
 sg13g2_fill_1 FILLER_26_1198 ();
 sg13g2_decap_4 FILLER_26_1213 ();
 sg13g2_fill_1 FILLER_26_1217 ();
 sg13g2_decap_8 FILLER_26_1244 ();
 sg13g2_decap_8 FILLER_26_1251 ();
 sg13g2_fill_1 FILLER_26_1258 ();
 sg13g2_decap_8 FILLER_26_1316 ();
 sg13g2_decap_8 FILLER_26_1323 ();
 sg13g2_decap_8 FILLER_26_1335 ();
 sg13g2_fill_2 FILLER_26_1373 ();
 sg13g2_fill_1 FILLER_26_1375 ();
 sg13g2_decap_8 FILLER_26_1394 ();
 sg13g2_decap_8 FILLER_26_1401 ();
 sg13g2_decap_8 FILLER_26_1408 ();
 sg13g2_decap_8 FILLER_26_1425 ();
 sg13g2_decap_4 FILLER_26_1432 ();
 sg13g2_fill_2 FILLER_26_1436 ();
 sg13g2_fill_1 FILLER_26_1442 ();
 sg13g2_decap_4 FILLER_26_1451 ();
 sg13g2_decap_4 FILLER_26_1459 ();
 sg13g2_fill_1 FILLER_26_1463 ();
 sg13g2_fill_1 FILLER_26_1495 ();
 sg13g2_decap_8 FILLER_26_1522 ();
 sg13g2_decap_8 FILLER_26_1529 ();
 sg13g2_decap_8 FILLER_26_1536 ();
 sg13g2_decap_8 FILLER_26_1543 ();
 sg13g2_decap_8 FILLER_26_1550 ();
 sg13g2_decap_8 FILLER_26_1557 ();
 sg13g2_decap_4 FILLER_26_1564 ();
 sg13g2_fill_1 FILLER_26_1603 ();
 sg13g2_fill_1 FILLER_26_1628 ();
 sg13g2_fill_1 FILLER_26_1638 ();
 sg13g2_decap_4 FILLER_26_1669 ();
 sg13g2_fill_1 FILLER_26_1678 ();
 sg13g2_decap_8 FILLER_26_1704 ();
 sg13g2_fill_2 FILLER_26_1711 ();
 sg13g2_decap_8 FILLER_26_1717 ();
 sg13g2_decap_8 FILLER_26_1724 ();
 sg13g2_decap_4 FILLER_26_1731 ();
 sg13g2_fill_2 FILLER_26_1735 ();
 sg13g2_fill_2 FILLER_26_1742 ();
 sg13g2_fill_1 FILLER_26_1744 ();
 sg13g2_decap_8 FILLER_26_1753 ();
 sg13g2_fill_2 FILLER_26_1760 ();
 sg13g2_decap_8 FILLER_26_1766 ();
 sg13g2_fill_1 FILLER_26_1773 ();
 sg13g2_decap_8 FILLER_26_1784 ();
 sg13g2_decap_4 FILLER_26_1791 ();
 sg13g2_fill_1 FILLER_26_1795 ();
 sg13g2_fill_1 FILLER_26_1822 ();
 sg13g2_fill_2 FILLER_26_1827 ();
 sg13g2_fill_2 FILLER_26_1860 ();
 sg13g2_decap_4 FILLER_26_1888 ();
 sg13g2_fill_2 FILLER_26_1919 ();
 sg13g2_decap_8 FILLER_26_1963 ();
 sg13g2_fill_1 FILLER_26_1979 ();
 sg13g2_fill_2 FILLER_26_2015 ();
 sg13g2_fill_1 FILLER_26_2017 ();
 sg13g2_fill_2 FILLER_26_2049 ();
 sg13g2_fill_1 FILLER_26_2051 ();
 sg13g2_fill_2 FILLER_26_2056 ();
 sg13g2_fill_1 FILLER_26_2058 ();
 sg13g2_fill_1 FILLER_26_2064 ();
 sg13g2_decap_8 FILLER_26_2081 ();
 sg13g2_decap_8 FILLER_26_2088 ();
 sg13g2_fill_1 FILLER_26_2095 ();
 sg13g2_decap_8 FILLER_26_2099 ();
 sg13g2_decap_4 FILLER_26_2106 ();
 sg13g2_fill_1 FILLER_26_2110 ();
 sg13g2_decap_8 FILLER_26_2116 ();
 sg13g2_decap_4 FILLER_26_2123 ();
 sg13g2_fill_2 FILLER_26_2127 ();
 sg13g2_fill_1 FILLER_26_2161 ();
 sg13g2_fill_1 FILLER_26_2168 ();
 sg13g2_fill_2 FILLER_26_2173 ();
 sg13g2_fill_1 FILLER_26_2182 ();
 sg13g2_fill_2 FILLER_26_2192 ();
 sg13g2_decap_8 FILLER_26_2247 ();
 sg13g2_decap_8 FILLER_26_2254 ();
 sg13g2_decap_4 FILLER_26_2261 ();
 sg13g2_fill_2 FILLER_26_2265 ();
 sg13g2_fill_2 FILLER_26_2282 ();
 sg13g2_decap_4 FILLER_26_2310 ();
 sg13g2_decap_8 FILLER_26_2336 ();
 sg13g2_decap_4 FILLER_26_2343 ();
 sg13g2_fill_2 FILLER_26_2347 ();
 sg13g2_decap_4 FILLER_26_2353 ();
 sg13g2_decap_8 FILLER_26_2362 ();
 sg13g2_decap_8 FILLER_26_2395 ();
 sg13g2_decap_8 FILLER_26_2402 ();
 sg13g2_decap_8 FILLER_26_2409 ();
 sg13g2_decap_8 FILLER_26_2416 ();
 sg13g2_decap_8 FILLER_26_2423 ();
 sg13g2_decap_8 FILLER_26_2430 ();
 sg13g2_decap_8 FILLER_26_2437 ();
 sg13g2_fill_1 FILLER_26_2536 ();
 sg13g2_decap_8 FILLER_26_2563 ();
 sg13g2_decap_8 FILLER_26_2570 ();
 sg13g2_decap_8 FILLER_26_2577 ();
 sg13g2_decap_8 FILLER_26_2584 ();
 sg13g2_decap_8 FILLER_26_2591 ();
 sg13g2_decap_8 FILLER_26_2598 ();
 sg13g2_decap_8 FILLER_26_2605 ();
 sg13g2_decap_8 FILLER_26_2612 ();
 sg13g2_decap_8 FILLER_26_2619 ();
 sg13g2_decap_8 FILLER_26_2626 ();
 sg13g2_decap_8 FILLER_26_2633 ();
 sg13g2_decap_8 FILLER_26_2640 ();
 sg13g2_decap_8 FILLER_26_2647 ();
 sg13g2_decap_8 FILLER_26_2654 ();
 sg13g2_decap_8 FILLER_26_2661 ();
 sg13g2_fill_2 FILLER_26_2668 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_55 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_decap_4 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_8 FILLER_27_110 ();
 sg13g2_decap_8 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_decap_4 FILLER_27_135 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_decap_4 FILLER_27_187 ();
 sg13g2_decap_4 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_4 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_301 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_decap_4 FILLER_27_374 ();
 sg13g2_decap_4 FILLER_27_386 ();
 sg13g2_fill_2 FILLER_27_395 ();
 sg13g2_decap_4 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_410 ();
 sg13g2_decap_4 FILLER_27_417 ();
 sg13g2_decap_8 FILLER_27_467 ();
 sg13g2_decap_8 FILLER_27_474 ();
 sg13g2_fill_1 FILLER_27_481 ();
 sg13g2_decap_4 FILLER_27_521 ();
 sg13g2_fill_1 FILLER_27_525 ();
 sg13g2_fill_1 FILLER_27_530 ();
 sg13g2_decap_8 FILLER_27_535 ();
 sg13g2_fill_2 FILLER_27_564 ();
 sg13g2_fill_2 FILLER_27_574 ();
 sg13g2_fill_1 FILLER_27_576 ();
 sg13g2_fill_1 FILLER_27_620 ();
 sg13g2_decap_4 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_635 ();
 sg13g2_fill_2 FILLER_27_642 ();
 sg13g2_fill_1 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_decap_8 FILLER_27_657 ();
 sg13g2_decap_8 FILLER_27_664 ();
 sg13g2_decap_8 FILLER_27_671 ();
 sg13g2_fill_1 FILLER_27_678 ();
 sg13g2_decap_8 FILLER_27_687 ();
 sg13g2_decap_8 FILLER_27_694 ();
 sg13g2_decap_8 FILLER_27_701 ();
 sg13g2_fill_2 FILLER_27_708 ();
 sg13g2_decap_4 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_4 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_813 ();
 sg13g2_decap_8 FILLER_27_820 ();
 sg13g2_decap_4 FILLER_27_827 ();
 sg13g2_fill_1 FILLER_27_831 ();
 sg13g2_fill_2 FILLER_27_837 ();
 sg13g2_fill_1 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_858 ();
 sg13g2_fill_1 FILLER_27_865 ();
 sg13g2_decap_4 FILLER_27_871 ();
 sg13g2_fill_1 FILLER_27_879 ();
 sg13g2_decap_4 FILLER_27_912 ();
 sg13g2_fill_2 FILLER_27_930 ();
 sg13g2_decap_8 FILLER_27_948 ();
 sg13g2_fill_2 FILLER_27_955 ();
 sg13g2_fill_2 FILLER_27_963 ();
 sg13g2_fill_2 FILLER_27_991 ();
 sg13g2_fill_1 FILLER_27_993 ();
 sg13g2_fill_1 FILLER_27_1000 ();
 sg13g2_fill_2 FILLER_27_1006 ();
 sg13g2_fill_1 FILLER_27_1008 ();
 sg13g2_decap_4 FILLER_27_1013 ();
 sg13g2_fill_1 FILLER_27_1052 ();
 sg13g2_decap_8 FILLER_27_1059 ();
 sg13g2_fill_2 FILLER_27_1071 ();
 sg13g2_decap_8 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1092 ();
 sg13g2_fill_1 FILLER_27_1099 ();
 sg13g2_fill_1 FILLER_27_1104 ();
 sg13g2_fill_2 FILLER_27_1110 ();
 sg13g2_fill_1 FILLER_27_1138 ();
 sg13g2_decap_4 FILLER_27_1174 ();
 sg13g2_fill_2 FILLER_27_1178 ();
 sg13g2_decap_4 FILLER_27_1222 ();
 sg13g2_fill_2 FILLER_27_1226 ();
 sg13g2_decap_8 FILLER_27_1241 ();
 sg13g2_decap_8 FILLER_27_1248 ();
 sg13g2_decap_8 FILLER_27_1255 ();
 sg13g2_fill_1 FILLER_27_1262 ();
 sg13g2_decap_8 FILLER_27_1272 ();
 sg13g2_fill_2 FILLER_27_1279 ();
 sg13g2_fill_1 FILLER_27_1281 ();
 sg13g2_fill_1 FILLER_27_1306 ();
 sg13g2_fill_2 FILLER_27_1325 ();
 sg13g2_decap_8 FILLER_27_1376 ();
 sg13g2_decap_8 FILLER_27_1383 ();
 sg13g2_decap_8 FILLER_27_1390 ();
 sg13g2_fill_1 FILLER_27_1397 ();
 sg13g2_fill_1 FILLER_27_1401 ();
 sg13g2_fill_2 FILLER_27_1408 ();
 sg13g2_fill_1 FILLER_27_1410 ();
 sg13g2_decap_4 FILLER_27_1416 ();
 sg13g2_fill_2 FILLER_27_1420 ();
 sg13g2_decap_8 FILLER_27_1430 ();
 sg13g2_decap_8 FILLER_27_1437 ();
 sg13g2_decap_8 FILLER_27_1444 ();
 sg13g2_decap_8 FILLER_27_1451 ();
 sg13g2_decap_8 FILLER_27_1468 ();
 sg13g2_decap_8 FILLER_27_1475 ();
 sg13g2_decap_8 FILLER_27_1482 ();
 sg13g2_decap_8 FILLER_27_1489 ();
 sg13g2_decap_4 FILLER_27_1496 ();
 sg13g2_fill_1 FILLER_27_1500 ();
 sg13g2_fill_1 FILLER_27_1509 ();
 sg13g2_decap_8 FILLER_27_1515 ();
 sg13g2_fill_2 FILLER_27_1522 ();
 sg13g2_fill_1 FILLER_27_1524 ();
 sg13g2_decap_8 FILLER_27_1577 ();
 sg13g2_fill_1 FILLER_27_1584 ();
 sg13g2_fill_1 FILLER_27_1600 ();
 sg13g2_decap_8 FILLER_27_1643 ();
 sg13g2_decap_8 FILLER_27_1650 ();
 sg13g2_decap_8 FILLER_27_1657 ();
 sg13g2_decap_8 FILLER_27_1664 ();
 sg13g2_decap_8 FILLER_27_1671 ();
 sg13g2_fill_2 FILLER_27_1682 ();
 sg13g2_fill_1 FILLER_27_1684 ();
 sg13g2_decap_4 FILLER_27_1728 ();
 sg13g2_fill_2 FILLER_27_1732 ();
 sg13g2_fill_2 FILLER_27_1739 ();
 sg13g2_fill_1 FILLER_27_1741 ();
 sg13g2_decap_4 FILLER_27_1794 ();
 sg13g2_decap_4 FILLER_27_1829 ();
 sg13g2_fill_2 FILLER_27_1833 ();
 sg13g2_fill_2 FILLER_27_1840 ();
 sg13g2_fill_1 FILLER_27_1842 ();
 sg13g2_fill_2 FILLER_27_1847 ();
 sg13g2_fill_1 FILLER_27_1849 ();
 sg13g2_fill_2 FILLER_27_1855 ();
 sg13g2_decap_8 FILLER_27_1868 ();
 sg13g2_fill_2 FILLER_27_1875 ();
 sg13g2_decap_4 FILLER_27_1882 ();
 sg13g2_fill_1 FILLER_27_1891 ();
 sg13g2_decap_4 FILLER_27_1930 ();
 sg13g2_decap_8 FILLER_27_1938 ();
 sg13g2_decap_8 FILLER_27_1945 ();
 sg13g2_fill_2 FILLER_27_1952 ();
 sg13g2_fill_1 FILLER_27_1954 ();
 sg13g2_decap_8 FILLER_27_1960 ();
 sg13g2_decap_8 FILLER_27_1967 ();
 sg13g2_fill_2 FILLER_27_2004 ();
 sg13g2_decap_8 FILLER_27_2078 ();
 sg13g2_decap_8 FILLER_27_2085 ();
 sg13g2_decap_4 FILLER_27_2092 ();
 sg13g2_decap_8 FILLER_27_2102 ();
 sg13g2_fill_1 FILLER_27_2109 ();
 sg13g2_decap_8 FILLER_27_2114 ();
 sg13g2_fill_2 FILLER_27_2121 ();
 sg13g2_fill_2 FILLER_27_2133 ();
 sg13g2_fill_1 FILLER_27_2135 ();
 sg13g2_fill_1 FILLER_27_2150 ();
 sg13g2_fill_1 FILLER_27_2163 ();
 sg13g2_decap_4 FILLER_27_2216 ();
 sg13g2_decap_8 FILLER_27_2226 ();
 sg13g2_decap_8 FILLER_27_2270 ();
 sg13g2_fill_2 FILLER_27_2277 ();
 sg13g2_fill_1 FILLER_27_2288 ();
 sg13g2_decap_8 FILLER_27_2295 ();
 sg13g2_decap_8 FILLER_27_2302 ();
 sg13g2_fill_2 FILLER_27_2309 ();
 sg13g2_decap_8 FILLER_27_2314 ();
 sg13g2_decap_8 FILLER_27_2326 ();
 sg13g2_decap_8 FILLER_27_2333 ();
 sg13g2_decap_8 FILLER_27_2340 ();
 sg13g2_fill_2 FILLER_27_2347 ();
 sg13g2_fill_2 FILLER_27_2380 ();
 sg13g2_decap_8 FILLER_27_2400 ();
 sg13g2_decap_8 FILLER_27_2407 ();
 sg13g2_decap_8 FILLER_27_2414 ();
 sg13g2_decap_4 FILLER_27_2421 ();
 sg13g2_fill_2 FILLER_27_2494 ();
 sg13g2_fill_1 FILLER_27_2500 ();
 sg13g2_fill_2 FILLER_27_2511 ();
 sg13g2_fill_1 FILLER_27_2513 ();
 sg13g2_decap_8 FILLER_27_2567 ();
 sg13g2_decap_8 FILLER_27_2574 ();
 sg13g2_decap_8 FILLER_27_2581 ();
 sg13g2_decap_8 FILLER_27_2588 ();
 sg13g2_decap_8 FILLER_27_2595 ();
 sg13g2_decap_8 FILLER_27_2602 ();
 sg13g2_decap_8 FILLER_27_2609 ();
 sg13g2_decap_8 FILLER_27_2616 ();
 sg13g2_decap_8 FILLER_27_2623 ();
 sg13g2_decap_8 FILLER_27_2630 ();
 sg13g2_decap_8 FILLER_27_2637 ();
 sg13g2_decap_8 FILLER_27_2644 ();
 sg13g2_decap_8 FILLER_27_2651 ();
 sg13g2_decap_8 FILLER_27_2658 ();
 sg13g2_decap_4 FILLER_27_2665 ();
 sg13g2_fill_1 FILLER_27_2669 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_11 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_90 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_fill_1 FILLER_28_390 ();
 sg13g2_fill_1 FILLER_28_404 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_4 FILLER_28_481 ();
 sg13g2_decap_8 FILLER_28_505 ();
 sg13g2_fill_2 FILLER_28_512 ();
 sg13g2_fill_1 FILLER_28_514 ();
 sg13g2_decap_8 FILLER_28_520 ();
 sg13g2_fill_1 FILLER_28_532 ();
 sg13g2_fill_2 FILLER_28_541 ();
 sg13g2_fill_2 FILLER_28_554 ();
 sg13g2_fill_2 FILLER_28_561 ();
 sg13g2_fill_1 FILLER_28_571 ();
 sg13g2_fill_2 FILLER_28_580 ();
 sg13g2_decap_4 FILLER_28_610 ();
 sg13g2_fill_1 FILLER_28_614 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_8 FILLER_28_636 ();
 sg13g2_decap_4 FILLER_28_669 ();
 sg13g2_fill_2 FILLER_28_673 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_fill_1 FILLER_28_728 ();
 sg13g2_fill_1 FILLER_28_742 ();
 sg13g2_decap_4 FILLER_28_747 ();
 sg13g2_fill_1 FILLER_28_751 ();
 sg13g2_fill_2 FILLER_28_756 ();
 sg13g2_fill_1 FILLER_28_847 ();
 sg13g2_fill_1 FILLER_28_856 ();
 sg13g2_fill_1 FILLER_28_883 ();
 sg13g2_fill_1 FILLER_28_892 ();
 sg13g2_fill_2 FILLER_28_899 ();
 sg13g2_fill_1 FILLER_28_927 ();
 sg13g2_fill_2 FILLER_28_954 ();
 sg13g2_fill_2 FILLER_28_998 ();
 sg13g2_fill_1 FILLER_28_1016 ();
 sg13g2_fill_1 FILLER_28_1022 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_fill_1 FILLER_28_1029 ();
 sg13g2_fill_2 FILLER_28_1039 ();
 sg13g2_fill_1 FILLER_28_1041 ();
 sg13g2_decap_4 FILLER_28_1077 ();
 sg13g2_decap_8 FILLER_28_1096 ();
 sg13g2_decap_8 FILLER_28_1103 ();
 sg13g2_decap_8 FILLER_28_1110 ();
 sg13g2_decap_8 FILLER_28_1117 ();
 sg13g2_decap_4 FILLER_28_1124 ();
 sg13g2_fill_1 FILLER_28_1128 ();
 sg13g2_decap_4 FILLER_28_1138 ();
 sg13g2_fill_1 FILLER_28_1147 ();
 sg13g2_decap_8 FILLER_28_1152 ();
 sg13g2_decap_8 FILLER_28_1159 ();
 sg13g2_decap_8 FILLER_28_1166 ();
 sg13g2_fill_1 FILLER_28_1173 ();
 sg13g2_decap_4 FILLER_28_1189 ();
 sg13g2_decap_8 FILLER_28_1242 ();
 sg13g2_decap_8 FILLER_28_1249 ();
 sg13g2_decap_8 FILLER_28_1256 ();
 sg13g2_decap_8 FILLER_28_1263 ();
 sg13g2_decap_8 FILLER_28_1270 ();
 sg13g2_fill_2 FILLER_28_1277 ();
 sg13g2_fill_1 FILLER_28_1300 ();
 sg13g2_fill_2 FILLER_28_1322 ();
 sg13g2_fill_1 FILLER_28_1324 ();
 sg13g2_decap_8 FILLER_28_1329 ();
 sg13g2_decap_4 FILLER_28_1336 ();
 sg13g2_fill_2 FILLER_28_1340 ();
 sg13g2_decap_8 FILLER_28_1372 ();
 sg13g2_decap_8 FILLER_28_1379 ();
 sg13g2_fill_2 FILLER_28_1386 ();
 sg13g2_fill_1 FILLER_28_1405 ();
 sg13g2_decap_8 FILLER_28_1437 ();
 sg13g2_decap_8 FILLER_28_1444 ();
 sg13g2_decap_4 FILLER_28_1451 ();
 sg13g2_decap_8 FILLER_28_1481 ();
 sg13g2_decap_8 FILLER_28_1488 ();
 sg13g2_fill_2 FILLER_28_1495 ();
 sg13g2_decap_4 FILLER_28_1510 ();
 sg13g2_decap_4 FILLER_28_1533 ();
 sg13g2_fill_1 FILLER_28_1546 ();
 sg13g2_fill_2 FILLER_28_1560 ();
 sg13g2_fill_2 FILLER_28_1575 ();
 sg13g2_decap_8 FILLER_28_1582 ();
 sg13g2_fill_2 FILLER_28_1589 ();
 sg13g2_fill_2 FILLER_28_1595 ();
 sg13g2_fill_2 FILLER_28_1608 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_decap_8 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1652 ();
 sg13g2_decap_8 FILLER_28_1659 ();
 sg13g2_decap_8 FILLER_28_1666 ();
 sg13g2_decap_8 FILLER_28_1673 ();
 sg13g2_decap_8 FILLER_28_1680 ();
 sg13g2_fill_2 FILLER_28_1733 ();
 sg13g2_fill_2 FILLER_28_1761 ();
 sg13g2_fill_2 FILLER_28_1776 ();
 sg13g2_decap_8 FILLER_28_1787 ();
 sg13g2_fill_2 FILLER_28_1799 ();
 sg13g2_fill_1 FILLER_28_1801 ();
 sg13g2_decap_4 FILLER_28_1811 ();
 sg13g2_fill_1 FILLER_28_1815 ();
 sg13g2_decap_8 FILLER_28_1826 ();
 sg13g2_decap_8 FILLER_28_1833 ();
 sg13g2_fill_1 FILLER_28_1883 ();
 sg13g2_decap_8 FILLER_28_1896 ();
 sg13g2_decap_8 FILLER_28_1903 ();
 sg13g2_decap_4 FILLER_28_1910 ();
 sg13g2_decap_8 FILLER_28_1926 ();
 sg13g2_fill_2 FILLER_28_1933 ();
 sg13g2_fill_1 FILLER_28_1935 ();
 sg13g2_decap_4 FILLER_28_1941 ();
 sg13g2_fill_1 FILLER_28_1945 ();
 sg13g2_decap_8 FILLER_28_1964 ();
 sg13g2_decap_8 FILLER_28_1971 ();
 sg13g2_fill_2 FILLER_28_1978 ();
 sg13g2_decap_4 FILLER_28_1985 ();
 sg13g2_fill_1 FILLER_28_1989 ();
 sg13g2_decap_4 FILLER_28_1995 ();
 sg13g2_decap_4 FILLER_28_2042 ();
 sg13g2_fill_2 FILLER_28_2051 ();
 sg13g2_fill_1 FILLER_28_2053 ();
 sg13g2_fill_2 FILLER_28_2084 ();
 sg13g2_fill_1 FILLER_28_2086 ();
 sg13g2_decap_4 FILLER_28_2095 ();
 sg13g2_fill_2 FILLER_28_2099 ();
 sg13g2_decap_4 FILLER_28_2109 ();
 sg13g2_decap_8 FILLER_28_2228 ();
 sg13g2_fill_1 FILLER_28_2235 ();
 sg13g2_fill_1 FILLER_28_2241 ();
 sg13g2_fill_2 FILLER_28_2246 ();
 sg13g2_fill_1 FILLER_28_2248 ();
 sg13g2_decap_8 FILLER_28_2275 ();
 sg13g2_fill_1 FILLER_28_2282 ();
 sg13g2_decap_8 FILLER_28_2295 ();
 sg13g2_fill_2 FILLER_28_2317 ();
 sg13g2_decap_8 FILLER_28_2349 ();
 sg13g2_decap_8 FILLER_28_2356 ();
 sg13g2_decap_8 FILLER_28_2363 ();
 sg13g2_decap_8 FILLER_28_2422 ();
 sg13g2_decap_4 FILLER_28_2429 ();
 sg13g2_fill_2 FILLER_28_2433 ();
 sg13g2_decap_8 FILLER_28_2506 ();
 sg13g2_fill_2 FILLER_28_2513 ();
 sg13g2_fill_1 FILLER_28_2537 ();
 sg13g2_decap_8 FILLER_28_2564 ();
 sg13g2_decap_8 FILLER_28_2571 ();
 sg13g2_decap_8 FILLER_28_2578 ();
 sg13g2_decap_8 FILLER_28_2585 ();
 sg13g2_decap_8 FILLER_28_2592 ();
 sg13g2_decap_8 FILLER_28_2599 ();
 sg13g2_decap_8 FILLER_28_2606 ();
 sg13g2_decap_8 FILLER_28_2613 ();
 sg13g2_decap_8 FILLER_28_2620 ();
 sg13g2_decap_8 FILLER_28_2627 ();
 sg13g2_decap_8 FILLER_28_2634 ();
 sg13g2_decap_8 FILLER_28_2641 ();
 sg13g2_decap_8 FILLER_28_2648 ();
 sg13g2_decap_8 FILLER_28_2655 ();
 sg13g2_decap_8 FILLER_28_2662 ();
 sg13g2_fill_1 FILLER_28_2669 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_11 ();
 sg13g2_fill_2 FILLER_29_31 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_decap_4 FILLER_29_145 ();
 sg13g2_decap_4 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_4 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_229 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_4 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_decap_4 FILLER_29_359 ();
 sg13g2_decap_4 FILLER_29_371 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_fill_2 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_475 ();
 sg13g2_decap_8 FILLER_29_482 ();
 sg13g2_decap_8 FILLER_29_489 ();
 sg13g2_decap_8 FILLER_29_496 ();
 sg13g2_decap_8 FILLER_29_503 ();
 sg13g2_decap_4 FILLER_29_510 ();
 sg13g2_fill_2 FILLER_29_514 ();
 sg13g2_fill_2 FILLER_29_521 ();
 sg13g2_fill_1 FILLER_29_523 ();
 sg13g2_fill_1 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_fill_2 FILLER_29_571 ();
 sg13g2_fill_1 FILLER_29_573 ();
 sg13g2_decap_8 FILLER_29_582 ();
 sg13g2_fill_2 FILLER_29_589 ();
 sg13g2_decap_4 FILLER_29_602 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_decap_8 FILLER_29_657 ();
 sg13g2_decap_8 FILLER_29_668 ();
 sg13g2_decap_4 FILLER_29_675 ();
 sg13g2_fill_1 FILLER_29_679 ();
 sg13g2_fill_2 FILLER_29_684 ();
 sg13g2_fill_2 FILLER_29_691 ();
 sg13g2_decap_8 FILLER_29_719 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_fill_1 FILLER_29_733 ();
 sg13g2_decap_4 FILLER_29_738 ();
 sg13g2_fill_1 FILLER_29_742 ();
 sg13g2_fill_1 FILLER_29_748 ();
 sg13g2_fill_1 FILLER_29_779 ();
 sg13g2_fill_1 FILLER_29_784 ();
 sg13g2_decap_4 FILLER_29_789 ();
 sg13g2_fill_1 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_4 FILLER_29_812 ();
 sg13g2_fill_2 FILLER_29_816 ();
 sg13g2_decap_4 FILLER_29_852 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_fill_1 FILLER_29_862 ();
 sg13g2_fill_2 FILLER_29_867 ();
 sg13g2_fill_1 FILLER_29_869 ();
 sg13g2_fill_1 FILLER_29_896 ();
 sg13g2_fill_2 FILLER_29_927 ();
 sg13g2_fill_2 FILLER_29_933 ();
 sg13g2_fill_1 FILLER_29_935 ();
 sg13g2_fill_2 FILLER_29_953 ();
 sg13g2_fill_1 FILLER_29_973 ();
 sg13g2_decap_4 FILLER_29_983 ();
 sg13g2_fill_1 FILLER_29_987 ();
 sg13g2_fill_1 FILLER_29_993 ();
 sg13g2_fill_2 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1028 ();
 sg13g2_fill_2 FILLER_29_1035 ();
 sg13g2_decap_8 FILLER_29_1042 ();
 sg13g2_decap_8 FILLER_29_1049 ();
 sg13g2_decap_4 FILLER_29_1056 ();
 sg13g2_fill_2 FILLER_29_1060 ();
 sg13g2_decap_4 FILLER_29_1067 ();
 sg13g2_fill_2 FILLER_29_1071 ();
 sg13g2_decap_8 FILLER_29_1085 ();
 sg13g2_decap_8 FILLER_29_1092 ();
 sg13g2_fill_1 FILLER_29_1099 ();
 sg13g2_decap_4 FILLER_29_1105 ();
 sg13g2_fill_2 FILLER_29_1109 ();
 sg13g2_fill_1 FILLER_29_1122 ();
 sg13g2_decap_4 FILLER_29_1130 ();
 sg13g2_decap_4 FILLER_29_1144 ();
 sg13g2_decap_8 FILLER_29_1183 ();
 sg13g2_decap_8 FILLER_29_1190 ();
 sg13g2_decap_4 FILLER_29_1197 ();
 sg13g2_decap_4 FILLER_29_1206 ();
 sg13g2_decap_4 FILLER_29_1240 ();
 sg13g2_fill_1 FILLER_29_1244 ();
 sg13g2_fill_2 FILLER_29_1297 ();
 sg13g2_fill_1 FILLER_29_1299 ();
 sg13g2_decap_8 FILLER_29_1326 ();
 sg13g2_decap_4 FILLER_29_1333 ();
 sg13g2_fill_2 FILLER_29_1337 ();
 sg13g2_fill_2 FILLER_29_1362 ();
 sg13g2_fill_1 FILLER_29_1364 ();
 sg13g2_decap_8 FILLER_29_1420 ();
 sg13g2_decap_8 FILLER_29_1466 ();
 sg13g2_fill_2 FILLER_29_1473 ();
 sg13g2_fill_2 FILLER_29_1501 ();
 sg13g2_fill_1 FILLER_29_1503 ();
 sg13g2_fill_2 FILLER_29_1543 ();
 sg13g2_fill_1 FILLER_29_1545 ();
 sg13g2_fill_2 FILLER_29_1587 ();
 sg13g2_fill_1 FILLER_29_1589 ();
 sg13g2_fill_2 FILLER_29_1613 ();
 sg13g2_decap_8 FILLER_29_1641 ();
 sg13g2_decap_8 FILLER_29_1648 ();
 sg13g2_fill_2 FILLER_29_1655 ();
 sg13g2_fill_1 FILLER_29_1657 ();
 sg13g2_decap_8 FILLER_29_1673 ();
 sg13g2_decap_8 FILLER_29_1680 ();
 sg13g2_fill_1 FILLER_29_1687 ();
 sg13g2_fill_1 FILLER_29_1706 ();
 sg13g2_fill_2 FILLER_29_1733 ();
 sg13g2_fill_1 FILLER_29_1735 ();
 sg13g2_fill_2 FILLER_29_1741 ();
 sg13g2_fill_1 FILLER_29_1769 ();
 sg13g2_decap_4 FILLER_29_1782 ();
 sg13g2_fill_1 FILLER_29_1791 ();
 sg13g2_fill_1 FILLER_29_1812 ();
 sg13g2_decap_8 FILLER_29_1839 ();
 sg13g2_fill_2 FILLER_29_1846 ();
 sg13g2_fill_1 FILLER_29_1848 ();
 sg13g2_decap_8 FILLER_29_1867 ();
 sg13g2_decap_8 FILLER_29_1874 ();
 sg13g2_fill_2 FILLER_29_1881 ();
 sg13g2_fill_1 FILLER_29_1883 ();
 sg13g2_fill_1 FILLER_29_1927 ();
 sg13g2_fill_2 FILLER_29_1933 ();
 sg13g2_fill_1 FILLER_29_1935 ();
 sg13g2_fill_1 FILLER_29_1971 ();
 sg13g2_fill_2 FILLER_29_1980 ();
 sg13g2_fill_1 FILLER_29_1982 ();
 sg13g2_decap_4 FILLER_29_1988 ();
 sg13g2_fill_2 FILLER_29_1992 ();
 sg13g2_fill_2 FILLER_29_2006 ();
 sg13g2_fill_1 FILLER_29_2013 ();
 sg13g2_fill_2 FILLER_29_2040 ();
 sg13g2_decap_8 FILLER_29_2073 ();
 sg13g2_fill_2 FILLER_29_2085 ();
 sg13g2_fill_2 FILLER_29_2120 ();
 sg13g2_fill_2 FILLER_29_2168 ();
 sg13g2_decap_4 FILLER_29_2208 ();
 sg13g2_fill_2 FILLER_29_2212 ();
 sg13g2_decap_4 FILLER_29_2253 ();
 sg13g2_fill_1 FILLER_29_2261 ();
 sg13g2_decap_4 FILLER_29_2293 ();
 sg13g2_fill_2 FILLER_29_2305 ();
 sg13g2_fill_1 FILLER_29_2314 ();
 sg13g2_fill_1 FILLER_29_2346 ();
 sg13g2_fill_1 FILLER_29_2351 ();
 sg13g2_decap_8 FILLER_29_2392 ();
 sg13g2_decap_8 FILLER_29_2399 ();
 sg13g2_fill_1 FILLER_29_2406 ();
 sg13g2_decap_8 FILLER_29_2413 ();
 sg13g2_decap_8 FILLER_29_2420 ();
 sg13g2_decap_8 FILLER_29_2427 ();
 sg13g2_fill_1 FILLER_29_2434 ();
 sg13g2_fill_2 FILLER_29_2439 ();
 sg13g2_fill_2 FILLER_29_2467 ();
 sg13g2_fill_2 FILLER_29_2473 ();
 sg13g2_decap_8 FILLER_29_2501 ();
 sg13g2_fill_2 FILLER_29_2508 ();
 sg13g2_fill_2 FILLER_29_2544 ();
 sg13g2_decap_8 FILLER_29_2554 ();
 sg13g2_decap_8 FILLER_29_2561 ();
 sg13g2_decap_8 FILLER_29_2568 ();
 sg13g2_decap_8 FILLER_29_2575 ();
 sg13g2_decap_8 FILLER_29_2582 ();
 sg13g2_decap_8 FILLER_29_2589 ();
 sg13g2_decap_8 FILLER_29_2596 ();
 sg13g2_decap_8 FILLER_29_2603 ();
 sg13g2_decap_8 FILLER_29_2610 ();
 sg13g2_decap_8 FILLER_29_2617 ();
 sg13g2_decap_8 FILLER_29_2624 ();
 sg13g2_decap_8 FILLER_29_2631 ();
 sg13g2_decap_8 FILLER_29_2638 ();
 sg13g2_decap_8 FILLER_29_2645 ();
 sg13g2_decap_8 FILLER_29_2652 ();
 sg13g2_decap_8 FILLER_29_2659 ();
 sg13g2_decap_4 FILLER_29_2666 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_decap_8 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_40 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_61 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_decap_8 FILLER_30_142 ();
 sg13g2_decap_8 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_4 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_4 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_4 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_decap_4 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_429 ();
 sg13g2_decap_4 FILLER_30_436 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_fill_1 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_503 ();
 sg13g2_decap_8 FILLER_30_510 ();
 sg13g2_decap_8 FILLER_30_517 ();
 sg13g2_fill_2 FILLER_30_524 ();
 sg13g2_fill_1 FILLER_30_538 ();
 sg13g2_decap_4 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_fill_1 FILLER_30_574 ();
 sg13g2_fill_1 FILLER_30_583 ();
 sg13g2_fill_1 FILLER_30_592 ();
 sg13g2_fill_2 FILLER_30_601 ();
 sg13g2_fill_2 FILLER_30_608 ();
 sg13g2_fill_2 FILLER_30_619 ();
 sg13g2_decap_8 FILLER_30_629 ();
 sg13g2_decap_4 FILLER_30_641 ();
 sg13g2_fill_1 FILLER_30_645 ();
 sg13g2_fill_2 FILLER_30_649 ();
 sg13g2_decap_4 FILLER_30_656 ();
 sg13g2_fill_1 FILLER_30_660 ();
 sg13g2_decap_8 FILLER_30_675 ();
 sg13g2_decap_8 FILLER_30_682 ();
 sg13g2_fill_2 FILLER_30_689 ();
 sg13g2_fill_1 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_722 ();
 sg13g2_decap_8 FILLER_30_729 ();
 sg13g2_decap_8 FILLER_30_736 ();
 sg13g2_fill_2 FILLER_30_743 ();
 sg13g2_fill_1 FILLER_30_745 ();
 sg13g2_decap_8 FILLER_30_794 ();
 sg13g2_decap_8 FILLER_30_801 ();
 sg13g2_decap_8 FILLER_30_808 ();
 sg13g2_decap_8 FILLER_30_815 ();
 sg13g2_decap_4 FILLER_30_822 ();
 sg13g2_fill_2 FILLER_30_826 ();
 sg13g2_decap_4 FILLER_30_838 ();
 sg13g2_fill_2 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_874 ();
 sg13g2_fill_1 FILLER_30_881 ();
 sg13g2_fill_1 FILLER_30_887 ();
 sg13g2_fill_2 FILLER_30_894 ();
 sg13g2_fill_1 FILLER_30_900 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_fill_2 FILLER_30_931 ();
 sg13g2_fill_2 FILLER_30_974 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1007 ();
 sg13g2_decap_4 FILLER_30_1014 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_fill_2 FILLER_30_1029 ();
 sg13g2_fill_2 FILLER_30_1063 ();
 sg13g2_fill_1 FILLER_30_1065 ();
 sg13g2_fill_2 FILLER_30_1090 ();
 sg13g2_decap_4 FILLER_30_1096 ();
 sg13g2_decap_8 FILLER_30_1108 ();
 sg13g2_decap_4 FILLER_30_1115 ();
 sg13g2_fill_2 FILLER_30_1128 ();
 sg13g2_decap_8 FILLER_30_1141 ();
 sg13g2_decap_8 FILLER_30_1148 ();
 sg13g2_decap_8 FILLER_30_1155 ();
 sg13g2_fill_1 FILLER_30_1162 ();
 sg13g2_fill_2 FILLER_30_1177 ();
 sg13g2_fill_1 FILLER_30_1179 ();
 sg13g2_decap_8 FILLER_30_1210 ();
 sg13g2_decap_8 FILLER_30_1217 ();
 sg13g2_fill_2 FILLER_30_1224 ();
 sg13g2_fill_2 FILLER_30_1238 ();
 sg13g2_decap_8 FILLER_30_1245 ();
 sg13g2_decap_4 FILLER_30_1264 ();
 sg13g2_fill_1 FILLER_30_1268 ();
 sg13g2_decap_8 FILLER_30_1273 ();
 sg13g2_fill_1 FILLER_30_1280 ();
 sg13g2_decap_8 FILLER_30_1312 ();
 sg13g2_decap_8 FILLER_30_1319 ();
 sg13g2_decap_8 FILLER_30_1326 ();
 sg13g2_decap_8 FILLER_30_1338 ();
 sg13g2_fill_1 FILLER_30_1345 ();
 sg13g2_decap_4 FILLER_30_1350 ();
 sg13g2_fill_1 FILLER_30_1354 ();
 sg13g2_fill_2 FILLER_30_1397 ();
 sg13g2_decap_4 FILLER_30_1409 ();
 sg13g2_fill_1 FILLER_30_1413 ();
 sg13g2_decap_4 FILLER_30_1419 ();
 sg13g2_fill_1 FILLER_30_1423 ();
 sg13g2_decap_8 FILLER_30_1429 ();
 sg13g2_fill_2 FILLER_30_1436 ();
 sg13g2_fill_1 FILLER_30_1438 ();
 sg13g2_fill_1 FILLER_30_1443 ();
 sg13g2_fill_2 FILLER_30_1478 ();
 sg13g2_decap_8 FILLER_30_1485 ();
 sg13g2_decap_8 FILLER_30_1492 ();
 sg13g2_fill_2 FILLER_30_1499 ();
 sg13g2_fill_1 FILLER_30_1501 ();
 sg13g2_fill_2 FILLER_30_1511 ();
 sg13g2_fill_1 FILLER_30_1513 ();
 sg13g2_fill_1 FILLER_30_1535 ();
 sg13g2_fill_2 FILLER_30_1588 ();
 sg13g2_fill_1 FILLER_30_1590 ();
 sg13g2_fill_1 FILLER_30_1655 ();
 sg13g2_fill_1 FILLER_30_1662 ();
 sg13g2_fill_1 FILLER_30_1689 ();
 sg13g2_fill_2 FILLER_30_1694 ();
 sg13g2_fill_2 FILLER_30_1701 ();
 sg13g2_decap_8 FILLER_30_1707 ();
 sg13g2_fill_2 FILLER_30_1714 ();
 sg13g2_fill_1 FILLER_30_1768 ();
 sg13g2_fill_2 FILLER_30_1773 ();
 sg13g2_fill_1 FILLER_30_1775 ();
 sg13g2_fill_1 FILLER_30_1802 ();
 sg13g2_decap_4 FILLER_30_1809 ();
 sg13g2_decap_4 FILLER_30_1839 ();
 sg13g2_decap_8 FILLER_30_1868 ();
 sg13g2_decap_8 FILLER_30_1875 ();
 sg13g2_decap_8 FILLER_30_1882 ();
 sg13g2_fill_2 FILLER_30_1889 ();
 sg13g2_decap_8 FILLER_30_1899 ();
 sg13g2_fill_2 FILLER_30_1906 ();
 sg13g2_fill_1 FILLER_30_1908 ();
 sg13g2_decap_8 FILLER_30_1935 ();
 sg13g2_fill_2 FILLER_30_1942 ();
 sg13g2_decap_8 FILLER_30_1950 ();
 sg13g2_decap_8 FILLER_30_1957 ();
 sg13g2_decap_8 FILLER_30_1964 ();
 sg13g2_fill_1 FILLER_30_1971 ();
 sg13g2_decap_8 FILLER_30_1976 ();
 sg13g2_decap_8 FILLER_30_1983 ();
 sg13g2_decap_8 FILLER_30_1990 ();
 sg13g2_fill_1 FILLER_30_1997 ();
 sg13g2_decap_4 FILLER_30_2002 ();
 sg13g2_fill_2 FILLER_30_2006 ();
 sg13g2_decap_4 FILLER_30_2021 ();
 sg13g2_decap_8 FILLER_30_2029 ();
 sg13g2_fill_1 FILLER_30_2044 ();
 sg13g2_decap_4 FILLER_30_2055 ();
 sg13g2_fill_1 FILLER_30_2063 ();
 sg13g2_decap_8 FILLER_30_2090 ();
 sg13g2_decap_8 FILLER_30_2097 ();
 sg13g2_decap_4 FILLER_30_2104 ();
 sg13g2_fill_1 FILLER_30_2108 ();
 sg13g2_fill_2 FILLER_30_2145 ();
 sg13g2_decap_8 FILLER_30_2196 ();
 sg13g2_decap_8 FILLER_30_2203 ();
 sg13g2_decap_8 FILLER_30_2210 ();
 sg13g2_decap_8 FILLER_30_2217 ();
 sg13g2_decap_4 FILLER_30_2224 ();
 sg13g2_fill_1 FILLER_30_2228 ();
 sg13g2_decap_4 FILLER_30_2259 ();
 sg13g2_fill_1 FILLER_30_2263 ();
 sg13g2_decap_8 FILLER_30_2268 ();
 sg13g2_decap_8 FILLER_30_2275 ();
 sg13g2_decap_8 FILLER_30_2282 ();
 sg13g2_fill_1 FILLER_30_2294 ();
 sg13g2_decap_4 FILLER_30_2300 ();
 sg13g2_fill_1 FILLER_30_2304 ();
 sg13g2_decap_8 FILLER_30_2309 ();
 sg13g2_decap_8 FILLER_30_2316 ();
 sg13g2_decap_8 FILLER_30_2323 ();
 sg13g2_decap_8 FILLER_30_2330 ();
 sg13g2_fill_2 FILLER_30_2337 ();
 sg13g2_fill_1 FILLER_30_2339 ();
 sg13g2_decap_8 FILLER_30_2392 ();
 sg13g2_decap_8 FILLER_30_2399 ();
 sg13g2_decap_8 FILLER_30_2406 ();
 sg13g2_decap_8 FILLER_30_2413 ();
 sg13g2_decap_4 FILLER_30_2420 ();
 sg13g2_fill_1 FILLER_30_2424 ();
 sg13g2_fill_2 FILLER_30_2469 ();
 sg13g2_fill_2 FILLER_30_2475 ();
 sg13g2_fill_1 FILLER_30_2503 ();
 sg13g2_decap_8 FILLER_30_2508 ();
 sg13g2_decap_4 FILLER_30_2515 ();
 sg13g2_decap_8 FILLER_30_2549 ();
 sg13g2_decap_8 FILLER_30_2556 ();
 sg13g2_decap_8 FILLER_30_2563 ();
 sg13g2_decap_8 FILLER_30_2570 ();
 sg13g2_decap_8 FILLER_30_2577 ();
 sg13g2_decap_8 FILLER_30_2584 ();
 sg13g2_decap_8 FILLER_30_2591 ();
 sg13g2_decap_8 FILLER_30_2598 ();
 sg13g2_decap_8 FILLER_30_2605 ();
 sg13g2_decap_8 FILLER_30_2612 ();
 sg13g2_decap_8 FILLER_30_2619 ();
 sg13g2_decap_8 FILLER_30_2626 ();
 sg13g2_decap_8 FILLER_30_2633 ();
 sg13g2_decap_8 FILLER_30_2640 ();
 sg13g2_decap_8 FILLER_30_2647 ();
 sg13g2_decap_8 FILLER_30_2654 ();
 sg13g2_decap_8 FILLER_30_2661 ();
 sg13g2_fill_2 FILLER_30_2668 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_27 ();
 sg13g2_decap_8 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_40 ();
 sg13g2_decap_4 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_191 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_4 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_299 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_decap_8 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_2 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_8 FILLER_31_404 ();
 sg13g2_decap_8 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_8 FILLER_31_425 ();
 sg13g2_decap_8 FILLER_31_436 ();
 sg13g2_decap_8 FILLER_31_474 ();
 sg13g2_decap_8 FILLER_31_481 ();
 sg13g2_fill_1 FILLER_31_510 ();
 sg13g2_decap_8 FILLER_31_516 ();
 sg13g2_decap_4 FILLER_31_523 ();
 sg13g2_fill_2 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_4 FILLER_31_556 ();
 sg13g2_fill_1 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_571 ();
 sg13g2_fill_1 FILLER_31_578 ();
 sg13g2_decap_8 FILLER_31_592 ();
 sg13g2_decap_8 FILLER_31_599 ();
 sg13g2_fill_1 FILLER_31_606 ();
 sg13g2_decap_4 FILLER_31_622 ();
 sg13g2_decap_4 FILLER_31_629 ();
 sg13g2_fill_1 FILLER_31_633 ();
 sg13g2_fill_1 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_fill_1 FILLER_31_711 ();
 sg13g2_fill_1 FILLER_31_742 ();
 sg13g2_fill_1 FILLER_31_754 ();
 sg13g2_fill_2 FILLER_31_765 ();
 sg13g2_fill_1 FILLER_31_771 ();
 sg13g2_fill_1 FILLER_31_789 ();
 sg13g2_fill_2 FILLER_31_802 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_fill_1 FILLER_31_839 ();
 sg13g2_decap_4 FILLER_31_866 ();
 sg13g2_fill_2 FILLER_31_894 ();
 sg13g2_decap_8 FILLER_31_900 ();
 sg13g2_fill_2 FILLER_31_907 ();
 sg13g2_decap_8 FILLER_31_914 ();
 sg13g2_decap_4 FILLER_31_921 ();
 sg13g2_decap_4 FILLER_31_930 ();
 sg13g2_decap_4 FILLER_31_938 ();
 sg13g2_decap_4 FILLER_31_972 ();
 sg13g2_decap_8 FILLER_31_988 ();
 sg13g2_decap_8 FILLER_31_995 ();
 sg13g2_decap_8 FILLER_31_1002 ();
 sg13g2_decap_4 FILLER_31_1009 ();
 sg13g2_decap_4 FILLER_31_1017 ();
 sg13g2_fill_2 FILLER_31_1021 ();
 sg13g2_decap_8 FILLER_31_1031 ();
 sg13g2_fill_2 FILLER_31_1038 ();
 sg13g2_fill_1 FILLER_31_1040 ();
 sg13g2_decap_8 FILLER_31_1067 ();
 sg13g2_decap_4 FILLER_31_1074 ();
 sg13g2_fill_1 FILLER_31_1078 ();
 sg13g2_fill_1 FILLER_31_1136 ();
 sg13g2_decap_8 FILLER_31_1183 ();
 sg13g2_decap_8 FILLER_31_1193 ();
 sg13g2_decap_4 FILLER_31_1200 ();
 sg13g2_fill_2 FILLER_31_1204 ();
 sg13g2_decap_8 FILLER_31_1247 ();
 sg13g2_decap_8 FILLER_31_1254 ();
 sg13g2_fill_2 FILLER_31_1261 ();
 sg13g2_fill_1 FILLER_31_1263 ();
 sg13g2_fill_2 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1277 ();
 sg13g2_decap_4 FILLER_31_1284 ();
 sg13g2_fill_2 FILLER_31_1302 ();
 sg13g2_fill_1 FILLER_31_1367 ();
 sg13g2_fill_2 FILLER_31_1372 ();
 sg13g2_fill_1 FILLER_31_1380 ();
 sg13g2_decap_8 FILLER_31_1438 ();
 sg13g2_decap_8 FILLER_31_1445 ();
 sg13g2_decap_8 FILLER_31_1452 ();
 sg13g2_decap_8 FILLER_31_1459 ();
 sg13g2_decap_8 FILLER_31_1466 ();
 sg13g2_decap_8 FILLER_31_1473 ();
 sg13g2_fill_2 FILLER_31_1480 ();
 sg13g2_fill_1 FILLER_31_1482 ();
 sg13g2_fill_2 FILLER_31_1513 ();
 sg13g2_fill_1 FILLER_31_1515 ();
 sg13g2_decap_4 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1555 ();
 sg13g2_fill_2 FILLER_31_1562 ();
 sg13g2_fill_2 FILLER_31_1572 ();
 sg13g2_fill_2 FILLER_31_1693 ();
 sg13g2_fill_1 FILLER_31_1695 ();
 sg13g2_decap_8 FILLER_31_1709 ();
 sg13g2_fill_1 FILLER_31_1721 ();
 sg13g2_decap_8 FILLER_31_1726 ();
 sg13g2_fill_1 FILLER_31_1738 ();
 sg13g2_decap_4 FILLER_31_1743 ();
 sg13g2_fill_1 FILLER_31_1747 ();
 sg13g2_decap_4 FILLER_31_1757 ();
 sg13g2_fill_1 FILLER_31_1761 ();
 sg13g2_decap_8 FILLER_31_1767 ();
 sg13g2_decap_8 FILLER_31_1779 ();
 sg13g2_decap_4 FILLER_31_1786 ();
 sg13g2_fill_2 FILLER_31_1790 ();
 sg13g2_fill_2 FILLER_31_1801 ();
 sg13g2_fill_1 FILLER_31_1803 ();
 sg13g2_fill_2 FILLER_31_1808 ();
 sg13g2_fill_1 FILLER_31_1810 ();
 sg13g2_decap_8 FILLER_31_1819 ();
 sg13g2_decap_4 FILLER_31_1826 ();
 sg13g2_fill_2 FILLER_31_1850 ();
 sg13g2_fill_2 FILLER_31_1855 ();
 sg13g2_fill_1 FILLER_31_1857 ();
 sg13g2_decap_8 FILLER_31_1863 ();
 sg13g2_fill_2 FILLER_31_1870 ();
 sg13g2_fill_1 FILLER_31_1872 ();
 sg13g2_decap_8 FILLER_31_1877 ();
 sg13g2_decap_8 FILLER_31_1884 ();
 sg13g2_decap_4 FILLER_31_1891 ();
 sg13g2_fill_1 FILLER_31_1895 ();
 sg13g2_decap_8 FILLER_31_1901 ();
 sg13g2_decap_8 FILLER_31_1908 ();
 sg13g2_decap_4 FILLER_31_1915 ();
 sg13g2_fill_1 FILLER_31_1919 ();
 sg13g2_decap_4 FILLER_31_1951 ();
 sg13g2_fill_1 FILLER_31_1955 ();
 sg13g2_decap_8 FILLER_31_1974 ();
 sg13g2_fill_2 FILLER_31_1981 ();
 sg13g2_fill_1 FILLER_31_1983 ();
 sg13g2_decap_8 FILLER_31_2024 ();
 sg13g2_decap_8 FILLER_31_2031 ();
 sg13g2_decap_8 FILLER_31_2038 ();
 sg13g2_decap_8 FILLER_31_2045 ();
 sg13g2_decap_8 FILLER_31_2052 ();
 sg13g2_decap_8 FILLER_31_2059 ();
 sg13g2_decap_8 FILLER_31_2066 ();
 sg13g2_decap_8 FILLER_31_2073 ();
 sg13g2_decap_8 FILLER_31_2080 ();
 sg13g2_fill_1 FILLER_31_2087 ();
 sg13g2_decap_4 FILLER_31_2092 ();
 sg13g2_fill_1 FILLER_31_2122 ();
 sg13g2_fill_2 FILLER_31_2151 ();
 sg13g2_decap_4 FILLER_31_2158 ();
 sg13g2_fill_1 FILLER_31_2162 ();
 sg13g2_decap_4 FILLER_31_2167 ();
 sg13g2_fill_2 FILLER_31_2171 ();
 sg13g2_decap_8 FILLER_31_2198 ();
 sg13g2_decap_4 FILLER_31_2205 ();
 sg13g2_fill_1 FILLER_31_2209 ();
 sg13g2_decap_4 FILLER_31_2219 ();
 sg13g2_fill_2 FILLER_31_2223 ();
 sg13g2_decap_8 FILLER_31_2251 ();
 sg13g2_decap_8 FILLER_31_2258 ();
 sg13g2_decap_4 FILLER_31_2265 ();
 sg13g2_decap_4 FILLER_31_2295 ();
 sg13g2_fill_1 FILLER_31_2299 ();
 sg13g2_decap_8 FILLER_31_2309 ();
 sg13g2_fill_2 FILLER_31_2316 ();
 sg13g2_decap_8 FILLER_31_2401 ();
 sg13g2_decap_8 FILLER_31_2408 ();
 sg13g2_fill_2 FILLER_31_2415 ();
 sg13g2_fill_2 FILLER_31_2437 ();
 sg13g2_fill_1 FILLER_31_2453 ();
 sg13g2_fill_2 FILLER_31_2467 ();
 sg13g2_fill_2 FILLER_31_2477 ();
 sg13g2_fill_2 FILLER_31_2505 ();
 sg13g2_decap_8 FILLER_31_2517 ();
 sg13g2_fill_1 FILLER_31_2524 ();
 sg13g2_decap_4 FILLER_31_2529 ();
 sg13g2_decap_8 FILLER_31_2537 ();
 sg13g2_decap_8 FILLER_31_2544 ();
 sg13g2_decap_8 FILLER_31_2551 ();
 sg13g2_decap_8 FILLER_31_2558 ();
 sg13g2_decap_8 FILLER_31_2565 ();
 sg13g2_decap_8 FILLER_31_2572 ();
 sg13g2_decap_8 FILLER_31_2579 ();
 sg13g2_decap_8 FILLER_31_2586 ();
 sg13g2_decap_8 FILLER_31_2593 ();
 sg13g2_decap_8 FILLER_31_2600 ();
 sg13g2_decap_8 FILLER_31_2607 ();
 sg13g2_decap_8 FILLER_31_2614 ();
 sg13g2_decap_8 FILLER_31_2621 ();
 sg13g2_decap_8 FILLER_31_2628 ();
 sg13g2_decap_8 FILLER_31_2635 ();
 sg13g2_decap_8 FILLER_31_2642 ();
 sg13g2_decap_8 FILLER_31_2649 ();
 sg13g2_decap_8 FILLER_31_2656 ();
 sg13g2_decap_8 FILLER_31_2663 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_34 ();
 sg13g2_decap_8 FILLER_32_41 ();
 sg13g2_decap_8 FILLER_32_48 ();
 sg13g2_decap_4 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_59 ();
 sg13g2_decap_4 FILLER_32_87 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_4 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_decap_8 FILLER_32_288 ();
 sg13g2_decap_4 FILLER_32_295 ();
 sg13g2_fill_2 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_1 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_2 FILLER_32_429 ();
 sg13g2_fill_1 FILLER_32_431 ();
 sg13g2_decap_8 FILLER_32_437 ();
 sg13g2_fill_1 FILLER_32_444 ();
 sg13g2_decap_4 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_456 ();
 sg13g2_fill_2 FILLER_32_463 ();
 sg13g2_fill_2 FILLER_32_468 ();
 sg13g2_fill_2 FILLER_32_477 ();
 sg13g2_fill_2 FILLER_32_484 ();
 sg13g2_fill_1 FILLER_32_486 ();
 sg13g2_fill_2 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_fill_2 FILLER_32_530 ();
 sg13g2_decap_4 FILLER_32_584 ();
 sg13g2_fill_2 FILLER_32_597 ();
 sg13g2_fill_1 FILLER_32_599 ();
 sg13g2_decap_4 FILLER_32_612 ();
 sg13g2_fill_2 FILLER_32_616 ();
 sg13g2_fill_1 FILLER_32_626 ();
 sg13g2_decap_4 FILLER_32_635 ();
 sg13g2_fill_2 FILLER_32_649 ();
 sg13g2_fill_1 FILLER_32_651 ();
 sg13g2_decap_4 FILLER_32_662 ();
 sg13g2_decap_8 FILLER_32_670 ();
 sg13g2_decap_8 FILLER_32_684 ();
 sg13g2_decap_8 FILLER_32_691 ();
 sg13g2_fill_2 FILLER_32_698 ();
 sg13g2_fill_2 FILLER_32_710 ();
 sg13g2_fill_2 FILLER_32_749 ();
 sg13g2_fill_1 FILLER_32_751 ();
 sg13g2_fill_2 FILLER_32_784 ();
 sg13g2_fill_1 FILLER_32_792 ();
 sg13g2_fill_1 FILLER_32_797 ();
 sg13g2_fill_1 FILLER_32_824 ();
 sg13g2_fill_1 FILLER_32_877 ();
 sg13g2_decap_4 FILLER_32_925 ();
 sg13g2_decap_4 FILLER_32_934 ();
 sg13g2_fill_1 FILLER_32_943 ();
 sg13g2_decap_8 FILLER_32_970 ();
 sg13g2_fill_1 FILLER_32_977 ();
 sg13g2_fill_1 FILLER_32_1009 ();
 sg13g2_fill_1 FILLER_32_1016 ();
 sg13g2_fill_2 FILLER_32_1023 ();
 sg13g2_decap_8 FILLER_32_1037 ();
 sg13g2_decap_4 FILLER_32_1044 ();
 sg13g2_fill_2 FILLER_32_1048 ();
 sg13g2_fill_2 FILLER_32_1065 ();
 sg13g2_fill_1 FILLER_32_1072 ();
 sg13g2_decap_8 FILLER_32_1115 ();
 sg13g2_decap_8 FILLER_32_1122 ();
 sg13g2_decap_8 FILLER_32_1143 ();
 sg13g2_decap_4 FILLER_32_1150 ();
 sg13g2_fill_1 FILLER_32_1154 ();
 sg13g2_decap_4 FILLER_32_1160 ();
 sg13g2_fill_1 FILLER_32_1173 ();
 sg13g2_fill_1 FILLER_32_1203 ();
 sg13g2_decap_8 FILLER_32_1209 ();
 sg13g2_fill_2 FILLER_32_1216 ();
 sg13g2_fill_2 FILLER_32_1226 ();
 sg13g2_decap_4 FILLER_32_1254 ();
 sg13g2_fill_1 FILLER_32_1319 ();
 sg13g2_fill_1 FILLER_32_1340 ();
 sg13g2_fill_2 FILLER_32_1346 ();
 sg13g2_fill_1 FILLER_32_1348 ();
 sg13g2_fill_1 FILLER_32_1381 ();
 sg13g2_fill_1 FILLER_32_1389 ();
 sg13g2_fill_1 FILLER_32_1399 ();
 sg13g2_fill_1 FILLER_32_1422 ();
 sg13g2_fill_2 FILLER_32_1449 ();
 sg13g2_fill_1 FILLER_32_1451 ();
 sg13g2_decap_4 FILLER_32_1456 ();
 sg13g2_fill_1 FILLER_32_1465 ();
 sg13g2_fill_1 FILLER_32_1470 ();
 sg13g2_fill_1 FILLER_32_1475 ();
 sg13g2_fill_2 FILLER_32_1506 ();
 sg13g2_fill_1 FILLER_32_1513 ();
 sg13g2_decap_8 FILLER_32_1518 ();
 sg13g2_decap_4 FILLER_32_1525 ();
 sg13g2_fill_1 FILLER_32_1529 ();
 sg13g2_decap_8 FILLER_32_1535 ();
 sg13g2_decap_8 FILLER_32_1542 ();
 sg13g2_decap_8 FILLER_32_1549 ();
 sg13g2_fill_1 FILLER_32_1556 ();
 sg13g2_decap_8 FILLER_32_1561 ();
 sg13g2_fill_2 FILLER_32_1568 ();
 sg13g2_fill_1 FILLER_32_1581 ();
 sg13g2_decap_8 FILLER_32_1590 ();
 sg13g2_decap_8 FILLER_32_1597 ();
 sg13g2_decap_8 FILLER_32_1604 ();
 sg13g2_fill_1 FILLER_32_1615 ();
 sg13g2_fill_2 FILLER_32_1625 ();
 sg13g2_decap_8 FILLER_32_1631 ();
 sg13g2_decap_4 FILLER_32_1638 ();
 sg13g2_fill_2 FILLER_32_1651 ();
 sg13g2_fill_1 FILLER_32_1653 ();
 sg13g2_decap_8 FILLER_32_1660 ();
 sg13g2_decap_8 FILLER_32_1667 ();
 sg13g2_decap_4 FILLER_32_1674 ();
 sg13g2_fill_1 FILLER_32_1683 ();
 sg13g2_fill_1 FILLER_32_1688 ();
 sg13g2_decap_8 FILLER_32_1715 ();
 sg13g2_decap_8 FILLER_32_1722 ();
 sg13g2_decap_8 FILLER_32_1729 ();
 sg13g2_fill_1 FILLER_32_1736 ();
 sg13g2_decap_8 FILLER_32_1789 ();
 sg13g2_decap_8 FILLER_32_1796 ();
 sg13g2_decap_8 FILLER_32_1803 ();
 sg13g2_decap_8 FILLER_32_1810 ();
 sg13g2_decap_4 FILLER_32_1817 ();
 sg13g2_fill_1 FILLER_32_1821 ();
 sg13g2_fill_1 FILLER_32_1828 ();
 sg13g2_decap_8 FILLER_32_1894 ();
 sg13g2_decap_8 FILLER_32_1901 ();
 sg13g2_decap_8 FILLER_32_1908 ();
 sg13g2_decap_4 FILLER_32_1925 ();
 sg13g2_decap_4 FILLER_32_1939 ();
 sg13g2_fill_1 FILLER_32_1943 ();
 sg13g2_decap_4 FILLER_32_1948 ();
 sg13g2_fill_2 FILLER_32_1952 ();
 sg13g2_fill_2 FILLER_32_1958 ();
 sg13g2_fill_2 FILLER_32_1999 ();
 sg13g2_fill_1 FILLER_32_2001 ();
 sg13g2_fill_2 FILLER_32_2020 ();
 sg13g2_fill_1 FILLER_32_2022 ();
 sg13g2_decap_8 FILLER_32_2032 ();
 sg13g2_decap_8 FILLER_32_2039 ();
 sg13g2_decap_4 FILLER_32_2046 ();
 sg13g2_fill_1 FILLER_32_2050 ();
 sg13g2_decap_4 FILLER_32_2056 ();
 sg13g2_fill_1 FILLER_32_2060 ();
 sg13g2_decap_4 FILLER_32_2065 ();
 sg13g2_fill_2 FILLER_32_2069 ();
 sg13g2_decap_4 FILLER_32_2076 ();
 sg13g2_fill_1 FILLER_32_2080 ();
 sg13g2_fill_2 FILLER_32_2112 ();
 sg13g2_fill_1 FILLER_32_2127 ();
 sg13g2_decap_8 FILLER_32_2166 ();
 sg13g2_decap_8 FILLER_32_2173 ();
 sg13g2_decap_8 FILLER_32_2180 ();
 sg13g2_decap_8 FILLER_32_2224 ();
 sg13g2_decap_8 FILLER_32_2231 ();
 sg13g2_decap_8 FILLER_32_2238 ();
 sg13g2_decap_4 FILLER_32_2245 ();
 sg13g2_fill_2 FILLER_32_2320 ();
 sg13g2_fill_1 FILLER_32_2326 ();
 sg13g2_decap_8 FILLER_32_2340 ();
 sg13g2_fill_1 FILLER_32_2347 ();
 sg13g2_decap_8 FILLER_32_2406 ();
 sg13g2_decap_8 FILLER_32_2413 ();
 sg13g2_decap_4 FILLER_32_2420 ();
 sg13g2_fill_2 FILLER_32_2424 ();
 sg13g2_decap_4 FILLER_32_2429 ();
 sg13g2_fill_2 FILLER_32_2433 ();
 sg13g2_fill_2 FILLER_32_2478 ();
 sg13g2_fill_2 FILLER_32_2488 ();
 sg13g2_fill_1 FILLER_32_2490 ();
 sg13g2_decap_4 FILLER_32_2504 ();
 sg13g2_decap_8 FILLER_32_2522 ();
 sg13g2_decap_8 FILLER_32_2529 ();
 sg13g2_fill_2 FILLER_32_2536 ();
 sg13g2_decap_8 FILLER_32_2568 ();
 sg13g2_decap_8 FILLER_32_2575 ();
 sg13g2_decap_8 FILLER_32_2582 ();
 sg13g2_decap_8 FILLER_32_2589 ();
 sg13g2_decap_8 FILLER_32_2596 ();
 sg13g2_decap_8 FILLER_32_2603 ();
 sg13g2_decap_8 FILLER_32_2610 ();
 sg13g2_decap_8 FILLER_32_2617 ();
 sg13g2_decap_8 FILLER_32_2624 ();
 sg13g2_decap_8 FILLER_32_2631 ();
 sg13g2_decap_8 FILLER_32_2638 ();
 sg13g2_decap_8 FILLER_32_2645 ();
 sg13g2_decap_8 FILLER_32_2652 ();
 sg13g2_decap_8 FILLER_32_2659 ();
 sg13g2_decap_4 FILLER_32_2666 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_16 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_decap_4 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_decap_4 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_decap_4 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_decap_4 FILLER_33_332 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_4 FILLER_33_409 ();
 sg13g2_fill_1 FILLER_33_413 ();
 sg13g2_decap_4 FILLER_33_440 ();
 sg13g2_fill_1 FILLER_33_461 ();
 sg13g2_fill_2 FILLER_33_467 ();
 sg13g2_fill_2 FILLER_33_474 ();
 sg13g2_fill_1 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_482 ();
 sg13g2_fill_2 FILLER_33_489 ();
 sg13g2_fill_1 FILLER_33_491 ();
 sg13g2_fill_2 FILLER_33_497 ();
 sg13g2_decap_4 FILLER_33_514 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_fill_2 FILLER_33_537 ();
 sg13g2_fill_1 FILLER_33_547 ();
 sg13g2_fill_1 FILLER_33_555 ();
 sg13g2_fill_1 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_569 ();
 sg13g2_fill_1 FILLER_33_571 ();
 sg13g2_fill_2 FILLER_33_585 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_decap_4 FILLER_33_607 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_4 FILLER_33_623 ();
 sg13g2_fill_2 FILLER_33_663 ();
 sg13g2_fill_1 FILLER_33_670 ();
 sg13g2_decap_8 FILLER_33_708 ();
 sg13g2_decap_8 FILLER_33_715 ();
 sg13g2_decap_8 FILLER_33_722 ();
 sg13g2_fill_2 FILLER_33_729 ();
 sg13g2_decap_4 FILLER_33_735 ();
 sg13g2_fill_2 FILLER_33_739 ();
 sg13g2_decap_4 FILLER_33_745 ();
 sg13g2_fill_1 FILLER_33_749 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_4 FILLER_33_800 ();
 sg13g2_fill_2 FILLER_33_804 ();
 sg13g2_decap_4 FILLER_33_842 ();
 sg13g2_fill_2 FILLER_33_854 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_fill_1 FILLER_33_862 ();
 sg13g2_fill_2 FILLER_33_867 ();
 sg13g2_fill_1 FILLER_33_869 ();
 sg13g2_fill_1 FILLER_33_896 ();
 sg13g2_fill_1 FILLER_33_903 ();
 sg13g2_decap_4 FILLER_33_924 ();
 sg13g2_fill_1 FILLER_33_928 ();
 sg13g2_decap_8 FILLER_33_933 ();
 sg13g2_decap_8 FILLER_33_940 ();
 sg13g2_decap_8 FILLER_33_947 ();
 sg13g2_fill_1 FILLER_33_954 ();
 sg13g2_fill_2 FILLER_33_960 ();
 sg13g2_fill_1 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1006 ();
 sg13g2_decap_4 FILLER_33_1013 ();
 sg13g2_fill_2 FILLER_33_1017 ();
 sg13g2_fill_2 FILLER_33_1051 ();
 sg13g2_fill_1 FILLER_33_1059 ();
 sg13g2_fill_2 FILLER_33_1086 ();
 sg13g2_fill_2 FILLER_33_1093 ();
 sg13g2_decap_8 FILLER_33_1121 ();
 sg13g2_fill_1 FILLER_33_1128 ();
 sg13g2_fill_2 FILLER_33_1138 ();
 sg13g2_fill_2 FILLER_33_1188 ();
 sg13g2_decap_4 FILLER_33_1226 ();
 sg13g2_decap_4 FILLER_33_1236 ();
 sg13g2_fill_2 FILLER_33_1266 ();
 sg13g2_decap_4 FILLER_33_1272 ();
 sg13g2_decap_8 FILLER_33_1282 ();
 sg13g2_decap_4 FILLER_33_1289 ();
 sg13g2_fill_1 FILLER_33_1299 ();
 sg13g2_fill_1 FILLER_33_1366 ();
 sg13g2_fill_1 FILLER_33_1375 ();
 sg13g2_fill_2 FILLER_33_1399 ();
 sg13g2_decap_8 FILLER_33_1439 ();
 sg13g2_decap_8 FILLER_33_1446 ();
 sg13g2_fill_1 FILLER_33_1453 ();
 sg13g2_decap_4 FILLER_33_1489 ();
 sg13g2_fill_1 FILLER_33_1493 ();
 sg13g2_decap_8 FILLER_33_1533 ();
 sg13g2_decap_8 FILLER_33_1540 ();
 sg13g2_fill_2 FILLER_33_1594 ();
 sg13g2_fill_1 FILLER_33_1596 ();
 sg13g2_decap_8 FILLER_33_1629 ();
 sg13g2_decap_8 FILLER_33_1636 ();
 sg13g2_decap_8 FILLER_33_1643 ();
 sg13g2_fill_2 FILLER_33_1650 ();
 sg13g2_decap_8 FILLER_33_1656 ();
 sg13g2_decap_8 FILLER_33_1663 ();
 sg13g2_decap_4 FILLER_33_1670 ();
 sg13g2_fill_2 FILLER_33_1674 ();
 sg13g2_fill_1 FILLER_33_1680 ();
 sg13g2_decap_8 FILLER_33_1686 ();
 sg13g2_fill_2 FILLER_33_1693 ();
 sg13g2_fill_1 FILLER_33_1695 ();
 sg13g2_decap_8 FILLER_33_1715 ();
 sg13g2_decap_8 FILLER_33_1722 ();
 sg13g2_decap_8 FILLER_33_1729 ();
 sg13g2_decap_8 FILLER_33_1741 ();
 sg13g2_decap_8 FILLER_33_1748 ();
 sg13g2_decap_8 FILLER_33_1759 ();
 sg13g2_decap_8 FILLER_33_1766 ();
 sg13g2_decap_8 FILLER_33_1773 ();
 sg13g2_decap_8 FILLER_33_1810 ();
 sg13g2_decap_8 FILLER_33_1817 ();
 sg13g2_fill_1 FILLER_33_1824 ();
 sg13g2_fill_1 FILLER_33_1834 ();
 sg13g2_fill_1 FILLER_33_1861 ();
 sg13g2_fill_1 FILLER_33_1879 ();
 sg13g2_decap_8 FILLER_33_1884 ();
 sg13g2_decap_8 FILLER_33_1896 ();
 sg13g2_fill_2 FILLER_33_1903 ();
 sg13g2_fill_1 FILLER_33_1905 ();
 sg13g2_decap_8 FILLER_33_1937 ();
 sg13g2_decap_4 FILLER_33_1944 ();
 sg13g2_fill_1 FILLER_33_1958 ();
 sg13g2_decap_4 FILLER_33_1965 ();
 sg13g2_fill_1 FILLER_33_1969 ();
 sg13g2_fill_1 FILLER_33_1990 ();
 sg13g2_decap_4 FILLER_33_1995 ();
 sg13g2_decap_8 FILLER_33_2029 ();
 sg13g2_fill_2 FILLER_33_2036 ();
 sg13g2_decap_4 FILLER_33_2043 ();
 sg13g2_fill_1 FILLER_33_2047 ();
 sg13g2_fill_2 FILLER_33_2052 ();
 sg13g2_fill_1 FILLER_33_2054 ();
 sg13g2_fill_2 FILLER_33_2064 ();
 sg13g2_fill_1 FILLER_33_2066 ();
 sg13g2_fill_1 FILLER_33_2102 ();
 sg13g2_fill_2 FILLER_33_2109 ();
 sg13g2_fill_2 FILLER_33_2143 ();
 sg13g2_fill_2 FILLER_33_2153 ();
 sg13g2_decap_8 FILLER_33_2164 ();
 sg13g2_fill_1 FILLER_33_2171 ();
 sg13g2_decap_8 FILLER_33_2204 ();
 sg13g2_decap_8 FILLER_33_2211 ();
 sg13g2_decap_8 FILLER_33_2218 ();
 sg13g2_decap_4 FILLER_33_2225 ();
 sg13g2_fill_2 FILLER_33_2229 ();
 sg13g2_decap_4 FILLER_33_2236 ();
 sg13g2_fill_2 FILLER_33_2240 ();
 sg13g2_fill_2 FILLER_33_2246 ();
 sg13g2_fill_1 FILLER_33_2248 ();
 sg13g2_decap_4 FILLER_33_2265 ();
 sg13g2_fill_1 FILLER_33_2269 ();
 sg13g2_fill_2 FILLER_33_2275 ();
 sg13g2_fill_1 FILLER_33_2277 ();
 sg13g2_decap_8 FILLER_33_2301 ();
 sg13g2_decap_8 FILLER_33_2334 ();
 sg13g2_decap_8 FILLER_33_2341 ();
 sg13g2_decap_4 FILLER_33_2348 ();
 sg13g2_fill_1 FILLER_33_2352 ();
 sg13g2_fill_1 FILLER_33_2398 ();
 sg13g2_decap_4 FILLER_33_2425 ();
 sg13g2_fill_2 FILLER_33_2463 ();
 sg13g2_decap_8 FILLER_33_2508 ();
 sg13g2_decap_4 FILLER_33_2515 ();
 sg13g2_decap_8 FILLER_33_2553 ();
 sg13g2_decap_8 FILLER_33_2560 ();
 sg13g2_decap_8 FILLER_33_2567 ();
 sg13g2_decap_8 FILLER_33_2574 ();
 sg13g2_decap_8 FILLER_33_2581 ();
 sg13g2_decap_8 FILLER_33_2588 ();
 sg13g2_decap_8 FILLER_33_2595 ();
 sg13g2_decap_8 FILLER_33_2602 ();
 sg13g2_decap_8 FILLER_33_2609 ();
 sg13g2_decap_8 FILLER_33_2616 ();
 sg13g2_decap_8 FILLER_33_2623 ();
 sg13g2_decap_8 FILLER_33_2630 ();
 sg13g2_decap_8 FILLER_33_2637 ();
 sg13g2_decap_8 FILLER_33_2644 ();
 sg13g2_decap_8 FILLER_33_2651 ();
 sg13g2_decap_8 FILLER_33_2658 ();
 sg13g2_decap_4 FILLER_33_2665 ();
 sg13g2_fill_1 FILLER_33_2669 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_19 ();
 sg13g2_decap_4 FILLER_34_34 ();
 sg13g2_decap_4 FILLER_34_68 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_decap_8 FILLER_34_108 ();
 sg13g2_decap_8 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_271 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_344 ();
 sg13g2_decap_4 FILLER_34_365 ();
 sg13g2_decap_4 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_fill_2 FILLER_34_430 ();
 sg13g2_fill_1 FILLER_34_432 ();
 sg13g2_decap_8 FILLER_34_440 ();
 sg13g2_decap_8 FILLER_34_447 ();
 sg13g2_decap_8 FILLER_34_454 ();
 sg13g2_decap_8 FILLER_34_461 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_fill_1 FILLER_34_475 ();
 sg13g2_decap_8 FILLER_34_480 ();
 sg13g2_decap_4 FILLER_34_487 ();
 sg13g2_decap_4 FILLER_34_499 ();
 sg13g2_fill_1 FILLER_34_512 ();
 sg13g2_fill_1 FILLER_34_539 ();
 sg13g2_fill_1 FILLER_34_552 ();
 sg13g2_fill_1 FILLER_34_561 ();
 sg13g2_fill_2 FILLER_34_566 ();
 sg13g2_fill_1 FILLER_34_568 ();
 sg13g2_fill_1 FILLER_34_572 ();
 sg13g2_fill_1 FILLER_34_601 ();
 sg13g2_fill_2 FILLER_34_607 ();
 sg13g2_decap_8 FILLER_34_612 ();
 sg13g2_decap_8 FILLER_34_619 ();
 sg13g2_decap_8 FILLER_34_626 ();
 sg13g2_decap_8 FILLER_34_633 ();
 sg13g2_fill_2 FILLER_34_640 ();
 sg13g2_fill_1 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_687 ();
 sg13g2_decap_8 FILLER_34_694 ();
 sg13g2_decap_8 FILLER_34_701 ();
 sg13g2_decap_8 FILLER_34_708 ();
 sg13g2_decap_8 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_decap_4 FILLER_34_729 ();
 sg13g2_fill_1 FILLER_34_755 ();
 sg13g2_fill_2 FILLER_34_761 ();
 sg13g2_fill_1 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_fill_2 FILLER_34_817 ();
 sg13g2_fill_1 FILLER_34_819 ();
 sg13g2_decap_4 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_fill_2 FILLER_34_858 ();
 sg13g2_fill_1 FILLER_34_860 ();
 sg13g2_fill_1 FILLER_34_870 ();
 sg13g2_fill_2 FILLER_34_929 ();
 sg13g2_fill_2 FILLER_34_971 ();
 sg13g2_decap_8 FILLER_34_1018 ();
 sg13g2_decap_4 FILLER_34_1025 ();
 sg13g2_fill_1 FILLER_34_1029 ();
 sg13g2_fill_2 FILLER_34_1034 ();
 sg13g2_fill_1 FILLER_34_1036 ();
 sg13g2_fill_2 FILLER_34_1041 ();
 sg13g2_fill_2 FILLER_34_1048 ();
 sg13g2_fill_2 FILLER_34_1054 ();
 sg13g2_fill_1 FILLER_34_1056 ();
 sg13g2_fill_1 FILLER_34_1062 ();
 sg13g2_decap_8 FILLER_34_1067 ();
 sg13g2_decap_8 FILLER_34_1078 ();
 sg13g2_decap_8 FILLER_34_1085 ();
 sg13g2_fill_1 FILLER_34_1101 ();
 sg13g2_fill_1 FILLER_34_1108 ();
 sg13g2_decap_4 FILLER_34_1156 ();
 sg13g2_fill_1 FILLER_34_1163 ();
 sg13g2_decap_4 FILLER_34_1170 ();
 sg13g2_fill_1 FILLER_34_1174 ();
 sg13g2_fill_2 FILLER_34_1180 ();
 sg13g2_fill_1 FILLER_34_1182 ();
 sg13g2_decap_4 FILLER_34_1187 ();
 sg13g2_fill_1 FILLER_34_1191 ();
 sg13g2_decap_4 FILLER_34_1202 ();
 sg13g2_decap_8 FILLER_34_1219 ();
 sg13g2_fill_2 FILLER_34_1226 ();
 sg13g2_fill_1 FILLER_34_1228 ();
 sg13g2_fill_1 FILLER_34_1237 ();
 sg13g2_decap_8 FILLER_34_1247 ();
 sg13g2_decap_8 FILLER_34_1254 ();
 sg13g2_decap_8 FILLER_34_1261 ();
 sg13g2_decap_8 FILLER_34_1268 ();
 sg13g2_fill_1 FILLER_34_1316 ();
 sg13g2_decap_8 FILLER_34_1334 ();
 sg13g2_fill_2 FILLER_34_1341 ();
 sg13g2_decap_8 FILLER_34_1419 ();
 sg13g2_decap_8 FILLER_34_1426 ();
 sg13g2_decap_8 FILLER_34_1433 ();
 sg13g2_decap_8 FILLER_34_1440 ();
 sg13g2_decap_4 FILLER_34_1447 ();
 sg13g2_fill_2 FILLER_34_1492 ();
 sg13g2_decap_8 FILLER_34_1499 ();
 sg13g2_fill_2 FILLER_34_1510 ();
 sg13g2_fill_1 FILLER_34_1515 ();
 sg13g2_fill_1 FILLER_34_1522 ();
 sg13g2_decap_8 FILLER_34_1527 ();
 sg13g2_decap_8 FILLER_34_1534 ();
 sg13g2_fill_1 FILLER_34_1546 ();
 sg13g2_decap_8 FILLER_34_1552 ();
 sg13g2_fill_1 FILLER_34_1559 ();
 sg13g2_fill_1 FILLER_34_1577 ();
 sg13g2_fill_1 FILLER_34_1584 ();
 sg13g2_fill_1 FILLER_34_1591 ();
 sg13g2_fill_2 FILLER_34_1629 ();
 sg13g2_fill_1 FILLER_34_1631 ();
 sg13g2_fill_2 FILLER_34_1638 ();
 sg13g2_fill_1 FILLER_34_1640 ();
 sg13g2_fill_2 FILLER_34_1652 ();
 sg13g2_fill_1 FILLER_34_1654 ();
 sg13g2_decap_8 FILLER_34_1715 ();
 sg13g2_decap_8 FILLER_34_1722 ();
 sg13g2_decap_4 FILLER_34_1768 ();
 sg13g2_fill_2 FILLER_34_1772 ();
 sg13g2_fill_1 FILLER_34_1779 ();
 sg13g2_fill_2 FILLER_34_1806 ();
 sg13g2_fill_1 FILLER_34_1834 ();
 sg13g2_decap_8 FILLER_34_1843 ();
 sg13g2_fill_2 FILLER_34_1850 ();
 sg13g2_fill_1 FILLER_34_1852 ();
 sg13g2_fill_2 FILLER_34_1894 ();
 sg13g2_fill_1 FILLER_34_1896 ();
 sg13g2_decap_8 FILLER_34_1927 ();
 sg13g2_fill_1 FILLER_34_1934 ();
 sg13g2_decap_4 FILLER_34_1940 ();
 sg13g2_fill_2 FILLER_34_1944 ();
 sg13g2_decap_4 FILLER_34_1950 ();
 sg13g2_decap_8 FILLER_34_1958 ();
 sg13g2_fill_2 FILLER_34_1969 ();
 sg13g2_decap_8 FILLER_34_1984 ();
 sg13g2_decap_4 FILLER_34_1991 ();
 sg13g2_fill_1 FILLER_34_1995 ();
 sg13g2_fill_2 FILLER_34_2022 ();
 sg13g2_fill_1 FILLER_34_2024 ();
 sg13g2_decap_4 FILLER_34_2038 ();
 sg13g2_fill_2 FILLER_34_2068 ();
 sg13g2_fill_1 FILLER_34_2070 ();
 sg13g2_fill_1 FILLER_34_2076 ();
 sg13g2_fill_2 FILLER_34_2086 ();
 sg13g2_fill_1 FILLER_34_2117 ();
 sg13g2_decap_8 FILLER_34_2152 ();
 sg13g2_decap_4 FILLER_34_2159 ();
 sg13g2_fill_1 FILLER_34_2163 ();
 sg13g2_fill_1 FILLER_34_2169 ();
 sg13g2_decap_8 FILLER_34_2222 ();
 sg13g2_decap_8 FILLER_34_2229 ();
 sg13g2_fill_2 FILLER_34_2236 ();
 sg13g2_fill_1 FILLER_34_2238 ();
 sg13g2_decap_8 FILLER_34_2270 ();
 sg13g2_decap_4 FILLER_34_2277 ();
 sg13g2_fill_2 FILLER_34_2281 ();
 sg13g2_fill_1 FILLER_34_2291 ();
 sg13g2_fill_2 FILLER_34_2307 ();
 sg13g2_fill_1 FILLER_34_2327 ();
 sg13g2_fill_2 FILLER_34_2354 ();
 sg13g2_fill_1 FILLER_34_2390 ();
 sg13g2_decap_8 FILLER_34_2411 ();
 sg13g2_decap_4 FILLER_34_2418 ();
 sg13g2_fill_1 FILLER_34_2422 ();
 sg13g2_fill_2 FILLER_34_2469 ();
 sg13g2_fill_1 FILLER_34_2471 ();
 sg13g2_decap_8 FILLER_34_2476 ();
 sg13g2_decap_4 FILLER_34_2483 ();
 sg13g2_fill_1 FILLER_34_2487 ();
 sg13g2_fill_1 FILLER_34_2524 ();
 sg13g2_decap_8 FILLER_34_2551 ();
 sg13g2_decap_8 FILLER_34_2558 ();
 sg13g2_decap_8 FILLER_34_2565 ();
 sg13g2_decap_8 FILLER_34_2572 ();
 sg13g2_decap_8 FILLER_34_2579 ();
 sg13g2_decap_8 FILLER_34_2586 ();
 sg13g2_decap_8 FILLER_34_2593 ();
 sg13g2_decap_8 FILLER_34_2600 ();
 sg13g2_decap_8 FILLER_34_2607 ();
 sg13g2_decap_8 FILLER_34_2614 ();
 sg13g2_decap_8 FILLER_34_2621 ();
 sg13g2_decap_8 FILLER_34_2628 ();
 sg13g2_decap_8 FILLER_34_2635 ();
 sg13g2_decap_8 FILLER_34_2642 ();
 sg13g2_decap_8 FILLER_34_2649 ();
 sg13g2_decap_8 FILLER_34_2656 ();
 sg13g2_decap_8 FILLER_34_2663 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_16 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_decap_4 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_decap_8 FILLER_35_78 ();
 sg13g2_fill_2 FILLER_35_89 ();
 sg13g2_decap_8 FILLER_35_117 ();
 sg13g2_decap_4 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_131 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_decap_8 FILLER_35_157 ();
 sg13g2_decap_8 FILLER_35_164 ();
 sg13g2_decap_8 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_4 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_decap_8 FILLER_35_234 ();
 sg13g2_decap_8 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_35_415 ();
 sg13g2_fill_1 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_440 ();
 sg13g2_decap_8 FILLER_35_474 ();
 sg13g2_fill_2 FILLER_35_481 ();
 sg13g2_fill_1 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_decap_8 FILLER_35_540 ();
 sg13g2_decap_8 FILLER_35_547 ();
 sg13g2_decap_8 FILLER_35_554 ();
 sg13g2_decap_8 FILLER_35_561 ();
 sg13g2_decap_4 FILLER_35_568 ();
 sg13g2_decap_4 FILLER_35_626 ();
 sg13g2_fill_1 FILLER_35_630 ();
 sg13g2_fill_2 FILLER_35_641 ();
 sg13g2_fill_1 FILLER_35_651 ();
 sg13g2_decap_4 FILLER_35_667 ();
 sg13g2_fill_2 FILLER_35_671 ();
 sg13g2_fill_1 FILLER_35_678 ();
 sg13g2_decap_8 FILLER_35_689 ();
 sg13g2_fill_2 FILLER_35_726 ();
 sg13g2_fill_2 FILLER_35_754 ();
 sg13g2_fill_2 FILLER_35_782 ();
 sg13g2_fill_1 FILLER_35_784 ();
 sg13g2_fill_2 FILLER_35_811 ();
 sg13g2_fill_1 FILLER_35_813 ();
 sg13g2_decap_4 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_fill_2 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_fill_1 FILLER_35_868 ();
 sg13g2_fill_2 FILLER_35_879 ();
 sg13g2_decap_8 FILLER_35_885 ();
 sg13g2_decap_4 FILLER_35_892 ();
 sg13g2_fill_1 FILLER_35_896 ();
 sg13g2_decap_4 FILLER_35_912 ();
 sg13g2_fill_2 FILLER_35_916 ();
 sg13g2_fill_1 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_929 ();
 sg13g2_fill_1 FILLER_35_936 ();
 sg13g2_fill_1 FILLER_35_941 ();
 sg13g2_fill_2 FILLER_35_980 ();
 sg13g2_fill_1 FILLER_35_982 ();
 sg13g2_fill_1 FILLER_35_988 ();
 sg13g2_decap_4 FILLER_35_1001 ();
 sg13g2_fill_1 FILLER_35_1005 ();
 sg13g2_decap_4 FILLER_35_1012 ();
 sg13g2_fill_2 FILLER_35_1016 ();
 sg13g2_fill_2 FILLER_35_1029 ();
 sg13g2_decap_8 FILLER_35_1037 ();
 sg13g2_decap_4 FILLER_35_1044 ();
 sg13g2_decap_8 FILLER_35_1053 ();
 sg13g2_decap_8 FILLER_35_1064 ();
 sg13g2_decap_8 FILLER_35_1071 ();
 sg13g2_decap_8 FILLER_35_1078 ();
 sg13g2_decap_8 FILLER_35_1085 ();
 sg13g2_fill_1 FILLER_35_1096 ();
 sg13g2_fill_1 FILLER_35_1103 ();
 sg13g2_fill_1 FILLER_35_1119 ();
 sg13g2_fill_2 FILLER_35_1129 ();
 sg13g2_fill_2 FILLER_35_1134 ();
 sg13g2_fill_2 FILLER_35_1148 ();
 sg13g2_decap_4 FILLER_35_1155 ();
 sg13g2_fill_1 FILLER_35_1159 ();
 sg13g2_decap_8 FILLER_35_1164 ();
 sg13g2_fill_1 FILLER_35_1171 ();
 sg13g2_fill_2 FILLER_35_1198 ();
 sg13g2_fill_1 FILLER_35_1200 ();
 sg13g2_fill_1 FILLER_35_1207 ();
 sg13g2_fill_2 FILLER_35_1212 ();
 sg13g2_fill_1 FILLER_35_1214 ();
 sg13g2_fill_2 FILLER_35_1225 ();
 sg13g2_fill_1 FILLER_35_1236 ();
 sg13g2_fill_2 FILLER_35_1242 ();
 sg13g2_fill_1 FILLER_35_1250 ();
 sg13g2_decap_8 FILLER_35_1259 ();
 sg13g2_decap_8 FILLER_35_1266 ();
 sg13g2_decap_8 FILLER_35_1273 ();
 sg13g2_decap_8 FILLER_35_1280 ();
 sg13g2_decap_4 FILLER_35_1287 ();
 sg13g2_fill_2 FILLER_35_1291 ();
 sg13g2_fill_2 FILLER_35_1300 ();
 sg13g2_fill_1 FILLER_35_1311 ();
 sg13g2_fill_1 FILLER_35_1315 ();
 sg13g2_fill_2 FILLER_35_1320 ();
 sg13g2_fill_1 FILLER_35_1325 ();
 sg13g2_decap_8 FILLER_35_1336 ();
 sg13g2_fill_2 FILLER_35_1343 ();
 sg13g2_decap_4 FILLER_35_1393 ();
 sg13g2_fill_2 FILLER_35_1397 ();
 sg13g2_decap_8 FILLER_35_1402 ();
 sg13g2_fill_1 FILLER_35_1409 ();
 sg13g2_decap_4 FILLER_35_1430 ();
 sg13g2_decap_4 FILLER_35_1470 ();
 sg13g2_decap_8 FILLER_35_1479 ();
 sg13g2_decap_8 FILLER_35_1486 ();
 sg13g2_decap_8 FILLER_35_1493 ();
 sg13g2_fill_2 FILLER_35_1500 ();
 sg13g2_fill_1 FILLER_35_1502 ();
 sg13g2_fill_2 FILLER_35_1545 ();
 sg13g2_decap_8 FILLER_35_1583 ();
 sg13g2_decap_8 FILLER_35_1590 ();
 sg13g2_fill_1 FILLER_35_1632 ();
 sg13g2_decap_8 FILLER_35_1659 ();
 sg13g2_decap_8 FILLER_35_1666 ();
 sg13g2_decap_8 FILLER_35_1673 ();
 sg13g2_fill_2 FILLER_35_1680 ();
 sg13g2_fill_1 FILLER_35_1682 ();
 sg13g2_fill_1 FILLER_35_1692 ();
 sg13g2_fill_1 FILLER_35_1698 ();
 sg13g2_fill_2 FILLER_35_1703 ();
 sg13g2_fill_2 FILLER_35_1793 ();
 sg13g2_fill_2 FILLER_35_1803 ();
 sg13g2_fill_2 FILLER_35_1826 ();
 sg13g2_fill_1 FILLER_35_1828 ();
 sg13g2_decap_8 FILLER_35_1856 ();
 sg13g2_decap_8 FILLER_35_1863 ();
 sg13g2_fill_1 FILLER_35_1913 ();
 sg13g2_fill_2 FILLER_35_1923 ();
 sg13g2_fill_1 FILLER_35_1925 ();
 sg13g2_fill_2 FILLER_35_1956 ();
 sg13g2_fill_1 FILLER_35_1958 ();
 sg13g2_decap_8 FILLER_35_1994 ();
 sg13g2_fill_1 FILLER_35_2001 ();
 sg13g2_decap_8 FILLER_35_2011 ();
 sg13g2_fill_2 FILLER_35_2018 ();
 sg13g2_fill_1 FILLER_35_2069 ();
 sg13g2_fill_1 FILLER_35_2075 ();
 sg13g2_fill_1 FILLER_35_2081 ();
 sg13g2_fill_2 FILLER_35_2087 ();
 sg13g2_fill_1 FILLER_35_2089 ();
 sg13g2_decap_4 FILLER_35_2093 ();
 sg13g2_fill_1 FILLER_35_2109 ();
 sg13g2_fill_2 FILLER_35_2157 ();
 sg13g2_fill_1 FILLER_35_2182 ();
 sg13g2_fill_1 FILLER_35_2205 ();
 sg13g2_decap_4 FILLER_35_2216 ();
 sg13g2_fill_2 FILLER_35_2220 ();
 sg13g2_fill_2 FILLER_35_2227 ();
 sg13g2_fill_1 FILLER_35_2229 ();
 sg13g2_decap_8 FILLER_35_2234 ();
 sg13g2_decap_8 FILLER_35_2250 ();
 sg13g2_decap_8 FILLER_35_2257 ();
 sg13g2_fill_1 FILLER_35_2264 ();
 sg13g2_decap_8 FILLER_35_2269 ();
 sg13g2_decap_8 FILLER_35_2276 ();
 sg13g2_decap_4 FILLER_35_2283 ();
 sg13g2_decap_8 FILLER_35_2310 ();
 sg13g2_fill_1 FILLER_35_2317 ();
 sg13g2_decap_8 FILLER_35_2344 ();
 sg13g2_fill_2 FILLER_35_2351 ();
 sg13g2_fill_1 FILLER_35_2353 ();
 sg13g2_fill_2 FILLER_35_2360 ();
 sg13g2_fill_1 FILLER_35_2365 ();
 sg13g2_fill_1 FILLER_35_2369 ();
 sg13g2_fill_2 FILLER_35_2384 ();
 sg13g2_fill_1 FILLER_35_2389 ();
 sg13g2_fill_2 FILLER_35_2423 ();
 sg13g2_fill_1 FILLER_35_2425 ();
 sg13g2_fill_1 FILLER_35_2462 ();
 sg13g2_fill_1 FILLER_35_2489 ();
 sg13g2_decap_8 FILLER_35_2503 ();
 sg13g2_decap_4 FILLER_35_2510 ();
 sg13g2_fill_2 FILLER_35_2524 ();
 sg13g2_fill_2 FILLER_35_2534 ();
 sg13g2_fill_1 FILLER_35_2536 ();
 sg13g2_decap_8 FILLER_35_2541 ();
 sg13g2_decap_8 FILLER_35_2548 ();
 sg13g2_decap_8 FILLER_35_2555 ();
 sg13g2_decap_8 FILLER_35_2562 ();
 sg13g2_decap_8 FILLER_35_2569 ();
 sg13g2_decap_8 FILLER_35_2576 ();
 sg13g2_decap_8 FILLER_35_2583 ();
 sg13g2_decap_8 FILLER_35_2590 ();
 sg13g2_decap_8 FILLER_35_2597 ();
 sg13g2_decap_8 FILLER_35_2604 ();
 sg13g2_decap_8 FILLER_35_2611 ();
 sg13g2_decap_8 FILLER_35_2618 ();
 sg13g2_decap_8 FILLER_35_2625 ();
 sg13g2_decap_8 FILLER_35_2632 ();
 sg13g2_decap_8 FILLER_35_2639 ();
 sg13g2_decap_8 FILLER_35_2646 ();
 sg13g2_decap_8 FILLER_35_2653 ();
 sg13g2_decap_8 FILLER_35_2660 ();
 sg13g2_fill_2 FILLER_35_2667 ();
 sg13g2_fill_1 FILLER_35_2669 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_52 ();
 sg13g2_fill_2 FILLER_36_59 ();
 sg13g2_decap_4 FILLER_36_74 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_93 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_decap_4 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_decap_4 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_decap_4 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_decap_4 FILLER_36_349 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_decap_4 FILLER_36_431 ();
 sg13g2_fill_2 FILLER_36_435 ();
 sg13g2_fill_2 FILLER_36_477 ();
 sg13g2_fill_1 FILLER_36_479 ();
 sg13g2_decap_8 FILLER_36_531 ();
 sg13g2_fill_2 FILLER_36_538 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_fill_1 FILLER_36_607 ();
 sg13g2_fill_2 FILLER_36_613 ();
 sg13g2_fill_1 FILLER_36_615 ();
 sg13g2_fill_1 FILLER_36_646 ();
 sg13g2_fill_1 FILLER_36_655 ();
 sg13g2_decap_4 FILLER_36_691 ();
 sg13g2_fill_2 FILLER_36_726 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_fill_2 FILLER_36_764 ();
 sg13g2_fill_1 FILLER_36_766 ();
 sg13g2_fill_2 FILLER_36_771 ();
 sg13g2_fill_1 FILLER_36_773 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_fill_1 FILLER_36_791 ();
 sg13g2_decap_4 FILLER_36_810 ();
 sg13g2_decap_4 FILLER_36_823 ();
 sg13g2_fill_1 FILLER_36_827 ();
 sg13g2_decap_8 FILLER_36_863 ();
 sg13g2_decap_8 FILLER_36_870 ();
 sg13g2_decap_4 FILLER_36_877 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_decap_4 FILLER_36_893 ();
 sg13g2_fill_2 FILLER_36_897 ();
 sg13g2_decap_8 FILLER_36_916 ();
 sg13g2_decap_4 FILLER_36_923 ();
 sg13g2_fill_1 FILLER_36_927 ();
 sg13g2_fill_2 FILLER_36_933 ();
 sg13g2_fill_2 FILLER_36_951 ();
 sg13g2_fill_1 FILLER_36_953 ();
 sg13g2_fill_1 FILLER_36_960 ();
 sg13g2_fill_1 FILLER_36_967 ();
 sg13g2_fill_2 FILLER_36_984 ();
 sg13g2_fill_1 FILLER_36_986 ();
 sg13g2_fill_2 FILLER_36_998 ();
 sg13g2_fill_1 FILLER_36_1000 ();
 sg13g2_decap_4 FILLER_36_1037 ();
 sg13g2_fill_2 FILLER_36_1041 ();
 sg13g2_decap_8 FILLER_36_1069 ();
 sg13g2_decap_8 FILLER_36_1076 ();
 sg13g2_decap_4 FILLER_36_1083 ();
 sg13g2_fill_2 FILLER_36_1087 ();
 sg13g2_fill_2 FILLER_36_1120 ();
 sg13g2_fill_1 FILLER_36_1122 ();
 sg13g2_fill_2 FILLER_36_1137 ();
 sg13g2_fill_1 FILLER_36_1151 ();
 sg13g2_fill_2 FILLER_36_1187 ();
 sg13g2_decap_4 FILLER_36_1199 ();
 sg13g2_fill_1 FILLER_36_1203 ();
 sg13g2_fill_2 FILLER_36_1230 ();
 sg13g2_fill_1 FILLER_36_1232 ();
 sg13g2_fill_1 FILLER_36_1289 ();
 sg13g2_decap_8 FILLER_36_1295 ();
 sg13g2_decap_8 FILLER_36_1307 ();
 sg13g2_fill_1 FILLER_36_1314 ();
 sg13g2_fill_2 FILLER_36_1320 ();
 sg13g2_fill_1 FILLER_36_1322 ();
 sg13g2_fill_2 FILLER_36_1327 ();
 sg13g2_fill_1 FILLER_36_1339 ();
 sg13g2_fill_2 FILLER_36_1343 ();
 sg13g2_fill_1 FILLER_36_1354 ();
 sg13g2_decap_8 FILLER_36_1416 ();
 sg13g2_decap_8 FILLER_36_1423 ();
 sg13g2_decap_8 FILLER_36_1430 ();
 sg13g2_fill_2 FILLER_36_1437 ();
 sg13g2_fill_1 FILLER_36_1453 ();
 sg13g2_fill_1 FILLER_36_1489 ();
 sg13g2_decap_8 FILLER_36_1494 ();
 sg13g2_decap_8 FILLER_36_1501 ();
 sg13g2_decap_8 FILLER_36_1508 ();
 sg13g2_decap_8 FILLER_36_1515 ();
 sg13g2_fill_2 FILLER_36_1522 ();
 sg13g2_decap_8 FILLER_36_1559 ();
 sg13g2_decap_8 FILLER_36_1566 ();
 sg13g2_fill_1 FILLER_36_1573 ();
 sg13g2_fill_1 FILLER_36_1578 ();
 sg13g2_decap_8 FILLER_36_1583 ();
 sg13g2_decap_8 FILLER_36_1590 ();
 sg13g2_decap_8 FILLER_36_1597 ();
 sg13g2_decap_4 FILLER_36_1604 ();
 sg13g2_fill_2 FILLER_36_1608 ();
 sg13g2_fill_2 FILLER_36_1619 ();
 sg13g2_decap_8 FILLER_36_1647 ();
 sg13g2_decap_4 FILLER_36_1654 ();
 sg13g2_fill_2 FILLER_36_1666 ();
 sg13g2_decap_8 FILLER_36_1673 ();
 sg13g2_decap_4 FILLER_36_1680 ();
 sg13g2_fill_2 FILLER_36_1684 ();
 sg13g2_decap_8 FILLER_36_1715 ();
 sg13g2_decap_8 FILLER_36_1722 ();
 sg13g2_decap_8 FILLER_36_1729 ();
 sg13g2_fill_2 FILLER_36_1736 ();
 sg13g2_fill_2 FILLER_36_1743 ();
 sg13g2_fill_2 FILLER_36_1753 ();
 sg13g2_fill_1 FILLER_36_1755 ();
 sg13g2_fill_2 FILLER_36_1762 ();
 sg13g2_decap_4 FILLER_36_1787 ();
 sg13g2_fill_2 FILLER_36_1791 ();
 sg13g2_decap_8 FILLER_36_1805 ();
 sg13g2_fill_1 FILLER_36_1812 ();
 sg13g2_decap_8 FILLER_36_1853 ();
 sg13g2_decap_8 FILLER_36_1860 ();
 sg13g2_decap_8 FILLER_36_1867 ();
 sg13g2_decap_4 FILLER_36_1874 ();
 sg13g2_fill_2 FILLER_36_1878 ();
 sg13g2_fill_2 FILLER_36_1912 ();
 sg13g2_fill_2 FILLER_36_1919 ();
 sg13g2_fill_2 FILLER_36_1947 ();
 sg13g2_fill_2 FILLER_36_1955 ();
 sg13g2_fill_1 FILLER_36_1957 ();
 sg13g2_decap_8 FILLER_36_1963 ();
 sg13g2_fill_1 FILLER_36_1970 ();
 sg13g2_decap_8 FILLER_36_2002 ();
 sg13g2_decap_8 FILLER_36_2009 ();
 sg13g2_decap_4 FILLER_36_2016 ();
 sg13g2_fill_2 FILLER_36_2020 ();
 sg13g2_decap_8 FILLER_36_2048 ();
 sg13g2_decap_8 FILLER_36_2055 ();
 sg13g2_fill_2 FILLER_36_2062 ();
 sg13g2_fill_1 FILLER_36_2064 ();
 sg13g2_decap_4 FILLER_36_2071 ();
 sg13g2_fill_1 FILLER_36_2075 ();
 sg13g2_decap_4 FILLER_36_2139 ();
 sg13g2_fill_2 FILLER_36_2156 ();
 sg13g2_fill_2 FILLER_36_2194 ();
 sg13g2_fill_1 FILLER_36_2254 ();
 sg13g2_fill_2 FILLER_36_2261 ();
 sg13g2_fill_1 FILLER_36_2263 ();
 sg13g2_fill_1 FILLER_36_2327 ();
 sg13g2_decap_8 FILLER_36_2337 ();
 sg13g2_decap_8 FILLER_36_2344 ();
 sg13g2_fill_1 FILLER_36_2351 ();
 sg13g2_fill_1 FILLER_36_2389 ();
 sg13g2_fill_1 FILLER_36_2399 ();
 sg13g2_fill_1 FILLER_36_2429 ();
 sg13g2_fill_2 FILLER_36_2434 ();
 sg13g2_fill_1 FILLER_36_2445 ();
 sg13g2_fill_1 FILLER_36_2498 ();
 sg13g2_fill_2 FILLER_36_2506 ();
 sg13g2_fill_1 FILLER_36_2508 ();
 sg13g2_decap_8 FILLER_36_2535 ();
 sg13g2_decap_8 FILLER_36_2542 ();
 sg13g2_decap_8 FILLER_36_2549 ();
 sg13g2_decap_8 FILLER_36_2556 ();
 sg13g2_decap_8 FILLER_36_2563 ();
 sg13g2_decap_8 FILLER_36_2570 ();
 sg13g2_decap_8 FILLER_36_2577 ();
 sg13g2_decap_8 FILLER_36_2584 ();
 sg13g2_decap_8 FILLER_36_2591 ();
 sg13g2_decap_8 FILLER_36_2598 ();
 sg13g2_decap_8 FILLER_36_2605 ();
 sg13g2_decap_8 FILLER_36_2612 ();
 sg13g2_decap_8 FILLER_36_2619 ();
 sg13g2_decap_8 FILLER_36_2626 ();
 sg13g2_decap_8 FILLER_36_2633 ();
 sg13g2_decap_8 FILLER_36_2640 ();
 sg13g2_decap_8 FILLER_36_2647 ();
 sg13g2_decap_8 FILLER_36_2654 ();
 sg13g2_decap_8 FILLER_36_2661 ();
 sg13g2_fill_2 FILLER_36_2668 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_30 ();
 sg13g2_fill_1 FILLER_37_43 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_76 ();
 sg13g2_decap_8 FILLER_37_107 ();
 sg13g2_decap_8 FILLER_37_114 ();
 sg13g2_fill_2 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_decap_8 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_decap_4 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_decap_4 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_fill_2 FILLER_37_329 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_412 ();
 sg13g2_decap_8 FILLER_37_419 ();
 sg13g2_decap_4 FILLER_37_426 ();
 sg13g2_fill_1 FILLER_37_430 ();
 sg13g2_decap_8 FILLER_37_471 ();
 sg13g2_decap_8 FILLER_37_478 ();
 sg13g2_fill_2 FILLER_37_485 ();
 sg13g2_fill_1 FILLER_37_487 ();
 sg13g2_fill_2 FILLER_37_498 ();
 sg13g2_fill_1 FILLER_37_520 ();
 sg13g2_fill_2 FILLER_37_525 ();
 sg13g2_fill_1 FILLER_37_527 ();
 sg13g2_decap_4 FILLER_37_532 ();
 sg13g2_fill_1 FILLER_37_536 ();
 sg13g2_decap_8 FILLER_37_555 ();
 sg13g2_decap_8 FILLER_37_562 ();
 sg13g2_decap_4 FILLER_37_569 ();
 sg13g2_fill_1 FILLER_37_573 ();
 sg13g2_decap_4 FILLER_37_578 ();
 sg13g2_fill_1 FILLER_37_582 ();
 sg13g2_fill_2 FILLER_37_601 ();
 sg13g2_fill_1 FILLER_37_603 ();
 sg13g2_decap_4 FILLER_37_638 ();
 sg13g2_fill_2 FILLER_37_642 ();
 sg13g2_fill_1 FILLER_37_652 ();
 sg13g2_decap_8 FILLER_37_667 ();
 sg13g2_fill_2 FILLER_37_674 ();
 sg13g2_fill_1 FILLER_37_676 ();
 sg13g2_decap_8 FILLER_37_682 ();
 sg13g2_decap_8 FILLER_37_689 ();
 sg13g2_fill_1 FILLER_37_696 ();
 sg13g2_decap_4 FILLER_37_731 ();
 sg13g2_fill_1 FILLER_37_747 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_fill_2 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_fill_2 FILLER_37_776 ();
 sg13g2_decap_8 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_fill_2 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_873 ();
 sg13g2_fill_2 FILLER_37_880 ();
 sg13g2_fill_1 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_4 FILLER_37_924 ();
 sg13g2_fill_1 FILLER_37_928 ();
 sg13g2_decap_8 FILLER_37_933 ();
 sg13g2_fill_1 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_949 ();
 sg13g2_decap_8 FILLER_37_956 ();
 sg13g2_decap_8 FILLER_37_963 ();
 sg13g2_decap_8 FILLER_37_970 ();
 sg13g2_decap_8 FILLER_37_977 ();
 sg13g2_decap_8 FILLER_37_984 ();
 sg13g2_decap_4 FILLER_37_991 ();
 sg13g2_fill_1 FILLER_37_1004 ();
 sg13g2_fill_1 FILLER_37_1010 ();
 sg13g2_decap_4 FILLER_37_1020 ();
 sg13g2_fill_2 FILLER_37_1024 ();
 sg13g2_decap_8 FILLER_37_1043 ();
 sg13g2_fill_1 FILLER_37_1054 ();
 sg13g2_decap_4 FILLER_37_1086 ();
 sg13g2_fill_1 FILLER_37_1090 ();
 sg13g2_decap_4 FILLER_37_1099 ();
 sg13g2_fill_2 FILLER_37_1103 ();
 sg13g2_fill_1 FILLER_37_1142 ();
 sg13g2_decap_4 FILLER_37_1162 ();
 sg13g2_fill_2 FILLER_37_1166 ();
 sg13g2_fill_1 FILLER_37_1199 ();
 sg13g2_decap_4 FILLER_37_1206 ();
 sg13g2_fill_2 FILLER_37_1214 ();
 sg13g2_decap_8 FILLER_37_1219 ();
 sg13g2_fill_1 FILLER_37_1226 ();
 sg13g2_fill_1 FILLER_37_1232 ();
 sg13g2_fill_1 FILLER_37_1239 ();
 sg13g2_fill_2 FILLER_37_1246 ();
 sg13g2_decap_4 FILLER_37_1271 ();
 sg13g2_fill_1 FILLER_37_1275 ();
 sg13g2_fill_1 FILLER_37_1306 ();
 sg13g2_fill_1 FILLER_37_1345 ();
 sg13g2_fill_1 FILLER_37_1350 ();
 sg13g2_fill_1 FILLER_37_1356 ();
 sg13g2_fill_2 FILLER_37_1390 ();
 sg13g2_fill_2 FILLER_37_1405 ();
 sg13g2_fill_2 FILLER_37_1411 ();
 sg13g2_fill_1 FILLER_37_1413 ();
 sg13g2_fill_2 FILLER_37_1418 ();
 sg13g2_decap_8 FILLER_37_1449 ();
 sg13g2_fill_1 FILLER_37_1456 ();
 sg13g2_fill_2 FILLER_37_1505 ();
 sg13g2_decap_8 FILLER_37_1511 ();
 sg13g2_decap_4 FILLER_37_1518 ();
 sg13g2_fill_1 FILLER_37_1522 ();
 sg13g2_fill_2 FILLER_37_1534 ();
 sg13g2_fill_1 FILLER_37_1536 ();
 sg13g2_fill_2 FILLER_37_1550 ();
 sg13g2_fill_1 FILLER_37_1552 ();
 sg13g2_fill_2 FILLER_37_1562 ();
 sg13g2_fill_1 FILLER_37_1564 ();
 sg13g2_decap_8 FILLER_37_1594 ();
 sg13g2_decap_8 FILLER_37_1630 ();
 sg13g2_fill_1 FILLER_37_1637 ();
 sg13g2_decap_8 FILLER_37_1647 ();
 sg13g2_fill_2 FILLER_37_1667 ();
 sg13g2_decap_8 FILLER_37_1695 ();
 sg13g2_decap_4 FILLER_37_1702 ();
 sg13g2_fill_2 FILLER_37_1706 ();
 sg13g2_decap_4 FILLER_37_1734 ();
 sg13g2_fill_1 FILLER_37_1764 ();
 sg13g2_fill_2 FILLER_37_1791 ();
 sg13g2_fill_2 FILLER_37_1807 ();
 sg13g2_fill_1 FILLER_37_1816 ();
 sg13g2_decap_8 FILLER_37_1835 ();
 sg13g2_decap_8 FILLER_37_1842 ();
 sg13g2_decap_4 FILLER_37_1853 ();
 sg13g2_fill_2 FILLER_37_1862 ();
 sg13g2_decap_8 FILLER_37_1935 ();
 sg13g2_fill_2 FILLER_37_1942 ();
 sg13g2_fill_1 FILLER_37_1944 ();
 sg13g2_fill_2 FILLER_37_1953 ();
 sg13g2_fill_1 FILLER_37_1955 ();
 sg13g2_fill_2 FILLER_37_1980 ();
 sg13g2_fill_1 FILLER_37_2012 ();
 sg13g2_decap_8 FILLER_37_2018 ();
 sg13g2_fill_2 FILLER_37_2025 ();
 sg13g2_fill_1 FILLER_37_2027 ();
 sg13g2_decap_8 FILLER_37_2033 ();
 sg13g2_decap_4 FILLER_37_2040 ();
 sg13g2_fill_1 FILLER_37_2044 ();
 sg13g2_decap_4 FILLER_37_2050 ();
 sg13g2_fill_1 FILLER_37_2054 ();
 sg13g2_fill_2 FILLER_37_2059 ();
 sg13g2_fill_2 FILLER_37_2072 ();
 sg13g2_fill_2 FILLER_37_2077 ();
 sg13g2_fill_1 FILLER_37_2126 ();
 sg13g2_decap_8 FILLER_37_2153 ();
 sg13g2_fill_1 FILLER_37_2160 ();
 sg13g2_decap_4 FILLER_37_2165 ();
 sg13g2_fill_1 FILLER_37_2169 ();
 sg13g2_fill_2 FILLER_37_2174 ();
 sg13g2_fill_1 FILLER_37_2176 ();
 sg13g2_decap_8 FILLER_37_2222 ();
 sg13g2_fill_2 FILLER_37_2229 ();
 sg13g2_fill_1 FILLER_37_2245 ();
 sg13g2_fill_2 FILLER_37_2252 ();
 sg13g2_fill_1 FILLER_37_2254 ();
 sg13g2_fill_1 FILLER_37_2260 ();
 sg13g2_fill_2 FILLER_37_2291 ();
 sg13g2_fill_1 FILLER_37_2293 ();
 sg13g2_decap_4 FILLER_37_2337 ();
 sg13g2_fill_1 FILLER_37_2341 ();
 sg13g2_fill_2 FILLER_37_2348 ();
 sg13g2_fill_1 FILLER_37_2350 ();
 sg13g2_fill_2 FILLER_37_2369 ();
 sg13g2_fill_1 FILLER_37_2371 ();
 sg13g2_fill_1 FILLER_37_2378 ();
 sg13g2_fill_2 FILLER_37_2411 ();
 sg13g2_fill_2 FILLER_37_2437 ();
 sg13g2_fill_2 FILLER_37_2478 ();
 sg13g2_decap_8 FILLER_37_2542 ();
 sg13g2_decap_8 FILLER_37_2549 ();
 sg13g2_decap_8 FILLER_37_2556 ();
 sg13g2_decap_8 FILLER_37_2563 ();
 sg13g2_decap_8 FILLER_37_2570 ();
 sg13g2_decap_8 FILLER_37_2577 ();
 sg13g2_decap_8 FILLER_37_2584 ();
 sg13g2_decap_8 FILLER_37_2591 ();
 sg13g2_decap_8 FILLER_37_2598 ();
 sg13g2_decap_8 FILLER_37_2605 ();
 sg13g2_decap_8 FILLER_37_2612 ();
 sg13g2_decap_8 FILLER_37_2619 ();
 sg13g2_decap_8 FILLER_37_2626 ();
 sg13g2_decap_8 FILLER_37_2633 ();
 sg13g2_decap_8 FILLER_37_2640 ();
 sg13g2_decap_8 FILLER_37_2647 ();
 sg13g2_decap_8 FILLER_37_2654 ();
 sg13g2_decap_8 FILLER_37_2661 ();
 sg13g2_fill_2 FILLER_37_2668 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_15 ();
 sg13g2_fill_1 FILLER_38_24 ();
 sg13g2_fill_1 FILLER_38_29 ();
 sg13g2_decap_4 FILLER_38_44 ();
 sg13g2_fill_1 FILLER_38_48 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_65 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_decap_8 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_169 ();
 sg13g2_fill_2 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_209 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_409 ();
 sg13g2_decap_4 FILLER_38_416 ();
 sg13g2_fill_1 FILLER_38_420 ();
 sg13g2_decap_4 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_442 ();
 sg13g2_decap_8 FILLER_38_449 ();
 sg13g2_decap_8 FILLER_38_466 ();
 sg13g2_decap_8 FILLER_38_473 ();
 sg13g2_decap_8 FILLER_38_480 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_decap_4 FILLER_38_536 ();
 sg13g2_fill_2 FILLER_38_540 ();
 sg13g2_decap_8 FILLER_38_550 ();
 sg13g2_fill_2 FILLER_38_557 ();
 sg13g2_fill_1 FILLER_38_559 ();
 sg13g2_decap_8 FILLER_38_568 ();
 sg13g2_fill_2 FILLER_38_575 ();
 sg13g2_fill_2 FILLER_38_581 ();
 sg13g2_fill_1 FILLER_38_583 ();
 sg13g2_fill_2 FILLER_38_592 ();
 sg13g2_decap_4 FILLER_38_609 ();
 sg13g2_fill_1 FILLER_38_613 ();
 sg13g2_decap_8 FILLER_38_622 ();
 sg13g2_fill_2 FILLER_38_629 ();
 sg13g2_fill_2 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_682 ();
 sg13g2_decap_8 FILLER_38_689 ();
 sg13g2_decap_8 FILLER_38_696 ();
 sg13g2_fill_2 FILLER_38_703 ();
 sg13g2_decap_8 FILLER_38_713 ();
 sg13g2_fill_2 FILLER_38_720 ();
 sg13g2_decap_8 FILLER_38_734 ();
 sg13g2_decap_4 FILLER_38_741 ();
 sg13g2_fill_1 FILLER_38_745 ();
 sg13g2_decap_8 FILLER_38_751 ();
 sg13g2_decap_8 FILLER_38_758 ();
 sg13g2_decap_4 FILLER_38_765 ();
 sg13g2_fill_1 FILLER_38_769 ();
 sg13g2_fill_2 FILLER_38_835 ();
 sg13g2_decap_8 FILLER_38_878 ();
 sg13g2_decap_8 FILLER_38_885 ();
 sg13g2_decap_8 FILLER_38_892 ();
 sg13g2_fill_2 FILLER_38_899 ();
 sg13g2_fill_1 FILLER_38_901 ();
 sg13g2_decap_4 FILLER_38_918 ();
 sg13g2_decap_4 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_962 ();
 sg13g2_decap_4 FILLER_38_969 ();
 sg13g2_fill_2 FILLER_38_973 ();
 sg13g2_fill_1 FILLER_38_1042 ();
 sg13g2_decap_4 FILLER_38_1049 ();
 sg13g2_decap_8 FILLER_38_1062 ();
 sg13g2_decap_8 FILLER_38_1069 ();
 sg13g2_fill_2 FILLER_38_1076 ();
 sg13g2_decap_8 FILLER_38_1090 ();
 sg13g2_decap_8 FILLER_38_1097 ();
 sg13g2_fill_2 FILLER_38_1104 ();
 sg13g2_fill_1 FILLER_38_1106 ();
 sg13g2_fill_2 FILLER_38_1112 ();
 sg13g2_fill_1 FILLER_38_1114 ();
 sg13g2_decap_4 FILLER_38_1119 ();
 sg13g2_fill_2 FILLER_38_1123 ();
 sg13g2_decap_8 FILLER_38_1174 ();
 sg13g2_fill_2 FILLER_38_1211 ();
 sg13g2_decap_4 FILLER_38_1225 ();
 sg13g2_fill_1 FILLER_38_1229 ();
 sg13g2_fill_1 FILLER_38_1234 ();
 sg13g2_fill_1 FILLER_38_1240 ();
 sg13g2_fill_2 FILLER_38_1249 ();
 sg13g2_fill_1 FILLER_38_1255 ();
 sg13g2_fill_2 FILLER_38_1282 ();
 sg13g2_fill_2 FILLER_38_1296 ();
 sg13g2_fill_1 FILLER_38_1302 ();
 sg13g2_fill_1 FILLER_38_1365 ();
 sg13g2_fill_1 FILLER_38_1385 ();
 sg13g2_fill_2 FILLER_38_1425 ();
 sg13g2_decap_8 FILLER_38_1431 ();
 sg13g2_decap_8 FILLER_38_1438 ();
 sg13g2_decap_8 FILLER_38_1445 ();
 sg13g2_decap_8 FILLER_38_1452 ();
 sg13g2_fill_1 FILLER_38_1459 ();
 sg13g2_decap_4 FILLER_38_1494 ();
 sg13g2_decap_4 FILLER_38_1502 ();
 sg13g2_fill_2 FILLER_38_1506 ();
 sg13g2_decap_8 FILLER_38_1512 ();
 sg13g2_decap_8 FILLER_38_1519 ();
 sg13g2_decap_8 FILLER_38_1526 ();
 sg13g2_decap_8 FILLER_38_1533 ();
 sg13g2_fill_2 FILLER_38_1540 ();
 sg13g2_fill_2 FILLER_38_1573 ();
 sg13g2_decap_8 FILLER_38_1601 ();
 sg13g2_decap_8 FILLER_38_1608 ();
 sg13g2_decap_8 FILLER_38_1615 ();
 sg13g2_fill_2 FILLER_38_1622 ();
 sg13g2_fill_1 FILLER_38_1659 ();
 sg13g2_fill_2 FILLER_38_1669 ();
 sg13g2_decap_8 FILLER_38_1676 ();
 sg13g2_decap_4 FILLER_38_1683 ();
 sg13g2_fill_1 FILLER_38_1700 ();
 sg13g2_decap_4 FILLER_38_1727 ();
 sg13g2_fill_2 FILLER_38_1731 ();
 sg13g2_fill_2 FILLER_38_1751 ();
 sg13g2_fill_1 FILLER_38_1753 ();
 sg13g2_fill_1 FILLER_38_1759 ();
 sg13g2_decap_8 FILLER_38_1786 ();
 sg13g2_fill_2 FILLER_38_1793 ();
 sg13g2_fill_1 FILLER_38_1824 ();
 sg13g2_decap_4 FILLER_38_1857 ();
 sg13g2_decap_8 FILLER_38_1887 ();
 sg13g2_fill_1 FILLER_38_1894 ();
 sg13g2_decap_4 FILLER_38_1900 ();
 sg13g2_decap_4 FILLER_38_1908 ();
 sg13g2_decap_8 FILLER_38_1917 ();
 sg13g2_decap_8 FILLER_38_1924 ();
 sg13g2_decap_8 FILLER_38_1931 ();
 sg13g2_decap_8 FILLER_38_1938 ();
 sg13g2_fill_2 FILLER_38_1945 ();
 sg13g2_fill_1 FILLER_38_1947 ();
 sg13g2_decap_4 FILLER_38_1966 ();
 sg13g2_fill_1 FILLER_38_1970 ();
 sg13g2_fill_2 FILLER_38_1986 ();
 sg13g2_decap_8 FILLER_38_2000 ();
 sg13g2_fill_1 FILLER_38_2007 ();
 sg13g2_decap_8 FILLER_38_2016 ();
 sg13g2_decap_8 FILLER_38_2023 ();
 sg13g2_fill_1 FILLER_38_2074 ();
 sg13g2_fill_1 FILLER_38_2116 ();
 sg13g2_fill_2 FILLER_38_2123 ();
 sg13g2_fill_2 FILLER_38_2131 ();
 sg13g2_fill_2 FILLER_38_2159 ();
 sg13g2_fill_2 FILLER_38_2200 ();
 sg13g2_fill_1 FILLER_38_2202 ();
 sg13g2_fill_2 FILLER_38_2234 ();
 sg13g2_decap_8 FILLER_38_2267 ();
 sg13g2_decap_8 FILLER_38_2274 ();
 sg13g2_decap_8 FILLER_38_2281 ();
 sg13g2_decap_8 FILLER_38_2288 ();
 sg13g2_fill_2 FILLER_38_2295 ();
 sg13g2_fill_1 FILLER_38_2297 ();
 sg13g2_fill_2 FILLER_38_2310 ();
 sg13g2_fill_1 FILLER_38_2325 ();
 sg13g2_fill_2 FILLER_38_2391 ();
 sg13g2_fill_2 FILLER_38_2434 ();
 sg13g2_decap_4 FILLER_38_2473 ();
 sg13g2_fill_2 FILLER_38_2477 ();
 sg13g2_decap_4 FILLER_38_2522 ();
 sg13g2_fill_1 FILLER_38_2526 ();
 sg13g2_fill_1 FILLER_38_2531 ();
 sg13g2_decap_8 FILLER_38_2562 ();
 sg13g2_decap_8 FILLER_38_2569 ();
 sg13g2_decap_8 FILLER_38_2576 ();
 sg13g2_decap_8 FILLER_38_2583 ();
 sg13g2_decap_8 FILLER_38_2590 ();
 sg13g2_decap_8 FILLER_38_2597 ();
 sg13g2_decap_8 FILLER_38_2604 ();
 sg13g2_decap_8 FILLER_38_2611 ();
 sg13g2_decap_8 FILLER_38_2618 ();
 sg13g2_decap_8 FILLER_38_2625 ();
 sg13g2_decap_8 FILLER_38_2632 ();
 sg13g2_decap_8 FILLER_38_2639 ();
 sg13g2_decap_8 FILLER_38_2646 ();
 sg13g2_decap_8 FILLER_38_2653 ();
 sg13g2_decap_8 FILLER_38_2660 ();
 sg13g2_fill_2 FILLER_38_2667 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_4 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_25 ();
 sg13g2_decap_8 FILLER_39_34 ();
 sg13g2_decap_8 FILLER_39_41 ();
 sg13g2_fill_2 FILLER_39_48 ();
 sg13g2_fill_1 FILLER_39_50 ();
 sg13g2_decap_8 FILLER_39_171 ();
 sg13g2_fill_1 FILLER_39_178 ();
 sg13g2_decap_8 FILLER_39_183 ();
 sg13g2_fill_2 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_198 ();
 sg13g2_decap_4 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_decap_4 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_264 ();
 sg13g2_decap_4 FILLER_39_271 ();
 sg13g2_fill_1 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_291 ();
 sg13g2_fill_2 FILLER_39_297 ();
 sg13g2_fill_1 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_350 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_373 ();
 sg13g2_fill_1 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_fill_1 FILLER_39_400 ();
 sg13g2_decap_8 FILLER_39_410 ();
 sg13g2_decap_4 FILLER_39_417 ();
 sg13g2_fill_1 FILLER_39_421 ();
 sg13g2_fill_1 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_445 ();
 sg13g2_fill_2 FILLER_39_452 ();
 sg13g2_fill_1 FILLER_39_454 ();
 sg13g2_fill_2 FILLER_39_481 ();
 sg13g2_fill_1 FILLER_39_483 ();
 sg13g2_fill_2 FILLER_39_501 ();
 sg13g2_fill_1 FILLER_39_503 ();
 sg13g2_fill_1 FILLER_39_519 ();
 sg13g2_decap_4 FILLER_39_526 ();
 sg13g2_fill_2 FILLER_39_530 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_8 FILLER_39_543 ();
 sg13g2_decap_4 FILLER_39_550 ();
 sg13g2_fill_2 FILLER_39_554 ();
 sg13g2_decap_4 FILLER_39_569 ();
 sg13g2_fill_2 FILLER_39_573 ();
 sg13g2_decap_8 FILLER_39_579 ();
 sg13g2_fill_2 FILLER_39_586 ();
 sg13g2_fill_1 FILLER_39_588 ();
 sg13g2_decap_4 FILLER_39_594 ();
 sg13g2_fill_1 FILLER_39_598 ();
 sg13g2_decap_8 FILLER_39_604 ();
 sg13g2_decap_8 FILLER_39_611 ();
 sg13g2_decap_8 FILLER_39_618 ();
 sg13g2_decap_8 FILLER_39_625 ();
 sg13g2_decap_4 FILLER_39_636 ();
 sg13g2_fill_2 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_682 ();
 sg13g2_decap_8 FILLER_39_689 ();
 sg13g2_fill_2 FILLER_39_696 ();
 sg13g2_decap_4 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_fill_1 FILLER_39_849 ();
 sg13g2_decap_8 FILLER_39_902 ();
 sg13g2_decap_8 FILLER_39_909 ();
 sg13g2_decap_8 FILLER_39_916 ();
 sg13g2_decap_4 FILLER_39_923 ();
 sg13g2_fill_2 FILLER_39_931 ();
 sg13g2_fill_1 FILLER_39_939 ();
 sg13g2_fill_2 FILLER_39_946 ();
 sg13g2_fill_1 FILLER_39_948 ();
 sg13g2_fill_2 FILLER_39_957 ();
 sg13g2_fill_1 FILLER_39_965 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_4 FILLER_39_992 ();
 sg13g2_decap_4 FILLER_39_1001 ();
 sg13g2_fill_1 FILLER_39_1014 ();
 sg13g2_decap_8 FILLER_39_1068 ();
 sg13g2_fill_2 FILLER_39_1075 ();
 sg13g2_fill_1 FILLER_39_1077 ();
 sg13g2_decap_4 FILLER_39_1090 ();
 sg13g2_fill_1 FILLER_39_1094 ();
 sg13g2_decap_8 FILLER_39_1107 ();
 sg13g2_decap_8 FILLER_39_1114 ();
 sg13g2_fill_1 FILLER_39_1121 ();
 sg13g2_decap_4 FILLER_39_1127 ();
 sg13g2_fill_2 FILLER_39_1135 ();
 sg13g2_fill_1 FILLER_39_1137 ();
 sg13g2_decap_8 FILLER_39_1142 ();
 sg13g2_fill_1 FILLER_39_1149 ();
 sg13g2_decap_8 FILLER_39_1154 ();
 sg13g2_decap_8 FILLER_39_1161 ();
 sg13g2_decap_8 FILLER_39_1168 ();
 sg13g2_fill_2 FILLER_39_1175 ();
 sg13g2_decap_8 FILLER_39_1194 ();
 sg13g2_decap_4 FILLER_39_1201 ();
 sg13g2_fill_2 FILLER_39_1205 ();
 sg13g2_decap_4 FILLER_39_1211 ();
 sg13g2_fill_1 FILLER_39_1215 ();
 sg13g2_fill_1 FILLER_39_1242 ();
 sg13g2_fill_2 FILLER_39_1249 ();
 sg13g2_fill_2 FILLER_39_1256 ();
 sg13g2_fill_2 FILLER_39_1263 ();
 sg13g2_decap_8 FILLER_39_1269 ();
 sg13g2_decap_8 FILLER_39_1276 ();
 sg13g2_fill_2 FILLER_39_1283 ();
 sg13g2_fill_1 FILLER_39_1285 ();
 sg13g2_decap_8 FILLER_39_1290 ();
 sg13g2_decap_8 FILLER_39_1316 ();
 sg13g2_decap_8 FILLER_39_1329 ();
 sg13g2_fill_1 FILLER_39_1336 ();
 sg13g2_decap_8 FILLER_39_1342 ();
 sg13g2_fill_1 FILLER_39_1349 ();
 sg13g2_decap_8 FILLER_39_1354 ();
 sg13g2_fill_1 FILLER_39_1361 ();
 sg13g2_fill_2 FILLER_39_1369 ();
 sg13g2_fill_1 FILLER_39_1408 ();
 sg13g2_fill_1 FILLER_39_1457 ();
 sg13g2_fill_1 FILLER_39_1468 ();
 sg13g2_decap_8 FILLER_39_1495 ();
 sg13g2_fill_2 FILLER_39_1507 ();
 sg13g2_decap_4 FILLER_39_1535 ();
 sg13g2_fill_2 FILLER_39_1552 ();
 sg13g2_fill_1 FILLER_39_1588 ();
 sg13g2_decap_4 FILLER_39_1624 ();
 sg13g2_decap_8 FILLER_39_1663 ();
 sg13g2_fill_2 FILLER_39_1670 ();
 sg13g2_decap_8 FILLER_39_1678 ();
 sg13g2_fill_2 FILLER_39_1685 ();
 sg13g2_fill_2 FILLER_39_1693 ();
 sg13g2_fill_1 FILLER_39_1706 ();
 sg13g2_fill_2 FILLER_39_1720 ();
 sg13g2_fill_1 FILLER_39_1722 ();
 sg13g2_decap_4 FILLER_39_1738 ();
 sg13g2_fill_2 FILLER_39_1742 ();
 sg13g2_decap_8 FILLER_39_1754 ();
 sg13g2_decap_4 FILLER_39_1761 ();
 sg13g2_fill_1 FILLER_39_1765 ();
 sg13g2_fill_1 FILLER_39_1775 ();
 sg13g2_decap_8 FILLER_39_1786 ();
 sg13g2_decap_4 FILLER_39_1793 ();
 sg13g2_fill_2 FILLER_39_1797 ();
 sg13g2_decap_4 FILLER_39_1804 ();
 sg13g2_fill_1 FILLER_39_1808 ();
 sg13g2_fill_1 FILLER_39_1844 ();
 sg13g2_fill_2 FILLER_39_1881 ();
 sg13g2_decap_8 FILLER_39_1896 ();
 sg13g2_decap_8 FILLER_39_1903 ();
 sg13g2_decap_8 FILLER_39_1910 ();
 sg13g2_fill_1 FILLER_39_1917 ();
 sg13g2_decap_4 FILLER_39_1957 ();
 sg13g2_fill_1 FILLER_39_2001 ();
 sg13g2_fill_2 FILLER_39_2028 ();
 sg13g2_fill_1 FILLER_39_2040 ();
 sg13g2_decap_4 FILLER_39_2067 ();
 sg13g2_fill_2 FILLER_39_2108 ();
 sg13g2_decap_4 FILLER_39_2149 ();
 sg13g2_fill_1 FILLER_39_2153 ();
 sg13g2_decap_4 FILLER_39_2189 ();
 sg13g2_decap_8 FILLER_39_2207 ();
 sg13g2_decap_8 FILLER_39_2214 ();
 sg13g2_decap_8 FILLER_39_2221 ();
 sg13g2_decap_8 FILLER_39_2228 ();
 sg13g2_fill_2 FILLER_39_2235 ();
 sg13g2_decap_8 FILLER_39_2271 ();
 sg13g2_decap_8 FILLER_39_2278 ();
 sg13g2_decap_8 FILLER_39_2285 ();
 sg13g2_decap_4 FILLER_39_2292 ();
 sg13g2_fill_2 FILLER_39_2296 ();
 sg13g2_fill_1 FILLER_39_2358 ();
 sg13g2_fill_1 FILLER_39_2388 ();
 sg13g2_fill_1 FILLER_39_2393 ();
 sg13g2_fill_2 FILLER_39_2420 ();
 sg13g2_fill_2 FILLER_39_2428 ();
 sg13g2_decap_8 FILLER_39_2499 ();
 sg13g2_decap_8 FILLER_39_2506 ();
 sg13g2_decap_4 FILLER_39_2513 ();
 sg13g2_fill_1 FILLER_39_2517 ();
 sg13g2_decap_8 FILLER_39_2558 ();
 sg13g2_decap_8 FILLER_39_2565 ();
 sg13g2_decap_8 FILLER_39_2572 ();
 sg13g2_decap_8 FILLER_39_2579 ();
 sg13g2_decap_8 FILLER_39_2586 ();
 sg13g2_decap_8 FILLER_39_2593 ();
 sg13g2_decap_8 FILLER_39_2600 ();
 sg13g2_decap_8 FILLER_39_2607 ();
 sg13g2_decap_8 FILLER_39_2614 ();
 sg13g2_decap_8 FILLER_39_2621 ();
 sg13g2_decap_8 FILLER_39_2628 ();
 sg13g2_decap_8 FILLER_39_2635 ();
 sg13g2_decap_8 FILLER_39_2642 ();
 sg13g2_decap_8 FILLER_39_2649 ();
 sg13g2_decap_8 FILLER_39_2656 ();
 sg13g2_decap_8 FILLER_39_2663 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_2 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_78 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_4 FILLER_40_112 ();
 sg13g2_fill_1 FILLER_40_116 ();
 sg13g2_fill_2 FILLER_40_121 ();
 sg13g2_fill_2 FILLER_40_137 ();
 sg13g2_fill_1 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_148 ();
 sg13g2_decap_8 FILLER_40_187 ();
 sg13g2_decap_8 FILLER_40_194 ();
 sg13g2_decap_4 FILLER_40_201 ();
 sg13g2_fill_1 FILLER_40_234 ();
 sg13g2_decap_4 FILLER_40_244 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_decap_4 FILLER_40_311 ();
 sg13g2_fill_1 FILLER_40_315 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_326 ();
 sg13g2_fill_1 FILLER_40_330 ();
 sg13g2_decap_4 FILLER_40_340 ();
 sg13g2_fill_1 FILLER_40_352 ();
 sg13g2_fill_1 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_391 ();
 sg13g2_fill_2 FILLER_40_402 ();
 sg13g2_fill_1 FILLER_40_404 ();
 sg13g2_decap_8 FILLER_40_446 ();
 sg13g2_decap_8 FILLER_40_453 ();
 sg13g2_fill_2 FILLER_40_460 ();
 sg13g2_fill_1 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_473 ();
 sg13g2_decap_8 FILLER_40_480 ();
 sg13g2_decap_8 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_494 ();
 sg13g2_fill_2 FILLER_40_499 ();
 sg13g2_fill_2 FILLER_40_506 ();
 sg13g2_fill_1 FILLER_40_517 ();
 sg13g2_fill_2 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_552 ();
 sg13g2_decap_4 FILLER_40_557 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_4 FILLER_40_581 ();
 sg13g2_decap_4 FILLER_40_593 ();
 sg13g2_decap_8 FILLER_40_606 ();
 sg13g2_decap_8 FILLER_40_613 ();
 sg13g2_decap_8 FILLER_40_620 ();
 sg13g2_decap_4 FILLER_40_627 ();
 sg13g2_fill_2 FILLER_40_631 ();
 sg13g2_fill_1 FILLER_40_638 ();
 sg13g2_fill_1 FILLER_40_647 ();
 sg13g2_fill_1 FILLER_40_656 ();
 sg13g2_fill_2 FILLER_40_661 ();
 sg13g2_fill_1 FILLER_40_676 ();
 sg13g2_fill_2 FILLER_40_688 ();
 sg13g2_decap_8 FILLER_40_695 ();
 sg13g2_fill_2 FILLER_40_702 ();
 sg13g2_fill_2 FILLER_40_730 ();
 sg13g2_fill_1 FILLER_40_732 ();
 sg13g2_decap_8 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_40_744 ();
 sg13g2_fill_2 FILLER_40_763 ();
 sg13g2_fill_1 FILLER_40_765 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_fill_2 FILLER_40_781 ();
 sg13g2_fill_1 FILLER_40_797 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_fill_2 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_835 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_fill_1 FILLER_40_849 ();
 sg13g2_fill_2 FILLER_40_853 ();
 sg13g2_fill_1 FILLER_40_862 ();
 sg13g2_fill_2 FILLER_40_903 ();
 sg13g2_fill_1 FILLER_40_905 ();
 sg13g2_fill_1 FILLER_40_937 ();
 sg13g2_decap_8 FILLER_40_982 ();
 sg13g2_decap_8 FILLER_40_989 ();
 sg13g2_decap_4 FILLER_40_996 ();
 sg13g2_fill_2 FILLER_40_1012 ();
 sg13g2_fill_2 FILLER_40_1024 ();
 sg13g2_fill_1 FILLER_40_1026 ();
 sg13g2_decap_4 FILLER_40_1048 ();
 sg13g2_decap_4 FILLER_40_1088 ();
 sg13g2_fill_1 FILLER_40_1092 ();
 sg13g2_fill_1 FILLER_40_1111 ();
 sg13g2_decap_8 FILLER_40_1142 ();
 sg13g2_decap_4 FILLER_40_1149 ();
 sg13g2_fill_1 FILLER_40_1153 ();
 sg13g2_decap_4 FILLER_40_1159 ();
 sg13g2_fill_2 FILLER_40_1163 ();
 sg13g2_decap_8 FILLER_40_1174 ();
 sg13g2_decap_8 FILLER_40_1181 ();
 sg13g2_decap_8 FILLER_40_1188 ();
 sg13g2_decap_8 FILLER_40_1195 ();
 sg13g2_fill_1 FILLER_40_1207 ();
 sg13g2_decap_8 FILLER_40_1223 ();
 sg13g2_decap_8 FILLER_40_1256 ();
 sg13g2_decap_8 FILLER_40_1263 ();
 sg13g2_decap_4 FILLER_40_1270 ();
 sg13g2_decap_8 FILLER_40_1282 ();
 sg13g2_fill_1 FILLER_40_1289 ();
 sg13g2_fill_2 FILLER_40_1336 ();
 sg13g2_fill_2 FILLER_40_1342 ();
 sg13g2_fill_2 FILLER_40_1349 ();
 sg13g2_fill_2 FILLER_40_1380 ();
 sg13g2_decap_4 FILLER_40_1395 ();
 sg13g2_fill_1 FILLER_40_1399 ();
 sg13g2_fill_2 FILLER_40_1408 ();
 sg13g2_fill_1 FILLER_40_1410 ();
 sg13g2_fill_2 FILLER_40_1416 ();
 sg13g2_fill_1 FILLER_40_1418 ();
 sg13g2_fill_2 FILLER_40_1423 ();
 sg13g2_fill_1 FILLER_40_1451 ();
 sg13g2_decap_8 FILLER_40_1491 ();
 sg13g2_decap_8 FILLER_40_1498 ();
 sg13g2_decap_4 FILLER_40_1505 ();
 sg13g2_fill_1 FILLER_40_1509 ();
 sg13g2_decap_8 FILLER_40_1536 ();
 sg13g2_fill_2 FILLER_40_1543 ();
 sg13g2_fill_2 FILLER_40_1550 ();
 sg13g2_fill_2 FILLER_40_1569 ();
 sg13g2_fill_2 FILLER_40_1585 ();
 sg13g2_fill_2 FILLER_40_1592 ();
 sg13g2_fill_1 FILLER_40_1602 ();
 sg13g2_fill_2 FILLER_40_1608 ();
 sg13g2_fill_1 FILLER_40_1614 ();
 sg13g2_decap_8 FILLER_40_1624 ();
 sg13g2_decap_8 FILLER_40_1631 ();
 sg13g2_fill_1 FILLER_40_1638 ();
 sg13g2_decap_4 FILLER_40_1649 ();
 sg13g2_fill_1 FILLER_40_1653 ();
 sg13g2_decap_4 FILLER_40_1658 ();
 sg13g2_fill_1 FILLER_40_1662 ();
 sg13g2_fill_2 FILLER_40_1667 ();
 sg13g2_fill_2 FILLER_40_1681 ();
 sg13g2_fill_1 FILLER_40_1683 ();
 sg13g2_decap_4 FILLER_40_1698 ();
 sg13g2_fill_1 FILLER_40_1702 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_4 FILLER_40_1719 ();
 sg13g2_fill_1 FILLER_40_1723 ();
 sg13g2_decap_8 FILLER_40_1750 ();
 sg13g2_decap_8 FILLER_40_1757 ();
 sg13g2_decap_8 FILLER_40_1764 ();
 sg13g2_decap_8 FILLER_40_1771 ();
 sg13g2_decap_8 FILLER_40_1778 ();
 sg13g2_decap_8 FILLER_40_1785 ();
 sg13g2_decap_4 FILLER_40_1792 ();
 sg13g2_fill_1 FILLER_40_1796 ();
 sg13g2_fill_2 FILLER_40_1807 ();
 sg13g2_fill_1 FILLER_40_1809 ();
 sg13g2_fill_2 FILLER_40_1815 ();
 sg13g2_fill_1 FILLER_40_1817 ();
 sg13g2_decap_8 FILLER_40_1827 ();
 sg13g2_decap_4 FILLER_40_1834 ();
 sg13g2_fill_1 FILLER_40_1838 ();
 sg13g2_fill_1 FILLER_40_1843 ();
 sg13g2_fill_1 FILLER_40_1848 ();
 sg13g2_decap_4 FILLER_40_1854 ();
 sg13g2_fill_1 FILLER_40_1858 ();
 sg13g2_fill_2 FILLER_40_1885 ();
 sg13g2_fill_1 FILLER_40_1887 ();
 sg13g2_fill_2 FILLER_40_1921 ();
 sg13g2_fill_2 FILLER_40_1949 ();
 sg13g2_decap_8 FILLER_40_1960 ();
 sg13g2_decap_8 FILLER_40_1967 ();
 sg13g2_fill_1 FILLER_40_1974 ();
 sg13g2_fill_2 FILLER_40_1979 ();
 sg13g2_fill_2 FILLER_40_1989 ();
 sg13g2_fill_1 FILLER_40_1996 ();
 sg13g2_fill_1 FILLER_40_2001 ();
 sg13g2_decap_8 FILLER_40_2006 ();
 sg13g2_fill_1 FILLER_40_2013 ();
 sg13g2_fill_2 FILLER_40_2023 ();
 sg13g2_fill_2 FILLER_40_2029 ();
 sg13g2_decap_8 FILLER_40_2036 ();
 sg13g2_fill_1 FILLER_40_2043 ();
 sg13g2_decap_4 FILLER_40_2061 ();
 sg13g2_fill_2 FILLER_40_2065 ();
 sg13g2_decap_8 FILLER_40_2079 ();
 sg13g2_fill_2 FILLER_40_2086 ();
 sg13g2_fill_1 FILLER_40_2088 ();
 sg13g2_fill_2 FILLER_40_2099 ();
 sg13g2_fill_1 FILLER_40_2110 ();
 sg13g2_decap_4 FILLER_40_2124 ();
 sg13g2_fill_2 FILLER_40_2128 ();
 sg13g2_decap_8 FILLER_40_2147 ();
 sg13g2_decap_8 FILLER_40_2154 ();
 sg13g2_decap_8 FILLER_40_2161 ();
 sg13g2_decap_8 FILLER_40_2168 ();
 sg13g2_decap_8 FILLER_40_2175 ();
 sg13g2_decap_8 FILLER_40_2182 ();
 sg13g2_decap_8 FILLER_40_2189 ();
 sg13g2_decap_8 FILLER_40_2196 ();
 sg13g2_decap_8 FILLER_40_2203 ();
 sg13g2_decap_8 FILLER_40_2210 ();
 sg13g2_decap_8 FILLER_40_2221 ();
 sg13g2_decap_8 FILLER_40_2228 ();
 sg13g2_decap_4 FILLER_40_2235 ();
 sg13g2_fill_2 FILLER_40_2254 ();
 sg13g2_fill_1 FILLER_40_2256 ();
 sg13g2_decap_8 FILLER_40_2283 ();
 sg13g2_decap_4 FILLER_40_2290 ();
 sg13g2_decap_8 FILLER_40_2298 ();
 sg13g2_fill_1 FILLER_40_2305 ();
 sg13g2_decap_4 FILLER_40_2310 ();
 sg13g2_fill_2 FILLER_40_2314 ();
 sg13g2_decap_4 FILLER_40_2325 ();
 sg13g2_fill_2 FILLER_40_2329 ();
 sg13g2_decap_8 FILLER_40_2335 ();
 sg13g2_fill_2 FILLER_40_2342 ();
 sg13g2_fill_2 FILLER_40_2352 ();
 sg13g2_fill_1 FILLER_40_2354 ();
 sg13g2_decap_8 FILLER_40_2360 ();
 sg13g2_decap_8 FILLER_40_2367 ();
 sg13g2_decap_4 FILLER_40_2374 ();
 sg13g2_fill_1 FILLER_40_2378 ();
 sg13g2_decap_8 FILLER_40_2399 ();
 sg13g2_decap_8 FILLER_40_2406 ();
 sg13g2_decap_8 FILLER_40_2413 ();
 sg13g2_fill_2 FILLER_40_2420 ();
 sg13g2_decap_4 FILLER_40_2434 ();
 sg13g2_decap_4 FILLER_40_2442 ();
 sg13g2_fill_2 FILLER_40_2446 ();
 sg13g2_decap_8 FILLER_40_2452 ();
 sg13g2_decap_8 FILLER_40_2459 ();
 sg13g2_decap_4 FILLER_40_2466 ();
 sg13g2_fill_2 FILLER_40_2518 ();
 sg13g2_decap_8 FILLER_40_2554 ();
 sg13g2_decap_8 FILLER_40_2561 ();
 sg13g2_decap_8 FILLER_40_2568 ();
 sg13g2_decap_8 FILLER_40_2575 ();
 sg13g2_decap_8 FILLER_40_2582 ();
 sg13g2_decap_8 FILLER_40_2589 ();
 sg13g2_decap_8 FILLER_40_2596 ();
 sg13g2_decap_8 FILLER_40_2603 ();
 sg13g2_decap_8 FILLER_40_2610 ();
 sg13g2_decap_8 FILLER_40_2617 ();
 sg13g2_decap_8 FILLER_40_2624 ();
 sg13g2_decap_8 FILLER_40_2631 ();
 sg13g2_decap_8 FILLER_40_2638 ();
 sg13g2_decap_8 FILLER_40_2645 ();
 sg13g2_decap_8 FILLER_40_2652 ();
 sg13g2_decap_8 FILLER_40_2659 ();
 sg13g2_decap_4 FILLER_40_2666 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_58 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_decap_8 FILLER_41_99 ();
 sg13g2_decap_8 FILLER_41_106 ();
 sg13g2_decap_8 FILLER_41_113 ();
 sg13g2_decap_8 FILLER_41_120 ();
 sg13g2_decap_8 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_134 ();
 sg13g2_decap_8 FILLER_41_141 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_fill_1 FILLER_41_156 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_fill_2 FILLER_41_174 ();
 sg13g2_fill_1 FILLER_41_213 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_fill_1 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_4 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_249 ();
 sg13g2_fill_2 FILLER_41_274 ();
 sg13g2_fill_2 FILLER_41_297 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_fill_2 FILLER_41_354 ();
 sg13g2_decap_8 FILLER_41_360 ();
 sg13g2_fill_2 FILLER_41_367 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_decap_4 FILLER_41_373 ();
 sg13g2_decap_4 FILLER_41_381 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_41_444 ();
 sg13g2_fill_2 FILLER_41_451 ();
 sg13g2_decap_4 FILLER_41_487 ();
 sg13g2_fill_2 FILLER_41_491 ();
 sg13g2_decap_4 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_501 ();
 sg13g2_decap_4 FILLER_41_507 ();
 sg13g2_fill_1 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_521 ();
 sg13g2_fill_2 FILLER_41_528 ();
 sg13g2_decap_4 FILLER_41_547 ();
 sg13g2_fill_1 FILLER_41_551 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_fill_1 FILLER_41_588 ();
 sg13g2_fill_2 FILLER_41_598 ();
 sg13g2_fill_1 FILLER_41_604 ();
 sg13g2_decap_8 FILLER_41_610 ();
 sg13g2_decap_4 FILLER_41_617 ();
 sg13g2_fill_1 FILLER_41_626 ();
 sg13g2_fill_1 FILLER_41_708 ();
 sg13g2_decap_4 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_755 ();
 sg13g2_decap_8 FILLER_41_762 ();
 sg13g2_fill_1 FILLER_41_769 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_4 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_41_835 ();
 sg13g2_decap_4 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_855 ();
 sg13g2_fill_2 FILLER_41_862 ();
 sg13g2_fill_1 FILLER_41_864 ();
 sg13g2_decap_4 FILLER_41_870 ();
 sg13g2_fill_1 FILLER_41_874 ();
 sg13g2_decap_8 FILLER_41_885 ();
 sg13g2_decap_8 FILLER_41_892 ();
 sg13g2_fill_2 FILLER_41_899 ();
 sg13g2_decap_8 FILLER_41_905 ();
 sg13g2_fill_1 FILLER_41_917 ();
 sg13g2_fill_2 FILLER_41_928 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_fill_1 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_981 ();
 sg13g2_fill_1 FILLER_41_988 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_4 FILLER_41_1029 ();
 sg13g2_decap_8 FILLER_41_1039 ();
 sg13g2_decap_8 FILLER_41_1046 ();
 sg13g2_decap_4 FILLER_41_1053 ();
 sg13g2_decap_4 FILLER_41_1061 ();
 sg13g2_fill_1 FILLER_41_1065 ();
 sg13g2_fill_2 FILLER_41_1152 ();
 sg13g2_fill_1 FILLER_41_1158 ();
 sg13g2_fill_2 FILLER_41_1185 ();
 sg13g2_fill_2 FILLER_41_1213 ();
 sg13g2_decap_8 FILLER_41_1220 ();
 sg13g2_decap_4 FILLER_41_1227 ();
 sg13g2_decap_8 FILLER_41_1235 ();
 sg13g2_decap_4 FILLER_41_1242 ();
 sg13g2_fill_2 FILLER_41_1246 ();
 sg13g2_fill_2 FILLER_41_1257 ();
 sg13g2_fill_2 FILLER_41_1285 ();
 sg13g2_fill_1 FILLER_41_1287 ();
 sg13g2_fill_2 FILLER_41_1292 ();
 sg13g2_fill_1 FILLER_41_1294 ();
 sg13g2_fill_1 FILLER_41_1300 ();
 sg13g2_fill_2 FILLER_41_1347 ();
 sg13g2_fill_1 FILLER_41_1349 ();
 sg13g2_decap_8 FILLER_41_1356 ();
 sg13g2_decap_8 FILLER_41_1367 ();
 sg13g2_fill_2 FILLER_41_1389 ();
 sg13g2_fill_2 FILLER_41_1394 ();
 sg13g2_fill_2 FILLER_41_1405 ();
 sg13g2_fill_1 FILLER_41_1407 ();
 sg13g2_fill_2 FILLER_41_1429 ();
 sg13g2_fill_2 FILLER_41_1440 ();
 sg13g2_fill_2 FILLER_41_1454 ();
 sg13g2_decap_4 FILLER_41_1497 ();
 sg13g2_fill_1 FILLER_41_1501 ();
 sg13g2_fill_2 FILLER_41_1516 ();
 sg13g2_fill_1 FILLER_41_1544 ();
 sg13g2_decap_8 FILLER_41_1549 ();
 sg13g2_decap_8 FILLER_41_1556 ();
 sg13g2_decap_4 FILLER_41_1563 ();
 sg13g2_fill_1 FILLER_41_1567 ();
 sg13g2_fill_2 FILLER_41_1580 ();
 sg13g2_decap_8 FILLER_41_1612 ();
 sg13g2_decap_8 FILLER_41_1619 ();
 sg13g2_decap_8 FILLER_41_1626 ();
 sg13g2_decap_8 FILLER_41_1633 ();
 sg13g2_decap_4 FILLER_41_1640 ();
 sg13g2_fill_2 FILLER_41_1644 ();
 sg13g2_fill_2 FILLER_41_1677 ();
 sg13g2_fill_1 FILLER_41_1679 ();
 sg13g2_decap_8 FILLER_41_1712 ();
 sg13g2_decap_4 FILLER_41_1719 ();
 sg13g2_fill_2 FILLER_41_1723 ();
 sg13g2_fill_2 FILLER_41_1751 ();
 sg13g2_fill_1 FILLER_41_1753 ();
 sg13g2_decap_4 FILLER_41_1794 ();
 sg13g2_fill_2 FILLER_41_1798 ();
 sg13g2_decap_8 FILLER_41_1826 ();
 sg13g2_fill_1 FILLER_41_1833 ();
 sg13g2_decap_8 FILLER_41_1842 ();
 sg13g2_fill_2 FILLER_41_1849 ();
 sg13g2_fill_1 FILLER_41_1855 ();
 sg13g2_fill_2 FILLER_41_1865 ();
 sg13g2_fill_2 FILLER_41_1886 ();
 sg13g2_decap_4 FILLER_41_1894 ();
 sg13g2_fill_2 FILLER_41_1898 ();
 sg13g2_decap_8 FILLER_41_1904 ();
 sg13g2_decap_4 FILLER_41_1911 ();
 sg13g2_fill_2 FILLER_41_1919 ();
 sg13g2_fill_1 FILLER_41_1921 ();
 sg13g2_decap_4 FILLER_41_1931 ();
 sg13g2_fill_1 FILLER_41_1935 ();
 sg13g2_decap_4 FILLER_41_1945 ();
 sg13g2_decap_8 FILLER_41_1953 ();
 sg13g2_decap_4 FILLER_41_1960 ();
 sg13g2_fill_2 FILLER_41_1977 ();
 sg13g2_fill_1 FILLER_41_1979 ();
 sg13g2_decap_8 FILLER_41_1988 ();
 sg13g2_fill_2 FILLER_41_1995 ();
 sg13g2_fill_1 FILLER_41_1997 ();
 sg13g2_decap_8 FILLER_41_2003 ();
 sg13g2_decap_4 FILLER_41_2010 ();
 sg13g2_fill_2 FILLER_41_2023 ();
 sg13g2_fill_1 FILLER_41_2025 ();
 sg13g2_decap_4 FILLER_41_2030 ();
 sg13g2_fill_1 FILLER_41_2038 ();
 sg13g2_fill_2 FILLER_41_2043 ();
 sg13g2_fill_1 FILLER_41_2045 ();
 sg13g2_fill_1 FILLER_41_2050 ();
 sg13g2_decap_4 FILLER_41_2064 ();
 sg13g2_fill_1 FILLER_41_2068 ();
 sg13g2_fill_2 FILLER_41_2074 ();
 sg13g2_decap_8 FILLER_41_2080 ();
 sg13g2_decap_8 FILLER_41_2108 ();
 sg13g2_decap_8 FILLER_41_2115 ();
 sg13g2_fill_2 FILLER_41_2122 ();
 sg13g2_fill_1 FILLER_41_2124 ();
 sg13g2_decap_8 FILLER_41_2133 ();
 sg13g2_fill_2 FILLER_41_2140 ();
 sg13g2_decap_8 FILLER_41_2147 ();
 sg13g2_fill_1 FILLER_41_2154 ();
 sg13g2_decap_8 FILLER_41_2159 ();
 sg13g2_fill_1 FILLER_41_2166 ();
 sg13g2_decap_8 FILLER_41_2172 ();
 sg13g2_fill_1 FILLER_41_2179 ();
 sg13g2_fill_2 FILLER_41_2230 ();
 sg13g2_decap_4 FILLER_41_2258 ();
 sg13g2_fill_2 FILLER_41_2275 ();
 sg13g2_decap_8 FILLER_41_2281 ();
 sg13g2_decap_8 FILLER_41_2288 ();
 sg13g2_decap_8 FILLER_41_2295 ();
 sg13g2_decap_8 FILLER_41_2302 ();
 sg13g2_decap_4 FILLER_41_2309 ();
 sg13g2_fill_1 FILLER_41_2313 ();
 sg13g2_decap_8 FILLER_41_2333 ();
 sg13g2_fill_2 FILLER_41_2340 ();
 sg13g2_decap_8 FILLER_41_2361 ();
 sg13g2_decap_8 FILLER_41_2368 ();
 sg13g2_decap_8 FILLER_41_2375 ();
 sg13g2_fill_2 FILLER_41_2382 ();
 sg13g2_fill_1 FILLER_41_2384 ();
 sg13g2_decap_8 FILLER_41_2388 ();
 sg13g2_decap_8 FILLER_41_2395 ();
 sg13g2_decap_8 FILLER_41_2402 ();
 sg13g2_decap_8 FILLER_41_2409 ();
 sg13g2_decap_8 FILLER_41_2416 ();
 sg13g2_decap_8 FILLER_41_2423 ();
 sg13g2_decap_4 FILLER_41_2430 ();
 sg13g2_fill_2 FILLER_41_2434 ();
 sg13g2_decap_8 FILLER_41_2466 ();
 sg13g2_decap_4 FILLER_41_2473 ();
 sg13g2_fill_1 FILLER_41_2477 ();
 sg13g2_decap_8 FILLER_41_2513 ();
 sg13g2_fill_2 FILLER_41_2520 ();
 sg13g2_decap_4 FILLER_41_2528 ();
 sg13g2_decap_8 FILLER_41_2536 ();
 sg13g2_decap_8 FILLER_41_2543 ();
 sg13g2_decap_8 FILLER_41_2550 ();
 sg13g2_decap_8 FILLER_41_2557 ();
 sg13g2_decap_8 FILLER_41_2564 ();
 sg13g2_decap_8 FILLER_41_2571 ();
 sg13g2_decap_8 FILLER_41_2578 ();
 sg13g2_decap_8 FILLER_41_2585 ();
 sg13g2_decap_8 FILLER_41_2592 ();
 sg13g2_decap_8 FILLER_41_2599 ();
 sg13g2_decap_8 FILLER_41_2606 ();
 sg13g2_decap_8 FILLER_41_2613 ();
 sg13g2_decap_8 FILLER_41_2620 ();
 sg13g2_decap_8 FILLER_41_2627 ();
 sg13g2_decap_8 FILLER_41_2634 ();
 sg13g2_decap_8 FILLER_41_2641 ();
 sg13g2_decap_8 FILLER_41_2648 ();
 sg13g2_decap_8 FILLER_41_2655 ();
 sg13g2_decap_8 FILLER_41_2662 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_44 ();
 sg13g2_decap_4 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_55 ();
 sg13g2_decap_4 FILLER_42_68 ();
 sg13g2_fill_1 FILLER_42_72 ();
 sg13g2_decap_8 FILLER_42_103 ();
 sg13g2_decap_8 FILLER_42_110 ();
 sg13g2_decap_8 FILLER_42_117 ();
 sg13g2_decap_8 FILLER_42_124 ();
 sg13g2_decap_8 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_4 FILLER_42_182 ();
 sg13g2_decap_4 FILLER_42_189 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_fill_2 FILLER_42_226 ();
 sg13g2_decap_8 FILLER_42_233 ();
 sg13g2_decap_8 FILLER_42_240 ();
 sg13g2_decap_8 FILLER_42_247 ();
 sg13g2_decap_8 FILLER_42_254 ();
 sg13g2_decap_8 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_306 ();
 sg13g2_fill_1 FILLER_42_308 ();
 sg13g2_fill_2 FILLER_42_314 ();
 sg13g2_decap_8 FILLER_42_323 ();
 sg13g2_decap_8 FILLER_42_330 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_decap_8 FILLER_42_369 ();
 sg13g2_decap_8 FILLER_42_376 ();
 sg13g2_fill_2 FILLER_42_383 ();
 sg13g2_fill_1 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_419 ();
 sg13g2_decap_8 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_433 ();
 sg13g2_decap_8 FILLER_42_440 ();
 sg13g2_decap_8 FILLER_42_447 ();
 sg13g2_fill_2 FILLER_42_454 ();
 sg13g2_decap_8 FILLER_42_463 ();
 sg13g2_decap_4 FILLER_42_470 ();
 sg13g2_decap_4 FILLER_42_477 ();
 sg13g2_fill_1 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_506 ();
 sg13g2_decap_8 FILLER_42_513 ();
 sg13g2_fill_2 FILLER_42_520 ();
 sg13g2_fill_1 FILLER_42_522 ();
 sg13g2_decap_4 FILLER_42_527 ();
 sg13g2_fill_2 FILLER_42_540 ();
 sg13g2_fill_1 FILLER_42_542 ();
 sg13g2_decap_4 FILLER_42_547 ();
 sg13g2_fill_1 FILLER_42_551 ();
 sg13g2_decap_4 FILLER_42_557 ();
 sg13g2_fill_1 FILLER_42_561 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_fill_1 FILLER_42_574 ();
 sg13g2_fill_2 FILLER_42_583 ();
 sg13g2_fill_1 FILLER_42_607 ();
 sg13g2_fill_2 FILLER_42_614 ();
 sg13g2_fill_2 FILLER_42_621 ();
 sg13g2_fill_2 FILLER_42_634 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_fill_2 FILLER_42_721 ();
 sg13g2_decap_4 FILLER_42_727 ();
 sg13g2_fill_2 FILLER_42_731 ();
 sg13g2_decap_8 FILLER_42_737 ();
 sg13g2_decap_4 FILLER_42_744 ();
 sg13g2_fill_1 FILLER_42_748 ();
 sg13g2_decap_8 FILLER_42_755 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_4 FILLER_42_790 ();
 sg13g2_fill_2 FILLER_42_794 ();
 sg13g2_fill_2 FILLER_42_822 ();
 sg13g2_fill_1 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_864 ();
 sg13g2_decap_8 FILLER_42_871 ();
 sg13g2_decap_8 FILLER_42_878 ();
 sg13g2_decap_8 FILLER_42_885 ();
 sg13g2_decap_8 FILLER_42_892 ();
 sg13g2_fill_1 FILLER_42_899 ();
 sg13g2_decap_8 FILLER_42_905 ();
 sg13g2_decap_8 FILLER_42_912 ();
 sg13g2_decap_4 FILLER_42_919 ();
 sg13g2_fill_2 FILLER_42_923 ();
 sg13g2_decap_4 FILLER_42_956 ();
 sg13g2_fill_2 FILLER_42_970 ();
 sg13g2_decap_4 FILLER_42_981 ();
 sg13g2_fill_2 FILLER_42_985 ();
 sg13g2_decap_8 FILLER_42_996 ();
 sg13g2_decap_4 FILLER_42_1003 ();
 sg13g2_fill_2 FILLER_42_1007 ();
 sg13g2_fill_1 FILLER_42_1013 ();
 sg13g2_decap_8 FILLER_42_1018 ();
 sg13g2_decap_4 FILLER_42_1025 ();
 sg13g2_fill_1 FILLER_42_1029 ();
 sg13g2_decap_4 FILLER_42_1070 ();
 sg13g2_fill_1 FILLER_42_1074 ();
 sg13g2_fill_2 FILLER_42_1101 ();
 sg13g2_fill_1 FILLER_42_1103 ();
 sg13g2_fill_2 FILLER_42_1122 ();
 sg13g2_fill_2 FILLER_42_1128 ();
 sg13g2_fill_1 FILLER_42_1136 ();
 sg13g2_fill_1 FILLER_42_1143 ();
 sg13g2_fill_2 FILLER_42_1175 ();
 sg13g2_fill_1 FILLER_42_1186 ();
 sg13g2_fill_2 FILLER_42_1213 ();
 sg13g2_decap_8 FILLER_42_1219 ();
 sg13g2_fill_2 FILLER_42_1226 ();
 sg13g2_decap_4 FILLER_42_1254 ();
 sg13g2_fill_1 FILLER_42_1258 ();
 sg13g2_decap_4 FILLER_42_1290 ();
 sg13g2_fill_1 FILLER_42_1294 ();
 sg13g2_decap_8 FILLER_42_1303 ();
 sg13g2_decap_8 FILLER_42_1310 ();
 sg13g2_decap_4 FILLER_42_1317 ();
 sg13g2_fill_1 FILLER_42_1321 ();
 sg13g2_fill_1 FILLER_42_1327 ();
 sg13g2_fill_1 FILLER_42_1337 ();
 sg13g2_fill_2 FILLER_42_1343 ();
 sg13g2_fill_1 FILLER_42_1345 ();
 sg13g2_fill_2 FILLER_42_1350 ();
 sg13g2_fill_1 FILLER_42_1352 ();
 sg13g2_fill_2 FILLER_42_1361 ();
 sg13g2_decap_8 FILLER_42_1376 ();
 sg13g2_fill_1 FILLER_42_1394 ();
 sg13g2_fill_2 FILLER_42_1431 ();
 sg13g2_fill_2 FILLER_42_1454 ();
 sg13g2_fill_1 FILLER_42_1460 ();
 sg13g2_fill_2 FILLER_42_1469 ();
 sg13g2_fill_1 FILLER_42_1475 ();
 sg13g2_fill_1 FILLER_42_1490 ();
 sg13g2_decap_4 FILLER_42_1526 ();
 sg13g2_decap_4 FILLER_42_1535 ();
 sg13g2_fill_2 FILLER_42_1545 ();
 sg13g2_decap_4 FILLER_42_1552 ();
 sg13g2_fill_2 FILLER_42_1556 ();
 sg13g2_fill_2 FILLER_42_1576 ();
 sg13g2_decap_8 FILLER_42_1609 ();
 sg13g2_fill_2 FILLER_42_1616 ();
 sg13g2_fill_1 FILLER_42_1618 ();
 sg13g2_decap_8 FILLER_42_1645 ();
 sg13g2_decap_4 FILLER_42_1652 ();
 sg13g2_decap_8 FILLER_42_1713 ();
 sg13g2_decap_8 FILLER_42_1720 ();
 sg13g2_fill_2 FILLER_42_1727 ();
 sg13g2_decap_4 FILLER_42_1734 ();
 sg13g2_fill_2 FILLER_42_1747 ();
 sg13g2_fill_1 FILLER_42_1749 ();
 sg13g2_fill_2 FILLER_42_1754 ();
 sg13g2_decap_8 FILLER_42_1788 ();
 sg13g2_fill_1 FILLER_42_1795 ();
 sg13g2_fill_1 FILLER_42_1800 ();
 sg13g2_fill_1 FILLER_42_1832 ();
 sg13g2_decap_4 FILLER_42_1862 ();
 sg13g2_decap_8 FILLER_42_1897 ();
 sg13g2_decap_8 FILLER_42_1904 ();
 sg13g2_decap_8 FILLER_42_1916 ();
 sg13g2_fill_1 FILLER_42_1923 ();
 sg13g2_fill_1 FILLER_42_1933 ();
 sg13g2_fill_2 FILLER_42_1940 ();
 sg13g2_decap_8 FILLER_42_1957 ();
 sg13g2_fill_2 FILLER_42_1964 ();
 sg13g2_fill_1 FILLER_42_1966 ();
 sg13g2_decap_8 FILLER_42_1976 ();
 sg13g2_decap_8 FILLER_42_1983 ();
 sg13g2_decap_4 FILLER_42_1990 ();
 sg13g2_decap_8 FILLER_42_1999 ();
 sg13g2_decap_8 FILLER_42_2006 ();
 sg13g2_decap_8 FILLER_42_2013 ();
 sg13g2_decap_4 FILLER_42_2020 ();
 sg13g2_decap_8 FILLER_42_2034 ();
 sg13g2_decap_8 FILLER_42_2041 ();
 sg13g2_fill_2 FILLER_42_2056 ();
 sg13g2_fill_2 FILLER_42_2068 ();
 sg13g2_fill_1 FILLER_42_2070 ();
 sg13g2_decap_8 FILLER_42_2097 ();
 sg13g2_fill_2 FILLER_42_2104 ();
 sg13g2_decap_4 FILLER_42_2111 ();
 sg13g2_decap_8 FILLER_42_2120 ();
 sg13g2_decap_4 FILLER_42_2127 ();
 sg13g2_fill_1 FILLER_42_2141 ();
 sg13g2_fill_2 FILLER_42_2147 ();
 sg13g2_fill_1 FILLER_42_2149 ();
 sg13g2_fill_2 FILLER_42_2162 ();
 sg13g2_fill_1 FILLER_42_2164 ();
 sg13g2_decap_4 FILLER_42_2199 ();
 sg13g2_fill_2 FILLER_42_2203 ();
 sg13g2_decap_4 FILLER_42_2208 ();
 sg13g2_fill_1 FILLER_42_2212 ();
 sg13g2_fill_1 FILLER_42_2253 ();
 sg13g2_decap_8 FILLER_42_2280 ();
 sg13g2_decap_8 FILLER_42_2287 ();
 sg13g2_decap_8 FILLER_42_2294 ();
 sg13g2_fill_2 FILLER_42_2301 ();
 sg13g2_fill_1 FILLER_42_2303 ();
 sg13g2_fill_2 FILLER_42_2312 ();
 sg13g2_decap_8 FILLER_42_2318 ();
 sg13g2_decap_8 FILLER_42_2325 ();
 sg13g2_decap_4 FILLER_42_2332 ();
 sg13g2_fill_1 FILLER_42_2336 ();
 sg13g2_decap_8 FILLER_42_2398 ();
 sg13g2_decap_8 FILLER_42_2405 ();
 sg13g2_decap_8 FILLER_42_2412 ();
 sg13g2_decap_8 FILLER_42_2419 ();
 sg13g2_decap_4 FILLER_42_2426 ();
 sg13g2_fill_1 FILLER_42_2469 ();
 sg13g2_decap_8 FILLER_42_2500 ();
 sg13g2_decap_8 FILLER_42_2507 ();
 sg13g2_decap_8 FILLER_42_2514 ();
 sg13g2_decap_8 FILLER_42_2521 ();
 sg13g2_decap_8 FILLER_42_2528 ();
 sg13g2_decap_8 FILLER_42_2535 ();
 sg13g2_decap_8 FILLER_42_2542 ();
 sg13g2_decap_8 FILLER_42_2549 ();
 sg13g2_decap_8 FILLER_42_2556 ();
 sg13g2_decap_8 FILLER_42_2563 ();
 sg13g2_decap_8 FILLER_42_2570 ();
 sg13g2_decap_8 FILLER_42_2577 ();
 sg13g2_decap_8 FILLER_42_2584 ();
 sg13g2_decap_8 FILLER_42_2591 ();
 sg13g2_decap_8 FILLER_42_2598 ();
 sg13g2_decap_8 FILLER_42_2605 ();
 sg13g2_decap_8 FILLER_42_2612 ();
 sg13g2_decap_8 FILLER_42_2619 ();
 sg13g2_decap_8 FILLER_42_2626 ();
 sg13g2_decap_8 FILLER_42_2633 ();
 sg13g2_decap_8 FILLER_42_2640 ();
 sg13g2_decap_8 FILLER_42_2647 ();
 sg13g2_decap_8 FILLER_42_2654 ();
 sg13g2_decap_8 FILLER_42_2661 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_9 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_4 FILLER_43_49 ();
 sg13g2_decap_4 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_decap_8 FILLER_43_107 ();
 sg13g2_decap_8 FILLER_43_114 ();
 sg13g2_decap_8 FILLER_43_121 ();
 sg13g2_decap_4 FILLER_43_128 ();
 sg13g2_decap_8 FILLER_43_181 ();
 sg13g2_decap_8 FILLER_43_188 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_fill_2 FILLER_43_225 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_fill_2 FILLER_43_238 ();
 sg13g2_fill_1 FILLER_43_240 ();
 sg13g2_fill_1 FILLER_43_267 ();
 sg13g2_decap_8 FILLER_43_307 ();
 sg13g2_decap_8 FILLER_43_314 ();
 sg13g2_decap_4 FILLER_43_321 ();
 sg13g2_fill_1 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_decap_4 FILLER_43_360 ();
 sg13g2_fill_1 FILLER_43_364 ();
 sg13g2_fill_1 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_decap_4 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_415 ();
 sg13g2_decap_4 FILLER_43_426 ();
 sg13g2_fill_1 FILLER_43_430 ();
 sg13g2_fill_2 FILLER_43_495 ();
 sg13g2_fill_1 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_506 ();
 sg13g2_decap_4 FILLER_43_513 ();
 sg13g2_fill_2 FILLER_43_517 ();
 sg13g2_decap_4 FILLER_43_528 ();
 sg13g2_fill_1 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_decap_4 FILLER_43_569 ();
 sg13g2_fill_1 FILLER_43_573 ();
 sg13g2_fill_1 FILLER_43_604 ();
 sg13g2_decap_8 FILLER_43_627 ();
 sg13g2_decap_8 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_641 ();
 sg13g2_decap_4 FILLER_43_646 ();
 sg13g2_decap_8 FILLER_43_687 ();
 sg13g2_decap_8 FILLER_43_694 ();
 sg13g2_decap_4 FILLER_43_701 ();
 sg13g2_fill_1 FILLER_43_705 ();
 sg13g2_decap_8 FILLER_43_710 ();
 sg13g2_decap_8 FILLER_43_717 ();
 sg13g2_fill_2 FILLER_43_724 ();
 sg13g2_fill_2 FILLER_43_743 ();
 sg13g2_fill_1 FILLER_43_745 ();
 sg13g2_decap_8 FILLER_43_750 ();
 sg13g2_fill_2 FILLER_43_757 ();
 sg13g2_fill_1 FILLER_43_763 ();
 sg13g2_fill_1 FILLER_43_790 ();
 sg13g2_fill_1 FILLER_43_860 ();
 sg13g2_fill_2 FILLER_43_873 ();
 sg13g2_fill_1 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_885 ();
 sg13g2_decap_8 FILLER_43_892 ();
 sg13g2_decap_8 FILLER_43_899 ();
 sg13g2_decap_8 FILLER_43_906 ();
 sg13g2_decap_4 FILLER_43_913 ();
 sg13g2_fill_2 FILLER_43_917 ();
 sg13g2_fill_1 FILLER_43_932 ();
 sg13g2_decap_8 FILLER_43_937 ();
 sg13g2_fill_2 FILLER_43_944 ();
 sg13g2_fill_1 FILLER_43_946 ();
 sg13g2_fill_1 FILLER_43_983 ();
 sg13g2_fill_2 FILLER_43_988 ();
 sg13g2_decap_8 FILLER_43_999 ();
 sg13g2_fill_1 FILLER_43_1037 ();
 sg13g2_fill_2 FILLER_43_1074 ();
 sg13g2_decap_4 FILLER_43_1082 ();
 sg13g2_fill_2 FILLER_43_1086 ();
 sg13g2_decap_8 FILLER_43_1094 ();
 sg13g2_fill_1 FILLER_43_1101 ();
 sg13g2_fill_2 FILLER_43_1122 ();
 sg13g2_fill_1 FILLER_43_1124 ();
 sg13g2_fill_1 FILLER_43_1130 ();
 sg13g2_fill_2 FILLER_43_1140 ();
 sg13g2_decap_4 FILLER_43_1152 ();
 sg13g2_fill_2 FILLER_43_1162 ();
 sg13g2_fill_1 FILLER_43_1164 ();
 sg13g2_fill_1 FILLER_43_1180 ();
 sg13g2_decap_4 FILLER_43_1187 ();
 sg13g2_decap_8 FILLER_43_1196 ();
 sg13g2_decap_4 FILLER_43_1203 ();
 sg13g2_fill_1 FILLER_43_1212 ();
 sg13g2_fill_1 FILLER_43_1239 ();
 sg13g2_fill_2 FILLER_43_1266 ();
 sg13g2_decap_8 FILLER_43_1272 ();
 sg13g2_decap_8 FILLER_43_1279 ();
 sg13g2_fill_1 FILLER_43_1286 ();
 sg13g2_decap_4 FILLER_43_1291 ();
 sg13g2_fill_1 FILLER_43_1299 ();
 sg13g2_decap_8 FILLER_43_1310 ();
 sg13g2_decap_4 FILLER_43_1317 ();
 sg13g2_fill_1 FILLER_43_1321 ();
 sg13g2_fill_2 FILLER_43_1348 ();
 sg13g2_fill_1 FILLER_43_1385 ();
 sg13g2_fill_2 FILLER_43_1412 ();
 sg13g2_fill_2 FILLER_43_1425 ();
 sg13g2_fill_1 FILLER_43_1456 ();
 sg13g2_fill_2 FILLER_43_1462 ();
 sg13g2_fill_1 FILLER_43_1498 ();
 sg13g2_fill_2 FILLER_43_1525 ();
 sg13g2_fill_1 FILLER_43_1527 ();
 sg13g2_fill_2 FILLER_43_1542 ();
 sg13g2_fill_2 FILLER_43_1571 ();
 sg13g2_decap_8 FILLER_43_1610 ();
 sg13g2_decap_8 FILLER_43_1617 ();
 sg13g2_fill_2 FILLER_43_1624 ();
 sg13g2_decap_8 FILLER_43_1691 ();
 sg13g2_decap_8 FILLER_43_1698 ();
 sg13g2_decap_4 FILLER_43_1705 ();
 sg13g2_fill_1 FILLER_43_1769 ();
 sg13g2_decap_8 FILLER_43_1806 ();
 sg13g2_decap_8 FILLER_43_1813 ();
 sg13g2_fill_1 FILLER_43_1820 ();
 sg13g2_decap_4 FILLER_43_1825 ();
 sg13g2_decap_8 FILLER_43_1848 ();
 sg13g2_decap_8 FILLER_43_1855 ();
 sg13g2_decap_8 FILLER_43_1862 ();
 sg13g2_fill_2 FILLER_43_1869 ();
 sg13g2_fill_1 FILLER_43_1871 ();
 sg13g2_decap_8 FILLER_43_1876 ();
 sg13g2_decap_8 FILLER_43_1883 ();
 sg13g2_decap_8 FILLER_43_1890 ();
 sg13g2_decap_4 FILLER_43_1897 ();
 sg13g2_fill_1 FILLER_43_1905 ();
 sg13g2_fill_2 FILLER_43_1910 ();
 sg13g2_fill_1 FILLER_43_1912 ();
 sg13g2_fill_2 FILLER_43_1917 ();
 sg13g2_fill_1 FILLER_43_1948 ();
 sg13g2_fill_1 FILLER_43_1954 ();
 sg13g2_fill_2 FILLER_43_1960 ();
 sg13g2_fill_2 FILLER_43_1967 ();
 sg13g2_decap_8 FILLER_43_1995 ();
 sg13g2_decap_4 FILLER_43_2002 ();
 sg13g2_fill_1 FILLER_43_2006 ();
 sg13g2_decap_4 FILLER_43_2011 ();
 sg13g2_fill_1 FILLER_43_2015 ();
 sg13g2_decap_4 FILLER_43_2028 ();
 sg13g2_decap_4 FILLER_43_2037 ();
 sg13g2_fill_1 FILLER_43_2077 ();
 sg13g2_fill_2 FILLER_43_2108 ();
 sg13g2_fill_1 FILLER_43_2110 ();
 sg13g2_fill_2 FILLER_43_2141 ();
 sg13g2_fill_1 FILLER_43_2169 ();
 sg13g2_fill_2 FILLER_43_2215 ();
 sg13g2_fill_2 FILLER_43_2222 ();
 sg13g2_decap_4 FILLER_43_2294 ();
 sg13g2_fill_2 FILLER_43_2298 ();
 sg13g2_decap_4 FILLER_43_2304 ();
 sg13g2_fill_1 FILLER_43_2308 ();
 sg13g2_decap_8 FILLER_43_2335 ();
 sg13g2_fill_2 FILLER_43_2342 ();
 sg13g2_fill_1 FILLER_43_2344 ();
 sg13g2_fill_2 FILLER_43_2348 ();
 sg13g2_decap_8 FILLER_43_2354 ();
 sg13g2_fill_2 FILLER_43_2361 ();
 sg13g2_fill_1 FILLER_43_2363 ();
 sg13g2_fill_2 FILLER_43_2390 ();
 sg13g2_fill_2 FILLER_43_2418 ();
 sg13g2_fill_1 FILLER_43_2420 ();
 sg13g2_decap_8 FILLER_43_2451 ();
 sg13g2_decap_8 FILLER_43_2458 ();
 sg13g2_fill_2 FILLER_43_2475 ();
 sg13g2_decap_8 FILLER_43_2529 ();
 sg13g2_decap_8 FILLER_43_2536 ();
 sg13g2_decap_8 FILLER_43_2543 ();
 sg13g2_decap_8 FILLER_43_2550 ();
 sg13g2_decap_8 FILLER_43_2557 ();
 sg13g2_decap_8 FILLER_43_2564 ();
 sg13g2_decap_8 FILLER_43_2571 ();
 sg13g2_decap_8 FILLER_43_2578 ();
 sg13g2_decap_8 FILLER_43_2585 ();
 sg13g2_decap_8 FILLER_43_2592 ();
 sg13g2_decap_8 FILLER_43_2599 ();
 sg13g2_decap_8 FILLER_43_2606 ();
 sg13g2_decap_8 FILLER_43_2613 ();
 sg13g2_decap_8 FILLER_43_2620 ();
 sg13g2_decap_8 FILLER_43_2627 ();
 sg13g2_decap_8 FILLER_43_2634 ();
 sg13g2_decap_8 FILLER_43_2641 ();
 sg13g2_decap_8 FILLER_43_2648 ();
 sg13g2_decap_8 FILLER_43_2655 ();
 sg13g2_decap_8 FILLER_43_2662 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_8 ();
 sg13g2_fill_1 FILLER_44_10 ();
 sg13g2_fill_2 FILLER_44_19 ();
 sg13g2_fill_1 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_43 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_71 ();
 sg13g2_fill_2 FILLER_44_76 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_fill_2 FILLER_44_110 ();
 sg13g2_decap_8 FILLER_44_138 ();
 sg13g2_fill_2 FILLER_44_145 ();
 sg13g2_decap_8 FILLER_44_173 ();
 sg13g2_decap_8 FILLER_44_180 ();
 sg13g2_decap_8 FILLER_44_187 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_4 FILLER_44_208 ();
 sg13g2_fill_2 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_decap_8 FILLER_44_227 ();
 sg13g2_decap_8 FILLER_44_234 ();
 sg13g2_decap_4 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_fill_2 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_301 ();
 sg13g2_fill_2 FILLER_44_308 ();
 sg13g2_decap_4 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_324 ();
 sg13g2_decap_8 FILLER_44_331 ();
 sg13g2_decap_4 FILLER_44_338 ();
 sg13g2_fill_2 FILLER_44_342 ();
 sg13g2_fill_2 FILLER_44_348 ();
 sg13g2_fill_1 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_405 ();
 sg13g2_decap_8 FILLER_44_412 ();
 sg13g2_decap_8 FILLER_44_419 ();
 sg13g2_decap_8 FILLER_44_426 ();
 sg13g2_fill_1 FILLER_44_433 ();
 sg13g2_fill_2 FILLER_44_439 ();
 sg13g2_decap_4 FILLER_44_449 ();
 sg13g2_fill_2 FILLER_44_453 ();
 sg13g2_decap_8 FILLER_44_459 ();
 sg13g2_decap_8 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_473 ();
 sg13g2_fill_2 FILLER_44_480 ();
 sg13g2_fill_1 FILLER_44_482 ();
 sg13g2_fill_2 FILLER_44_500 ();
 sg13g2_decap_8 FILLER_44_512 ();
 sg13g2_fill_2 FILLER_44_519 ();
 sg13g2_decap_4 FILLER_44_530 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_decap_8 FILLER_44_564 ();
 sg13g2_decap_4 FILLER_44_571 ();
 sg13g2_fill_1 FILLER_44_575 ();
 sg13g2_fill_1 FILLER_44_581 ();
 sg13g2_fill_1 FILLER_44_594 ();
 sg13g2_fill_2 FILLER_44_600 ();
 sg13g2_fill_2 FILLER_44_606 ();
 sg13g2_fill_2 FILLER_44_612 ();
 sg13g2_decap_8 FILLER_44_622 ();
 sg13g2_decap_4 FILLER_44_629 ();
 sg13g2_fill_1 FILLER_44_633 ();
 sg13g2_fill_2 FILLER_44_639 ();
 sg13g2_fill_1 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_fill_2 FILLER_44_662 ();
 sg13g2_fill_1 FILLER_44_718 ();
 sg13g2_fill_2 FILLER_44_724 ();
 sg13g2_fill_1 FILLER_44_726 ();
 sg13g2_fill_2 FILLER_44_757 ();
 sg13g2_fill_1 FILLER_44_759 ();
 sg13g2_fill_1 FILLER_44_786 ();
 sg13g2_decap_4 FILLER_44_798 ();
 sg13g2_fill_1 FILLER_44_802 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_841 ();
 sg13g2_fill_2 FILLER_44_848 ();
 sg13g2_fill_2 FILLER_44_855 ();
 sg13g2_fill_2 FILLER_44_863 ();
 sg13g2_decap_4 FILLER_44_871 ();
 sg13g2_fill_1 FILLER_44_885 ();
 sg13g2_fill_1 FILLER_44_892 ();
 sg13g2_fill_1 FILLER_44_899 ();
 sg13g2_fill_2 FILLER_44_906 ();
 sg13g2_fill_1 FILLER_44_908 ();
 sg13g2_fill_1 FILLER_44_919 ();
 sg13g2_fill_2 FILLER_44_925 ();
 sg13g2_decap_8 FILLER_44_931 ();
 sg13g2_fill_2 FILLER_44_938 ();
 sg13g2_fill_1 FILLER_44_952 ();
 sg13g2_fill_2 FILLER_44_958 ();
 sg13g2_fill_1 FILLER_44_969 ();
 sg13g2_fill_2 FILLER_44_979 ();
 sg13g2_fill_1 FILLER_44_985 ();
 sg13g2_fill_2 FILLER_44_993 ();
 sg13g2_fill_1 FILLER_44_1019 ();
 sg13g2_decap_8 FILLER_44_1025 ();
 sg13g2_fill_1 FILLER_44_1032 ();
 sg13g2_fill_1 FILLER_44_1048 ();
 sg13g2_fill_1 FILLER_44_1067 ();
 sg13g2_fill_1 FILLER_44_1072 ();
 sg13g2_fill_1 FILLER_44_1102 ();
 sg13g2_fill_2 FILLER_44_1107 ();
 sg13g2_fill_1 FILLER_44_1109 ();
 sg13g2_decap_8 FILLER_44_1113 ();
 sg13g2_fill_2 FILLER_44_1120 ();
 sg13g2_fill_2 FILLER_44_1128 ();
 sg13g2_fill_1 FILLER_44_1130 ();
 sg13g2_decap_8 FILLER_44_1136 ();
 sg13g2_fill_1 FILLER_44_1143 ();
 sg13g2_decap_8 FILLER_44_1149 ();
 sg13g2_decap_8 FILLER_44_1156 ();
 sg13g2_decap_4 FILLER_44_1163 ();
 sg13g2_fill_1 FILLER_44_1167 ();
 sg13g2_decap_8 FILLER_44_1184 ();
 sg13g2_decap_4 FILLER_44_1191 ();
 sg13g2_fill_2 FILLER_44_1195 ();
 sg13g2_fill_1 FILLER_44_1202 ();
 sg13g2_decap_4 FILLER_44_1207 ();
 sg13g2_fill_2 FILLER_44_1211 ();
 sg13g2_decap_8 FILLER_44_1218 ();
 sg13g2_fill_2 FILLER_44_1225 ();
 sg13g2_fill_1 FILLER_44_1236 ();
 sg13g2_decap_8 FILLER_44_1263 ();
 sg13g2_decap_8 FILLER_44_1270 ();
 sg13g2_decap_4 FILLER_44_1277 ();
 sg13g2_decap_4 FILLER_44_1300 ();
 sg13g2_decap_8 FILLER_44_1309 ();
 sg13g2_decap_8 FILLER_44_1316 ();
 sg13g2_decap_8 FILLER_44_1323 ();
 sg13g2_fill_2 FILLER_44_1330 ();
 sg13g2_fill_1 FILLER_44_1332 ();
 sg13g2_fill_1 FILLER_44_1347 ();
 sg13g2_fill_1 FILLER_44_1364 ();
 sg13g2_decap_4 FILLER_44_1410 ();
 sg13g2_fill_2 FILLER_44_1428 ();
 sg13g2_fill_1 FILLER_44_1430 ();
 sg13g2_fill_1 FILLER_44_1450 ();
 sg13g2_decap_8 FILLER_44_1465 ();
 sg13g2_decap_8 FILLER_44_1472 ();
 sg13g2_fill_1 FILLER_44_1494 ();
 sg13g2_decap_4 FILLER_44_1507 ();
 sg13g2_fill_2 FILLER_44_1551 ();
 sg13g2_decap_4 FILLER_44_1624 ();
 sg13g2_fill_2 FILLER_44_1641 ();
 sg13g2_fill_1 FILLER_44_1643 ();
 sg13g2_decap_8 FILLER_44_1650 ();
 sg13g2_fill_2 FILLER_44_1657 ();
 sg13g2_decap_4 FILLER_44_1669 ();
 sg13g2_decap_8 FILLER_44_1686 ();
 sg13g2_decap_4 FILLER_44_1693 ();
 sg13g2_fill_2 FILLER_44_1697 ();
 sg13g2_decap_4 FILLER_44_1714 ();
 sg13g2_fill_2 FILLER_44_1718 ();
 sg13g2_fill_2 FILLER_44_1769 ();
 sg13g2_fill_1 FILLER_44_1771 ();
 sg13g2_decap_8 FILLER_44_1803 ();
 sg13g2_decap_4 FILLER_44_1810 ();
 sg13g2_fill_2 FILLER_44_1814 ();
 sg13g2_fill_2 FILLER_44_1822 ();
 sg13g2_fill_2 FILLER_44_1829 ();
 sg13g2_fill_1 FILLER_44_1831 ();
 sg13g2_decap_4 FILLER_44_1860 ();
 sg13g2_fill_1 FILLER_44_1864 ();
 sg13g2_fill_1 FILLER_44_1933 ();
 sg13g2_fill_1 FILLER_44_1939 ();
 sg13g2_fill_1 FILLER_44_1972 ();
 sg13g2_decap_4 FILLER_44_1983 ();
 sg13g2_fill_1 FILLER_44_2017 ();
 sg13g2_fill_2 FILLER_44_2069 ();
 sg13g2_fill_1 FILLER_44_2071 ();
 sg13g2_fill_1 FILLER_44_2077 ();
 sg13g2_fill_1 FILLER_44_2082 ();
 sg13g2_decap_8 FILLER_44_2089 ();
 sg13g2_fill_1 FILLER_44_2096 ();
 sg13g2_decap_8 FILLER_44_2105 ();
 sg13g2_decap_4 FILLER_44_2112 ();
 sg13g2_fill_1 FILLER_44_2116 ();
 sg13g2_decap_4 FILLER_44_2129 ();
 sg13g2_fill_2 FILLER_44_2133 ();
 sg13g2_decap_4 FILLER_44_2140 ();
 sg13g2_fill_2 FILLER_44_2144 ();
 sg13g2_decap_8 FILLER_44_2150 ();
 sg13g2_fill_1 FILLER_44_2196 ();
 sg13g2_fill_2 FILLER_44_2234 ();
 sg13g2_fill_1 FILLER_44_2241 ();
 sg13g2_fill_2 FILLER_44_2246 ();
 sg13g2_fill_2 FILLER_44_2254 ();
 sg13g2_fill_2 FILLER_44_2262 ();
 sg13g2_fill_2 FILLER_44_2268 ();
 sg13g2_fill_1 FILLER_44_2270 ();
 sg13g2_fill_1 FILLER_44_2280 ();
 sg13g2_fill_2 FILLER_44_2286 ();
 sg13g2_fill_2 FILLER_44_2297 ();
 sg13g2_fill_2 FILLER_44_2304 ();
 sg13g2_decap_4 FILLER_44_2332 ();
 sg13g2_fill_1 FILLER_44_2375 ();
 sg13g2_fill_2 FILLER_44_2380 ();
 sg13g2_decap_4 FILLER_44_2386 ();
 sg13g2_decap_8 FILLER_44_2395 ();
 sg13g2_decap_8 FILLER_44_2402 ();
 sg13g2_decap_8 FILLER_44_2409 ();
 sg13g2_decap_8 FILLER_44_2416 ();
 sg13g2_decap_8 FILLER_44_2423 ();
 sg13g2_fill_1 FILLER_44_2439 ();
 sg13g2_fill_1 FILLER_44_2445 ();
 sg13g2_decap_8 FILLER_44_2452 ();
 sg13g2_decap_4 FILLER_44_2459 ();
 sg13g2_fill_1 FILLER_44_2463 ();
 sg13g2_fill_2 FILLER_44_2470 ();
 sg13g2_decap_4 FILLER_44_2497 ();
 sg13g2_fill_1 FILLER_44_2501 ();
 sg13g2_fill_2 FILLER_44_2506 ();
 sg13g2_fill_1 FILLER_44_2508 ();
 sg13g2_decap_8 FILLER_44_2513 ();
 sg13g2_decap_8 FILLER_44_2550 ();
 sg13g2_decap_8 FILLER_44_2557 ();
 sg13g2_decap_8 FILLER_44_2564 ();
 sg13g2_decap_8 FILLER_44_2571 ();
 sg13g2_decap_8 FILLER_44_2578 ();
 sg13g2_decap_8 FILLER_44_2585 ();
 sg13g2_decap_8 FILLER_44_2592 ();
 sg13g2_decap_8 FILLER_44_2599 ();
 sg13g2_decap_8 FILLER_44_2606 ();
 sg13g2_decap_8 FILLER_44_2613 ();
 sg13g2_decap_8 FILLER_44_2620 ();
 sg13g2_decap_8 FILLER_44_2627 ();
 sg13g2_decap_8 FILLER_44_2634 ();
 sg13g2_decap_8 FILLER_44_2641 ();
 sg13g2_decap_8 FILLER_44_2648 ();
 sg13g2_decap_8 FILLER_44_2655 ();
 sg13g2_decap_8 FILLER_44_2662 ();
 sg13g2_fill_1 FILLER_44_2669 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_1 FILLER_45_38 ();
 sg13g2_fill_2 FILLER_45_45 ();
 sg13g2_fill_1 FILLER_45_52 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_86 ();
 sg13g2_decap_8 FILLER_45_93 ();
 sg13g2_decap_8 FILLER_45_100 ();
 sg13g2_decap_8 FILLER_45_107 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_1 FILLER_45_200 ();
 sg13g2_fill_2 FILLER_45_209 ();
 sg13g2_fill_1 FILLER_45_216 ();
 sg13g2_decap_8 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_233 ();
 sg13g2_decap_8 FILLER_45_240 ();
 sg13g2_decap_8 FILLER_45_247 ();
 sg13g2_decap_8 FILLER_45_254 ();
 sg13g2_decap_8 FILLER_45_261 ();
 sg13g2_decap_8 FILLER_45_268 ();
 sg13g2_decap_4 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_279 ();
 sg13g2_decap_4 FILLER_45_285 ();
 sg13g2_fill_1 FILLER_45_289 ();
 sg13g2_fill_2 FILLER_45_299 ();
 sg13g2_fill_1 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_decap_8 FILLER_45_327 ();
 sg13g2_decap_4 FILLER_45_334 ();
 sg13g2_fill_2 FILLER_45_338 ();
 sg13g2_fill_2 FILLER_45_354 ();
 sg13g2_decap_4 FILLER_45_359 ();
 sg13g2_fill_1 FILLER_45_363 ();
 sg13g2_fill_1 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_4 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_400 ();
 sg13g2_decap_4 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_45_415 ();
 sg13g2_decap_4 FILLER_45_422 ();
 sg13g2_fill_2 FILLER_45_426 ();
 sg13g2_fill_2 FILLER_45_434 ();
 sg13g2_fill_1 FILLER_45_436 ();
 sg13g2_decap_8 FILLER_45_456 ();
 sg13g2_decap_8 FILLER_45_463 ();
 sg13g2_decap_8 FILLER_45_470 ();
 sg13g2_decap_4 FILLER_45_477 ();
 sg13g2_fill_1 FILLER_45_481 ();
 sg13g2_decap_8 FILLER_45_492 ();
 sg13g2_fill_1 FILLER_45_499 ();
 sg13g2_fill_1 FILLER_45_510 ();
 sg13g2_fill_2 FILLER_45_521 ();
 sg13g2_fill_2 FILLER_45_528 ();
 sg13g2_decap_4 FILLER_45_552 ();
 sg13g2_fill_2 FILLER_45_556 ();
 sg13g2_fill_2 FILLER_45_563 ();
 sg13g2_decap_4 FILLER_45_570 ();
 sg13g2_fill_1 FILLER_45_574 ();
 sg13g2_fill_1 FILLER_45_580 ();
 sg13g2_fill_1 FILLER_45_586 ();
 sg13g2_decap_8 FILLER_45_606 ();
 sg13g2_decap_8 FILLER_45_613 ();
 sg13g2_decap_8 FILLER_45_628 ();
 sg13g2_decap_8 FILLER_45_635 ();
 sg13g2_decap_8 FILLER_45_642 ();
 sg13g2_decap_8 FILLER_45_649 ();
 sg13g2_decap_8 FILLER_45_656 ();
 sg13g2_decap_8 FILLER_45_663 ();
 sg13g2_decap_8 FILLER_45_670 ();
 sg13g2_decap_8 FILLER_45_677 ();
 sg13g2_decap_8 FILLER_45_684 ();
 sg13g2_decap_4 FILLER_45_691 ();
 sg13g2_fill_2 FILLER_45_700 ();
 sg13g2_fill_1 FILLER_45_702 ();
 sg13g2_decap_4 FILLER_45_734 ();
 sg13g2_fill_1 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_fill_1 FILLER_45_809 ();
 sg13g2_fill_2 FILLER_45_820 ();
 sg13g2_fill_1 FILLER_45_822 ();
 sg13g2_decap_4 FILLER_45_827 ();
 sg13g2_decap_8 FILLER_45_836 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_4 FILLER_45_868 ();
 sg13g2_fill_2 FILLER_45_872 ();
 sg13g2_decap_8 FILLER_45_880 ();
 sg13g2_fill_1 FILLER_45_887 ();
 sg13g2_fill_2 FILLER_45_894 ();
 sg13g2_fill_1 FILLER_45_911 ();
 sg13g2_decap_4 FILLER_45_919 ();
 sg13g2_fill_1 FILLER_45_923 ();
 sg13g2_fill_2 FILLER_45_965 ();
 sg13g2_fill_1 FILLER_45_967 ();
 sg13g2_decap_4 FILLER_45_977 ();
 sg13g2_fill_1 FILLER_45_992 ();
 sg13g2_decap_8 FILLER_45_1013 ();
 sg13g2_decap_8 FILLER_45_1020 ();
 sg13g2_decap_8 FILLER_45_1027 ();
 sg13g2_decap_4 FILLER_45_1034 ();
 sg13g2_fill_1 FILLER_45_1038 ();
 sg13g2_fill_2 FILLER_45_1043 ();
 sg13g2_decap_4 FILLER_45_1067 ();
 sg13g2_fill_1 FILLER_45_1071 ();
 sg13g2_decap_8 FILLER_45_1076 ();
 sg13g2_fill_1 FILLER_45_1098 ();
 sg13g2_fill_2 FILLER_45_1103 ();
 sg13g2_fill_1 FILLER_45_1109 ();
 sg13g2_fill_2 FILLER_45_1121 ();
 sg13g2_decap_8 FILLER_45_1134 ();
 sg13g2_decap_4 FILLER_45_1141 ();
 sg13g2_fill_1 FILLER_45_1145 ();
 sg13g2_decap_4 FILLER_45_1172 ();
 sg13g2_fill_2 FILLER_45_1176 ();
 sg13g2_decap_8 FILLER_45_1187 ();
 sg13g2_decap_8 FILLER_45_1225 ();
 sg13g2_decap_8 FILLER_45_1232 ();
 sg13g2_decap_4 FILLER_45_1245 ();
 sg13g2_decap_8 FILLER_45_1254 ();
 sg13g2_decap_8 FILLER_45_1261 ();
 sg13g2_decap_8 FILLER_45_1268 ();
 sg13g2_decap_8 FILLER_45_1275 ();
 sg13g2_decap_4 FILLER_45_1282 ();
 sg13g2_decap_4 FILLER_45_1291 ();
 sg13g2_fill_2 FILLER_45_1299 ();
 sg13g2_decap_8 FILLER_45_1307 ();
 sg13g2_decap_8 FILLER_45_1314 ();
 sg13g2_fill_2 FILLER_45_1321 ();
 sg13g2_fill_1 FILLER_45_1323 ();
 sg13g2_fill_2 FILLER_45_1364 ();
 sg13g2_fill_1 FILLER_45_1374 ();
 sg13g2_fill_2 FILLER_45_1394 ();
 sg13g2_fill_1 FILLER_45_1407 ();
 sg13g2_fill_2 FILLER_45_1412 ();
 sg13g2_fill_2 FILLER_45_1418 ();
 sg13g2_fill_2 FILLER_45_1424 ();
 sg13g2_fill_2 FILLER_45_1439 ();
 sg13g2_decap_8 FILLER_45_1446 ();
 sg13g2_decap_8 FILLER_45_1453 ();
 sg13g2_decap_4 FILLER_45_1460 ();
 sg13g2_decap_8 FILLER_45_1473 ();
 sg13g2_decap_8 FILLER_45_1480 ();
 sg13g2_decap_4 FILLER_45_1502 ();
 sg13g2_fill_2 FILLER_45_1506 ();
 sg13g2_decap_8 FILLER_45_1538 ();
 sg13g2_fill_2 FILLER_45_1545 ();
 sg13g2_fill_1 FILLER_45_1547 ();
 sg13g2_fill_2 FILLER_45_1559 ();
 sg13g2_fill_1 FILLER_45_1566 ();
 sg13g2_decap_8 FILLER_45_1572 ();
 sg13g2_decap_4 FILLER_45_1579 ();
 sg13g2_fill_1 FILLER_45_1588 ();
 sg13g2_fill_2 FILLER_45_1594 ();
 sg13g2_fill_1 FILLER_45_1596 ();
 sg13g2_fill_1 FILLER_45_1607 ();
 sg13g2_decap_8 FILLER_45_1612 ();
 sg13g2_decap_4 FILLER_45_1619 ();
 sg13g2_fill_2 FILLER_45_1623 ();
 sg13g2_decap_8 FILLER_45_1639 ();
 sg13g2_decap_8 FILLER_45_1646 ();
 sg13g2_decap_8 FILLER_45_1653 ();
 sg13g2_decap_4 FILLER_45_1660 ();
 sg13g2_decap_8 FILLER_45_1690 ();
 sg13g2_fill_2 FILLER_45_1697 ();
 sg13g2_decap_8 FILLER_45_1711 ();
 sg13g2_decap_8 FILLER_45_1718 ();
 sg13g2_decap_8 FILLER_45_1725 ();
 sg13g2_decap_8 FILLER_45_1732 ();
 sg13g2_decap_8 FILLER_45_1739 ();
 sg13g2_decap_8 FILLER_45_1746 ();
 sg13g2_fill_1 FILLER_45_1753 ();
 sg13g2_decap_8 FILLER_45_1776 ();
 sg13g2_fill_1 FILLER_45_1783 ();
 sg13g2_decap_4 FILLER_45_1788 ();
 sg13g2_fill_2 FILLER_45_1792 ();
 sg13g2_fill_1 FILLER_45_1805 ();
 sg13g2_decap_8 FILLER_45_1810 ();
 sg13g2_fill_1 FILLER_45_1939 ();
 sg13g2_fill_2 FILLER_45_1972 ();
 sg13g2_decap_8 FILLER_45_1979 ();
 sg13g2_decap_8 FILLER_45_1995 ();
 sg13g2_decap_8 FILLER_45_2002 ();
 sg13g2_decap_8 FILLER_45_2009 ();
 sg13g2_decap_8 FILLER_45_2016 ();
 sg13g2_fill_1 FILLER_45_2023 ();
 sg13g2_fill_1 FILLER_45_2041 ();
 sg13g2_decap_4 FILLER_45_2056 ();
 sg13g2_fill_2 FILLER_45_2060 ();
 sg13g2_decap_4 FILLER_45_2066 ();
 sg13g2_decap_4 FILLER_45_2074 ();
 sg13g2_fill_2 FILLER_45_2078 ();
 sg13g2_decap_8 FILLER_45_2084 ();
 sg13g2_decap_8 FILLER_45_2091 ();
 sg13g2_decap_8 FILLER_45_2098 ();
 sg13g2_fill_2 FILLER_45_2105 ();
 sg13g2_decap_4 FILLER_45_2111 ();
 sg13g2_fill_2 FILLER_45_2120 ();
 sg13g2_fill_1 FILLER_45_2122 ();
 sg13g2_fill_2 FILLER_45_2127 ();
 sg13g2_decap_4 FILLER_45_2160 ();
 sg13g2_fill_1 FILLER_45_2164 ();
 sg13g2_decap_8 FILLER_45_2170 ();
 sg13g2_decap_4 FILLER_45_2177 ();
 sg13g2_fill_1 FILLER_45_2186 ();
 sg13g2_decap_4 FILLER_45_2202 ();
 sg13g2_decap_8 FILLER_45_2211 ();
 sg13g2_fill_1 FILLER_45_2218 ();
 sg13g2_fill_1 FILLER_45_2245 ();
 sg13g2_decap_8 FILLER_45_2251 ();
 sg13g2_decap_8 FILLER_45_2258 ();
 sg13g2_decap_8 FILLER_45_2265 ();
 sg13g2_decap_4 FILLER_45_2298 ();
 sg13g2_decap_4 FILLER_45_2308 ();
 sg13g2_fill_1 FILLER_45_2312 ();
 sg13g2_fill_2 FILLER_45_2319 ();
 sg13g2_decap_8 FILLER_45_2330 ();
 sg13g2_decap_8 FILLER_45_2337 ();
 sg13g2_fill_2 FILLER_45_2344 ();
 sg13g2_decap_8 FILLER_45_2401 ();
 sg13g2_fill_2 FILLER_45_2408 ();
 sg13g2_fill_2 FILLER_45_2419 ();
 sg13g2_fill_2 FILLER_45_2458 ();
 sg13g2_fill_1 FILLER_45_2464 ();
 sg13g2_fill_2 FILLER_45_2473 ();
 sg13g2_fill_1 FILLER_45_2490 ();
 sg13g2_fill_2 FILLER_45_2529 ();
 sg13g2_decap_8 FILLER_45_2535 ();
 sg13g2_decap_8 FILLER_45_2542 ();
 sg13g2_decap_8 FILLER_45_2549 ();
 sg13g2_decap_8 FILLER_45_2556 ();
 sg13g2_decap_8 FILLER_45_2563 ();
 sg13g2_decap_8 FILLER_45_2570 ();
 sg13g2_decap_8 FILLER_45_2577 ();
 sg13g2_decap_8 FILLER_45_2584 ();
 sg13g2_decap_8 FILLER_45_2591 ();
 sg13g2_decap_8 FILLER_45_2598 ();
 sg13g2_decap_8 FILLER_45_2605 ();
 sg13g2_decap_8 FILLER_45_2612 ();
 sg13g2_decap_8 FILLER_45_2619 ();
 sg13g2_decap_8 FILLER_45_2626 ();
 sg13g2_decap_8 FILLER_45_2633 ();
 sg13g2_decap_8 FILLER_45_2640 ();
 sg13g2_decap_8 FILLER_45_2647 ();
 sg13g2_decap_8 FILLER_45_2654 ();
 sg13g2_decap_8 FILLER_45_2661 ();
 sg13g2_fill_2 FILLER_45_2668 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_16 ();
 sg13g2_fill_1 FILLER_46_33 ();
 sg13g2_fill_1 FILLER_46_73 ();
 sg13g2_decap_8 FILLER_46_79 ();
 sg13g2_decap_8 FILLER_46_86 ();
 sg13g2_decap_8 FILLER_46_93 ();
 sg13g2_decap_4 FILLER_46_100 ();
 sg13g2_fill_1 FILLER_46_104 ();
 sg13g2_decap_8 FILLER_46_121 ();
 sg13g2_decap_4 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_fill_1 FILLER_46_142 ();
 sg13g2_decap_8 FILLER_46_151 ();
 sg13g2_decap_8 FILLER_46_158 ();
 sg13g2_fill_2 FILLER_46_165 ();
 sg13g2_decap_8 FILLER_46_170 ();
 sg13g2_decap_8 FILLER_46_177 ();
 sg13g2_fill_2 FILLER_46_184 ();
 sg13g2_fill_2 FILLER_46_225 ();
 sg13g2_decap_8 FILLER_46_241 ();
 sg13g2_decap_8 FILLER_46_248 ();
 sg13g2_fill_2 FILLER_46_255 ();
 sg13g2_fill_1 FILLER_46_257 ();
 sg13g2_decap_4 FILLER_46_291 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_372 ();
 sg13g2_decap_4 FILLER_46_379 ();
 sg13g2_fill_1 FILLER_46_383 ();
 sg13g2_decap_4 FILLER_46_389 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_1 FILLER_46_402 ();
 sg13g2_fill_1 FILLER_46_411 ();
 sg13g2_fill_1 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_46_453 ();
 sg13g2_decap_8 FILLER_46_460 ();
 sg13g2_decap_8 FILLER_46_467 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_decap_8 FILLER_46_495 ();
 sg13g2_fill_2 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_558 ();
 sg13g2_decap_8 FILLER_46_606 ();
 sg13g2_decap_8 FILLER_46_613 ();
 sg13g2_decap_8 FILLER_46_620 ();
 sg13g2_decap_8 FILLER_46_627 ();
 sg13g2_decap_8 FILLER_46_634 ();
 sg13g2_decap_8 FILLER_46_641 ();
 sg13g2_decap_8 FILLER_46_648 ();
 sg13g2_decap_8 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_662 ();
 sg13g2_fill_2 FILLER_46_668 ();
 sg13g2_decap_8 FILLER_46_683 ();
 sg13g2_fill_2 FILLER_46_690 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_4 FILLER_46_707 ();
 sg13g2_fill_1 FILLER_46_711 ();
 sg13g2_fill_2 FILLER_46_756 ();
 sg13g2_fill_2 FILLER_46_764 ();
 sg13g2_fill_2 FILLER_46_783 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_4 FILLER_46_822 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_4 FILLER_46_883 ();
 sg13g2_fill_2 FILLER_46_897 ();
 sg13g2_decap_4 FILLER_46_920 ();
 sg13g2_fill_1 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_929 ();
 sg13g2_fill_1 FILLER_46_936 ();
 sg13g2_decap_8 FILLER_46_941 ();
 sg13g2_fill_2 FILLER_46_948 ();
 sg13g2_fill_2 FILLER_46_968 ();
 sg13g2_fill_1 FILLER_46_970 ();
 sg13g2_decap_4 FILLER_46_981 ();
 sg13g2_fill_2 FILLER_46_985 ();
 sg13g2_fill_2 FILLER_46_1008 ();
 sg13g2_fill_2 FILLER_46_1014 ();
 sg13g2_fill_1 FILLER_46_1016 ();
 sg13g2_fill_1 FILLER_46_1021 ();
 sg13g2_fill_1 FILLER_46_1027 ();
 sg13g2_fill_2 FILLER_46_1037 ();
 sg13g2_decap_8 FILLER_46_1050 ();
 sg13g2_fill_1 FILLER_46_1066 ();
 sg13g2_decap_8 FILLER_46_1104 ();
 sg13g2_decap_8 FILLER_46_1111 ();
 sg13g2_fill_2 FILLER_46_1118 ();
 sg13g2_decap_8 FILLER_46_1128 ();
 sg13g2_decap_8 FILLER_46_1135 ();
 sg13g2_fill_2 FILLER_46_1142 ();
 sg13g2_decap_8 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1155 ();
 sg13g2_fill_1 FILLER_46_1162 ();
 sg13g2_fill_2 FILLER_46_1176 ();
 sg13g2_fill_1 FILLER_46_1178 ();
 sg13g2_decap_4 FILLER_46_1188 ();
 sg13g2_fill_2 FILLER_46_1222 ();
 sg13g2_fill_1 FILLER_46_1224 ();
 sg13g2_fill_1 FILLER_46_1251 ();
 sg13g2_fill_1 FILLER_46_1270 ();
 sg13g2_fill_2 FILLER_46_1287 ();
 sg13g2_fill_1 FILLER_46_1289 ();
 sg13g2_fill_1 FILLER_46_1294 ();
 sg13g2_decap_8 FILLER_46_1307 ();
 sg13g2_decap_8 FILLER_46_1314 ();
 sg13g2_decap_8 FILLER_46_1321 ();
 sg13g2_fill_2 FILLER_46_1328 ();
 sg13g2_fill_1 FILLER_46_1359 ();
 sg13g2_decap_8 FILLER_46_1411 ();
 sg13g2_decap_8 FILLER_46_1440 ();
 sg13g2_fill_2 FILLER_46_1447 ();
 sg13g2_fill_1 FILLER_46_1459 ();
 sg13g2_fill_2 FILLER_46_1464 ();
 sg13g2_fill_2 FILLER_46_1501 ();
 sg13g2_fill_1 FILLER_46_1503 ();
 sg13g2_decap_8 FILLER_46_1509 ();
 sg13g2_decap_4 FILLER_46_1516 ();
 sg13g2_decap_8 FILLER_46_1531 ();
 sg13g2_decap_8 FILLER_46_1538 ();
 sg13g2_decap_8 FILLER_46_1545 ();
 sg13g2_decap_4 FILLER_46_1552 ();
 sg13g2_fill_1 FILLER_46_1559 ();
 sg13g2_fill_1 FILLER_46_1567 ();
 sg13g2_decap_8 FILLER_46_1573 ();
 sg13g2_decap_4 FILLER_46_1580 ();
 sg13g2_fill_1 FILLER_46_1599 ();
 sg13g2_decap_4 FILLER_46_1605 ();
 sg13g2_fill_2 FILLER_46_1609 ();
 sg13g2_fill_2 FILLER_46_1637 ();
 sg13g2_fill_2 FILLER_46_1642 ();
 sg13g2_fill_1 FILLER_46_1644 ();
 sg13g2_fill_1 FILLER_46_1650 ();
 sg13g2_decap_8 FILLER_46_1660 ();
 sg13g2_decap_4 FILLER_46_1667 ();
 sg13g2_fill_1 FILLER_46_1671 ();
 sg13g2_fill_1 FILLER_46_1677 ();
 sg13g2_decap_4 FILLER_46_1704 ();
 sg13g2_fill_1 FILLER_46_1713 ();
 sg13g2_fill_1 FILLER_46_1719 ();
 sg13g2_decap_8 FILLER_46_1729 ();
 sg13g2_decap_8 FILLER_46_1736 ();
 sg13g2_decap_8 FILLER_46_1743 ();
 sg13g2_decap_8 FILLER_46_1750 ();
 sg13g2_decap_8 FILLER_46_1757 ();
 sg13g2_decap_8 FILLER_46_1764 ();
 sg13g2_decap_8 FILLER_46_1771 ();
 sg13g2_decap_8 FILLER_46_1778 ();
 sg13g2_decap_8 FILLER_46_1785 ();
 sg13g2_decap_4 FILLER_46_1792 ();
 sg13g2_decap_8 FILLER_46_1822 ();
 sg13g2_fill_2 FILLER_46_1829 ();
 sg13g2_fill_1 FILLER_46_1831 ();
 sg13g2_fill_1 FILLER_46_1836 ();
 sg13g2_fill_2 FILLER_46_1843 ();
 sg13g2_decap_8 FILLER_46_1875 ();
 sg13g2_decap_8 FILLER_46_1882 ();
 sg13g2_decap_8 FILLER_46_1889 ();
 sg13g2_decap_8 FILLER_46_1896 ();
 sg13g2_fill_1 FILLER_46_1903 ();
 sg13g2_fill_1 FILLER_46_1917 ();
 sg13g2_fill_1 FILLER_46_1924 ();
 sg13g2_fill_1 FILLER_46_1943 ();
 sg13g2_decap_8 FILLER_46_1986 ();
 sg13g2_decap_4 FILLER_46_1993 ();
 sg13g2_decap_4 FILLER_46_2014 ();
 sg13g2_fill_2 FILLER_46_2018 ();
 sg13g2_decap_4 FILLER_46_2028 ();
 sg13g2_fill_1 FILLER_46_2032 ();
 sg13g2_fill_2 FILLER_46_2037 ();
 sg13g2_fill_1 FILLER_46_2039 ();
 sg13g2_decap_8 FILLER_46_2045 ();
 sg13g2_fill_2 FILLER_46_2052 ();
 sg13g2_decap_4 FILLER_46_2063 ();
 sg13g2_fill_1 FILLER_46_2067 ();
 sg13g2_decap_4 FILLER_46_2082 ();
 sg13g2_fill_2 FILLER_46_2090 ();
 sg13g2_decap_4 FILLER_46_2097 ();
 sg13g2_fill_1 FILLER_46_2105 ();
 sg13g2_fill_1 FILLER_46_2150 ();
 sg13g2_decap_4 FILLER_46_2156 ();
 sg13g2_fill_1 FILLER_46_2160 ();
 sg13g2_fill_2 FILLER_46_2191 ();
 sg13g2_decap_4 FILLER_46_2198 ();
 sg13g2_decap_4 FILLER_46_2206 ();
 sg13g2_fill_2 FILLER_46_2210 ();
 sg13g2_decap_4 FILLER_46_2216 ();
 sg13g2_fill_1 FILLER_46_2220 ();
 sg13g2_decap_8 FILLER_46_2230 ();
 sg13g2_fill_2 FILLER_46_2237 ();
 sg13g2_fill_1 FILLER_46_2239 ();
 sg13g2_fill_1 FILLER_46_2246 ();
 sg13g2_decap_4 FILLER_46_2251 ();
 sg13g2_fill_1 FILLER_46_2255 ();
 sg13g2_decap_4 FILLER_46_2260 ();
 sg13g2_fill_2 FILLER_46_2275 ();
 sg13g2_fill_1 FILLER_46_2277 ();
 sg13g2_fill_2 FILLER_46_2282 ();
 sg13g2_decap_4 FILLER_46_2288 ();
 sg13g2_fill_2 FILLER_46_2292 ();
 sg13g2_fill_2 FILLER_46_2352 ();
 sg13g2_decap_8 FILLER_46_2385 ();
 sg13g2_decap_8 FILLER_46_2392 ();
 sg13g2_fill_1 FILLER_46_2403 ();
 sg13g2_fill_2 FILLER_46_2463 ();
 sg13g2_decap_4 FILLER_46_2470 ();
 sg13g2_fill_1 FILLER_46_2474 ();
 sg13g2_decap_8 FILLER_46_2548 ();
 sg13g2_decap_8 FILLER_46_2555 ();
 sg13g2_decap_8 FILLER_46_2562 ();
 sg13g2_decap_8 FILLER_46_2569 ();
 sg13g2_decap_8 FILLER_46_2576 ();
 sg13g2_decap_8 FILLER_46_2583 ();
 sg13g2_decap_8 FILLER_46_2590 ();
 sg13g2_decap_8 FILLER_46_2597 ();
 sg13g2_decap_8 FILLER_46_2604 ();
 sg13g2_decap_8 FILLER_46_2611 ();
 sg13g2_decap_8 FILLER_46_2618 ();
 sg13g2_decap_8 FILLER_46_2625 ();
 sg13g2_decap_8 FILLER_46_2632 ();
 sg13g2_decap_8 FILLER_46_2639 ();
 sg13g2_decap_8 FILLER_46_2646 ();
 sg13g2_decap_8 FILLER_46_2653 ();
 sg13g2_decap_8 FILLER_46_2660 ();
 sg13g2_fill_2 FILLER_46_2667 ();
 sg13g2_fill_1 FILLER_46_2669 ();
 sg13g2_fill_1 FILLER_47_69 ();
 sg13g2_fill_2 FILLER_47_73 ();
 sg13g2_fill_1 FILLER_47_75 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_4 FILLER_47_95 ();
 sg13g2_fill_1 FILLER_47_99 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_115 ();
 sg13g2_decap_4 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_129 ();
 sg13g2_decap_8 FILLER_47_136 ();
 sg13g2_decap_8 FILLER_47_143 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_decap_4 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_161 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_fill_1 FILLER_47_190 ();
 sg13g2_decap_8 FILLER_47_239 ();
 sg13g2_decap_8 FILLER_47_277 ();
 sg13g2_decap_8 FILLER_47_284 ();
 sg13g2_decap_8 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_fill_1 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_387 ();
 sg13g2_decap_8 FILLER_47_394 ();
 sg13g2_decap_4 FILLER_47_401 ();
 sg13g2_fill_1 FILLER_47_405 ();
 sg13g2_fill_1 FILLER_47_427 ();
 sg13g2_fill_2 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_517 ();
 sg13g2_decap_8 FILLER_47_523 ();
 sg13g2_decap_8 FILLER_47_536 ();
 sg13g2_decap_8 FILLER_47_543 ();
 sg13g2_decap_8 FILLER_47_550 ();
 sg13g2_decap_8 FILLER_47_557 ();
 sg13g2_decap_4 FILLER_47_564 ();
 sg13g2_fill_2 FILLER_47_568 ();
 sg13g2_fill_2 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_fill_2 FILLER_47_609 ();
 sg13g2_fill_1 FILLER_47_611 ();
 sg13g2_decap_4 FILLER_47_617 ();
 sg13g2_fill_1 FILLER_47_621 ();
 sg13g2_fill_1 FILLER_47_635 ();
 sg13g2_decap_8 FILLER_47_648 ();
 sg13g2_decap_8 FILLER_47_697 ();
 sg13g2_decap_4 FILLER_47_712 ();
 sg13g2_fill_2 FILLER_47_729 ();
 sg13g2_fill_1 FILLER_47_731 ();
 sg13g2_fill_2 FILLER_47_739 ();
 sg13g2_fill_1 FILLER_47_753 ();
 sg13g2_fill_2 FILLER_47_774 ();
 sg13g2_fill_1 FILLER_47_799 ();
 sg13g2_fill_1 FILLER_47_849 ();
 sg13g2_fill_2 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_876 ();
 sg13g2_decap_8 FILLER_47_883 ();
 sg13g2_fill_2 FILLER_47_890 ();
 sg13g2_fill_2 FILLER_47_897 ();
 sg13g2_decap_8 FILLER_47_908 ();
 sg13g2_fill_2 FILLER_47_915 ();
 sg13g2_decap_8 FILLER_47_926 ();
 sg13g2_decap_8 FILLER_47_933 ();
 sg13g2_fill_1 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_972 ();
 sg13g2_decap_4 FILLER_47_979 ();
 sg13g2_decap_4 FILLER_47_988 ();
 sg13g2_fill_1 FILLER_47_1009 ();
 sg13g2_fill_1 FILLER_47_1025 ();
 sg13g2_fill_1 FILLER_47_1030 ();
 sg13g2_decap_8 FILLER_47_1036 ();
 sg13g2_fill_1 FILLER_47_1043 ();
 sg13g2_decap_4 FILLER_47_1049 ();
 sg13g2_decap_8 FILLER_47_1067 ();
 sg13g2_decap_4 FILLER_47_1074 ();
 sg13g2_fill_2 FILLER_47_1087 ();
 sg13g2_fill_1 FILLER_47_1089 ();
 sg13g2_decap_8 FILLER_47_1106 ();
 sg13g2_fill_2 FILLER_47_1119 ();
 sg13g2_fill_1 FILLER_47_1147 ();
 sg13g2_fill_2 FILLER_47_1159 ();
 sg13g2_fill_1 FILLER_47_1161 ();
 sg13g2_fill_1 FILLER_47_1172 ();
 sg13g2_fill_2 FILLER_47_1178 ();
 sg13g2_fill_1 FILLER_47_1180 ();
 sg13g2_decap_8 FILLER_47_1195 ();
 sg13g2_fill_2 FILLER_47_1214 ();
 sg13g2_fill_1 FILLER_47_1216 ();
 sg13g2_fill_1 FILLER_47_1222 ();
 sg13g2_fill_2 FILLER_47_1253 ();
 sg13g2_fill_1 FILLER_47_1255 ();
 sg13g2_decap_8 FILLER_47_1261 ();
 sg13g2_decap_4 FILLER_47_1279 ();
 sg13g2_fill_2 FILLER_47_1287 ();
 sg13g2_fill_2 FILLER_47_1315 ();
 sg13g2_fill_1 FILLER_47_1317 ();
 sg13g2_fill_1 FILLER_47_1344 ();
 sg13g2_decap_8 FILLER_47_1384 ();
 sg13g2_decap_8 FILLER_47_1391 ();
 sg13g2_fill_2 FILLER_47_1403 ();
 sg13g2_fill_1 FILLER_47_1405 ();
 sg13g2_fill_1 FILLER_47_1415 ();
 sg13g2_fill_1 FILLER_47_1470 ();
 sg13g2_fill_1 FILLER_47_1482 ();
 sg13g2_fill_1 FILLER_47_1503 ();
 sg13g2_decap_4 FILLER_47_1508 ();
 sg13g2_fill_1 FILLER_47_1517 ();
 sg13g2_fill_1 FILLER_47_1523 ();
 sg13g2_decap_4 FILLER_47_1529 ();
 sg13g2_fill_2 FILLER_47_1563 ();
 sg13g2_decap_4 FILLER_47_1572 ();
 sg13g2_fill_2 FILLER_47_1576 ();
 sg13g2_fill_1 FILLER_47_1629 ();
 sg13g2_decap_4 FILLER_47_1644 ();
 sg13g2_fill_2 FILLER_47_1679 ();
 sg13g2_fill_1 FILLER_47_1681 ();
 sg13g2_fill_1 FILLER_47_1704 ();
 sg13g2_fill_1 FILLER_47_1715 ();
 sg13g2_fill_2 FILLER_47_1720 ();
 sg13g2_fill_2 FILLER_47_1755 ();
 sg13g2_fill_1 FILLER_47_1757 ();
 sg13g2_decap_4 FILLER_47_1762 ();
 sg13g2_fill_2 FILLER_47_1766 ();
 sg13g2_decap_8 FILLER_47_1773 ();
 sg13g2_fill_1 FILLER_47_1780 ();
 sg13g2_decap_8 FILLER_47_1791 ();
 sg13g2_fill_2 FILLER_47_1798 ();
 sg13g2_fill_1 FILLER_47_1849 ();
 sg13g2_decap_8 FILLER_47_1880 ();
 sg13g2_decap_8 FILLER_47_1887 ();
 sg13g2_decap_8 FILLER_47_1894 ();
 sg13g2_decap_8 FILLER_47_1901 ();
 sg13g2_decap_8 FILLER_47_1908 ();
 sg13g2_decap_4 FILLER_47_1915 ();
 sg13g2_fill_1 FILLER_47_1919 ();
 sg13g2_fill_1 FILLER_47_1929 ();
 sg13g2_fill_1 FILLER_47_1936 ();
 sg13g2_fill_1 FILLER_47_1946 ();
 sg13g2_fill_1 FILLER_47_1956 ();
 sg13g2_decap_8 FILLER_47_1983 ();
 sg13g2_decap_8 FILLER_47_1990 ();
 sg13g2_decap_8 FILLER_47_1997 ();
 sg13g2_decap_8 FILLER_47_2004 ();
 sg13g2_decap_8 FILLER_47_2011 ();
 sg13g2_decap_8 FILLER_47_2018 ();
 sg13g2_decap_4 FILLER_47_2025 ();
 sg13g2_fill_2 FILLER_47_2029 ();
 sg13g2_fill_2 FILLER_47_2034 ();
 sg13g2_decap_8 FILLER_47_2041 ();
 sg13g2_decap_8 FILLER_47_2048 ();
 sg13g2_decap_8 FILLER_47_2055 ();
 sg13g2_decap_8 FILLER_47_2062 ();
 sg13g2_fill_1 FILLER_47_2069 ();
 sg13g2_fill_2 FILLER_47_2096 ();
 sg13g2_fill_1 FILLER_47_2098 ();
 sg13g2_fill_1 FILLER_47_2104 ();
 sg13g2_fill_1 FILLER_47_2164 ();
 sg13g2_fill_2 FILLER_47_2193 ();
 sg13g2_fill_2 FILLER_47_2221 ();
 sg13g2_fill_1 FILLER_47_2223 ();
 sg13g2_fill_2 FILLER_47_2239 ();
 sg13g2_decap_8 FILLER_47_2258 ();
 sg13g2_decap_4 FILLER_47_2265 ();
 sg13g2_fill_2 FILLER_47_2269 ();
 sg13g2_decap_8 FILLER_47_2297 ();
 sg13g2_fill_1 FILLER_47_2304 ();
 sg13g2_decap_4 FILLER_47_2309 ();
 sg13g2_fill_2 FILLER_47_2313 ();
 sg13g2_decap_8 FILLER_47_2320 ();
 sg13g2_decap_8 FILLER_47_2327 ();
 sg13g2_decap_8 FILLER_47_2334 ();
 sg13g2_decap_8 FILLER_47_2341 ();
 sg13g2_fill_2 FILLER_47_2348 ();
 sg13g2_fill_1 FILLER_47_2350 ();
 sg13g2_decap_4 FILLER_47_2386 ();
 sg13g2_fill_2 FILLER_47_2390 ();
 sg13g2_fill_1 FILLER_47_2456 ();
 sg13g2_fill_2 FILLER_47_2461 ();
 sg13g2_fill_2 FILLER_47_2470 ();
 sg13g2_fill_1 FILLER_47_2472 ();
 sg13g2_decap_4 FILLER_47_2499 ();
 sg13g2_decap_4 FILLER_47_2526 ();
 sg13g2_fill_1 FILLER_47_2530 ();
 sg13g2_decap_8 FILLER_47_2561 ();
 sg13g2_decap_8 FILLER_47_2568 ();
 sg13g2_decap_8 FILLER_47_2575 ();
 sg13g2_decap_8 FILLER_47_2582 ();
 sg13g2_decap_8 FILLER_47_2589 ();
 sg13g2_decap_8 FILLER_47_2596 ();
 sg13g2_decap_8 FILLER_47_2603 ();
 sg13g2_decap_8 FILLER_47_2610 ();
 sg13g2_decap_8 FILLER_47_2617 ();
 sg13g2_decap_8 FILLER_47_2624 ();
 sg13g2_decap_8 FILLER_47_2631 ();
 sg13g2_decap_8 FILLER_47_2638 ();
 sg13g2_decap_8 FILLER_47_2645 ();
 sg13g2_decap_8 FILLER_47_2652 ();
 sg13g2_decap_8 FILLER_47_2659 ();
 sg13g2_decap_4 FILLER_47_2666 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_decap_8 FILLER_48_9 ();
 sg13g2_decap_8 FILLER_48_32 ();
 sg13g2_decap_8 FILLER_48_48 ();
 sg13g2_decap_8 FILLER_48_55 ();
 sg13g2_fill_1 FILLER_48_62 ();
 sg13g2_decap_8 FILLER_48_68 ();
 sg13g2_decap_8 FILLER_48_75 ();
 sg13g2_decap_4 FILLER_48_125 ();
 sg13g2_fill_2 FILLER_48_133 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_decap_8 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_146 ();
 sg13g2_fill_2 FILLER_48_173 ();
 sg13g2_fill_2 FILLER_48_231 ();
 sg13g2_fill_2 FILLER_48_255 ();
 sg13g2_decap_8 FILLER_48_271 ();
 sg13g2_fill_2 FILLER_48_278 ();
 sg13g2_fill_1 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_286 ();
 sg13g2_decap_8 FILLER_48_293 ();
 sg13g2_decap_8 FILLER_48_300 ();
 sg13g2_fill_2 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_309 ();
 sg13g2_fill_2 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_fill_2 FILLER_48_396 ();
 sg13g2_fill_2 FILLER_48_451 ();
 sg13g2_fill_1 FILLER_48_453 ();
 sg13g2_decap_4 FILLER_48_465 ();
 sg13g2_decap_8 FILLER_48_477 ();
 sg13g2_decap_8 FILLER_48_484 ();
 sg13g2_decap_4 FILLER_48_491 ();
 sg13g2_fill_1 FILLER_48_495 ();
 sg13g2_fill_2 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_fill_2 FILLER_48_532 ();
 sg13g2_fill_1 FILLER_48_534 ();
 sg13g2_decap_4 FILLER_48_539 ();
 sg13g2_fill_2 FILLER_48_543 ();
 sg13g2_fill_2 FILLER_48_550 ();
 sg13g2_fill_1 FILLER_48_552 ();
 sg13g2_decap_8 FILLER_48_557 ();
 sg13g2_fill_2 FILLER_48_564 ();
 sg13g2_fill_1 FILLER_48_566 ();
 sg13g2_fill_2 FILLER_48_589 ();
 sg13g2_fill_1 FILLER_48_596 ();
 sg13g2_fill_2 FILLER_48_601 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_fill_1 FILLER_48_632 ();
 sg13g2_fill_1 FILLER_48_648 ();
 sg13g2_decap_4 FILLER_48_725 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_fill_1 FILLER_48_754 ();
 sg13g2_fill_1 FILLER_48_768 ();
 sg13g2_fill_2 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_783 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_4 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_833 ();
 sg13g2_fill_2 FILLER_48_852 ();
 sg13g2_fill_1 FILLER_48_854 ();
 sg13g2_fill_1 FILLER_48_864 ();
 sg13g2_decap_4 FILLER_48_869 ();
 sg13g2_fill_1 FILLER_48_873 ();
 sg13g2_fill_2 FILLER_48_878 ();
 sg13g2_fill_1 FILLER_48_884 ();
 sg13g2_fill_2 FILLER_48_889 ();
 sg13g2_fill_1 FILLER_48_891 ();
 sg13g2_decap_8 FILLER_48_906 ();
 sg13g2_decap_4 FILLER_48_913 ();
 sg13g2_decap_8 FILLER_48_923 ();
 sg13g2_decap_8 FILLER_48_947 ();
 sg13g2_decap_8 FILLER_48_954 ();
 sg13g2_decap_8 FILLER_48_961 ();
 sg13g2_fill_2 FILLER_48_968 ();
 sg13g2_fill_1 FILLER_48_988 ();
 sg13g2_fill_1 FILLER_48_994 ();
 sg13g2_fill_1 FILLER_48_1021 ();
 sg13g2_fill_2 FILLER_48_1060 ();
 sg13g2_fill_2 FILLER_48_1095 ();
 sg13g2_fill_1 FILLER_48_1097 ();
 sg13g2_fill_2 FILLER_48_1125 ();
 sg13g2_decap_8 FILLER_48_1137 ();
 sg13g2_decap_8 FILLER_48_1144 ();
 sg13g2_decap_4 FILLER_48_1151 ();
 sg13g2_decap_4 FILLER_48_1189 ();
 sg13g2_fill_2 FILLER_48_1212 ();
 sg13g2_fill_1 FILLER_48_1214 ();
 sg13g2_fill_2 FILLER_48_1239 ();
 sg13g2_fill_1 FILLER_48_1241 ();
 sg13g2_fill_1 FILLER_48_1259 ();
 sg13g2_fill_1 FILLER_48_1265 ();
 sg13g2_fill_1 FILLER_48_1274 ();
 sg13g2_decap_8 FILLER_48_1301 ();
 sg13g2_decap_4 FILLER_48_1308 ();
 sg13g2_fill_1 FILLER_48_1312 ();
 sg13g2_decap_8 FILLER_48_1323 ();
 sg13g2_fill_2 FILLER_48_1345 ();
 sg13g2_fill_1 FILLER_48_1367 ();
 sg13g2_decap_8 FILLER_48_1376 ();
 sg13g2_fill_2 FILLER_48_1383 ();
 sg13g2_fill_1 FILLER_48_1461 ();
 sg13g2_fill_2 FILLER_48_1505 ();
 sg13g2_fill_1 FILLER_48_1507 ();
 sg13g2_fill_2 FILLER_48_1531 ();
 sg13g2_fill_1 FILLER_48_1533 ();
 sg13g2_fill_1 FILLER_48_1579 ();
 sg13g2_fill_1 FILLER_48_1596 ();
 sg13g2_fill_2 FILLER_48_1732 ();
 sg13g2_fill_1 FILLER_48_1734 ();
 sg13g2_decap_4 FILLER_48_1740 ();
 sg13g2_decap_8 FILLER_48_1754 ();
 sg13g2_decap_4 FILLER_48_1761 ();
 sg13g2_fill_1 FILLER_48_1765 ();
 sg13g2_fill_2 FILLER_48_1791 ();
 sg13g2_fill_1 FILLER_48_1793 ();
 sg13g2_decap_8 FILLER_48_1807 ();
 sg13g2_fill_2 FILLER_48_1843 ();
 sg13g2_fill_1 FILLER_48_1853 ();
 sg13g2_fill_2 FILLER_48_1866 ();
 sg13g2_decap_8 FILLER_48_1881 ();
 sg13g2_decap_8 FILLER_48_1888 ();
 sg13g2_fill_2 FILLER_48_1895 ();
 sg13g2_fill_1 FILLER_48_1897 ();
 sg13g2_decap_4 FILLER_48_1903 ();
 sg13g2_fill_1 FILLER_48_1915 ();
 sg13g2_decap_4 FILLER_48_1974 ();
 sg13g2_fill_2 FILLER_48_1978 ();
 sg13g2_decap_8 FILLER_48_2020 ();
 sg13g2_fill_1 FILLER_48_2027 ();
 sg13g2_decap_8 FILLER_48_2037 ();
 sg13g2_decap_4 FILLER_48_2044 ();
 sg13g2_fill_1 FILLER_48_2048 ();
 sg13g2_fill_1 FILLER_48_2104 ();
 sg13g2_fill_2 FILLER_48_2137 ();
 sg13g2_decap_4 FILLER_48_2182 ();
 sg13g2_fill_1 FILLER_48_2186 ();
 sg13g2_decap_8 FILLER_48_2199 ();
 sg13g2_fill_2 FILLER_48_2206 ();
 sg13g2_fill_1 FILLER_48_2208 ();
 sg13g2_decap_8 FILLER_48_2278 ();
 sg13g2_decap_4 FILLER_48_2285 ();
 sg13g2_decap_8 FILLER_48_2295 ();
 sg13g2_decap_8 FILLER_48_2302 ();
 sg13g2_fill_2 FILLER_48_2317 ();
 sg13g2_fill_2 FILLER_48_2323 ();
 sg13g2_fill_1 FILLER_48_2325 ();
 sg13g2_decap_8 FILLER_48_2330 ();
 sg13g2_decap_8 FILLER_48_2350 ();
 sg13g2_decap_8 FILLER_48_2374 ();
 sg13g2_decap_8 FILLER_48_2381 ();
 sg13g2_decap_8 FILLER_48_2388 ();
 sg13g2_decap_8 FILLER_48_2395 ();
 sg13g2_decap_8 FILLER_48_2402 ();
 sg13g2_decap_4 FILLER_48_2409 ();
 sg13g2_fill_1 FILLER_48_2413 ();
 sg13g2_fill_1 FILLER_48_2422 ();
 sg13g2_fill_1 FILLER_48_2458 ();
 sg13g2_decap_8 FILLER_48_2497 ();
 sg13g2_decap_8 FILLER_48_2504 ();
 sg13g2_fill_2 FILLER_48_2511 ();
 sg13g2_decap_8 FILLER_48_2519 ();
 sg13g2_decap_8 FILLER_48_2526 ();
 sg13g2_decap_8 FILLER_48_2533 ();
 sg13g2_decap_8 FILLER_48_2544 ();
 sg13g2_decap_8 FILLER_48_2551 ();
 sg13g2_decap_8 FILLER_48_2558 ();
 sg13g2_decap_8 FILLER_48_2565 ();
 sg13g2_decap_8 FILLER_48_2572 ();
 sg13g2_decap_8 FILLER_48_2579 ();
 sg13g2_decap_8 FILLER_48_2586 ();
 sg13g2_decap_8 FILLER_48_2593 ();
 sg13g2_decap_8 FILLER_48_2600 ();
 sg13g2_decap_8 FILLER_48_2607 ();
 sg13g2_decap_8 FILLER_48_2614 ();
 sg13g2_decap_8 FILLER_48_2621 ();
 sg13g2_decap_8 FILLER_48_2628 ();
 sg13g2_decap_8 FILLER_48_2635 ();
 sg13g2_decap_8 FILLER_48_2642 ();
 sg13g2_decap_8 FILLER_48_2649 ();
 sg13g2_decap_8 FILLER_48_2656 ();
 sg13g2_decap_8 FILLER_48_2663 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_23 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_4 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_decap_4 FILLER_49_148 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_decap_8 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_191 ();
 sg13g2_decap_4 FILLER_49_198 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_fill_1 FILLER_49_229 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_decap_4 FILLER_49_311 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_decap_4 FILLER_49_368 ();
 sg13g2_fill_2 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_379 ();
 sg13g2_decap_4 FILLER_49_385 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_fill_2 FILLER_49_401 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_1 FILLER_49_424 ();
 sg13g2_fill_1 FILLER_49_436 ();
 sg13g2_fill_1 FILLER_49_442 ();
 sg13g2_fill_2 FILLER_49_447 ();
 sg13g2_decap_4 FILLER_49_462 ();
 sg13g2_decap_4 FILLER_49_510 ();
 sg13g2_fill_2 FILLER_49_514 ();
 sg13g2_decap_8 FILLER_49_526 ();
 sg13g2_decap_4 FILLER_49_533 ();
 sg13g2_fill_2 FILLER_49_549 ();
 sg13g2_decap_8 FILLER_49_555 ();
 sg13g2_decap_8 FILLER_49_562 ();
 sg13g2_fill_2 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_590 ();
 sg13g2_fill_2 FILLER_49_600 ();
 sg13g2_fill_1 FILLER_49_602 ();
 sg13g2_fill_1 FILLER_49_613 ();
 sg13g2_fill_1 FILLER_49_625 ();
 sg13g2_fill_2 FILLER_49_637 ();
 sg13g2_fill_2 FILLER_49_649 ();
 sg13g2_fill_1 FILLER_49_656 ();
 sg13g2_decap_4 FILLER_49_675 ();
 sg13g2_fill_1 FILLER_49_679 ();
 sg13g2_fill_2 FILLER_49_685 ();
 sg13g2_fill_2 FILLER_49_694 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_4 FILLER_49_707 ();
 sg13g2_fill_1 FILLER_49_711 ();
 sg13g2_decap_8 FILLER_49_720 ();
 sg13g2_decap_4 FILLER_49_727 ();
 sg13g2_fill_2 FILLER_49_731 ();
 sg13g2_decap_4 FILLER_49_738 ();
 sg13g2_fill_1 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_793 ();
 sg13g2_fill_2 FILLER_49_800 ();
 sg13g2_fill_1 FILLER_49_806 ();
 sg13g2_fill_2 FILLER_49_833 ();
 sg13g2_fill_1 FILLER_49_879 ();
 sg13g2_fill_2 FILLER_49_886 ();
 sg13g2_fill_1 FILLER_49_888 ();
 sg13g2_fill_1 FILLER_49_919 ();
 sg13g2_fill_1 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_934 ();
 sg13g2_fill_2 FILLER_49_947 ();
 sg13g2_decap_8 FILLER_49_961 ();
 sg13g2_fill_2 FILLER_49_976 ();
 sg13g2_fill_1 FILLER_49_978 ();
 sg13g2_fill_1 FILLER_49_1005 ();
 sg13g2_fill_2 FILLER_49_1026 ();
 sg13g2_fill_2 FILLER_49_1040 ();
 sg13g2_fill_2 FILLER_49_1050 ();
 sg13g2_decap_8 FILLER_49_1063 ();
 sg13g2_fill_1 FILLER_49_1070 ();
 sg13g2_decap_8 FILLER_49_1075 ();
 sg13g2_decap_4 FILLER_49_1082 ();
 sg13g2_fill_1 FILLER_49_1086 ();
 sg13g2_fill_1 FILLER_49_1123 ();
 sg13g2_decap_4 FILLER_49_1145 ();
 sg13g2_decap_8 FILLER_49_1154 ();
 sg13g2_decap_8 FILLER_49_1161 ();
 sg13g2_decap_8 FILLER_49_1188 ();
 sg13g2_fill_2 FILLER_49_1195 ();
 sg13g2_fill_1 FILLER_49_1207 ();
 sg13g2_fill_1 FILLER_49_1214 ();
 sg13g2_fill_1 FILLER_49_1235 ();
 sg13g2_fill_2 FILLER_49_1244 ();
 sg13g2_decap_8 FILLER_49_1261 ();
 sg13g2_decap_8 FILLER_49_1268 ();
 sg13g2_fill_2 FILLER_49_1275 ();
 sg13g2_fill_1 FILLER_49_1277 ();
 sg13g2_decap_4 FILLER_49_1291 ();
 sg13g2_fill_1 FILLER_49_1358 ();
 sg13g2_fill_2 FILLER_49_1364 ();
 sg13g2_fill_1 FILLER_49_1392 ();
 sg13g2_decap_8 FILLER_49_1485 ();
 sg13g2_decap_8 FILLER_49_1492 ();
 sg13g2_decap_8 FILLER_49_1499 ();
 sg13g2_decap_8 FILLER_49_1506 ();
 sg13g2_decap_8 FILLER_49_1513 ();
 sg13g2_decap_8 FILLER_49_1520 ();
 sg13g2_decap_8 FILLER_49_1527 ();
 sg13g2_decap_8 FILLER_49_1544 ();
 sg13g2_decap_4 FILLER_49_1551 ();
 sg13g2_fill_1 FILLER_49_1577 ();
 sg13g2_fill_2 FILLER_49_1583 ();
 sg13g2_fill_1 FILLER_49_1605 ();
 sg13g2_decap_8 FILLER_49_1648 ();
 sg13g2_decap_8 FILLER_49_1655 ();
 sg13g2_fill_2 FILLER_49_1685 ();
 sg13g2_fill_1 FILLER_49_1693 ();
 sg13g2_fill_2 FILLER_49_1700 ();
 sg13g2_decap_4 FILLER_49_1728 ();
 sg13g2_decap_4 FILLER_49_1740 ();
 sg13g2_fill_2 FILLER_49_1752 ();
 sg13g2_fill_1 FILLER_49_1764 ();
 sg13g2_fill_1 FILLER_49_1769 ();
 sg13g2_fill_1 FILLER_49_1798 ();
 sg13g2_fill_2 FILLER_49_1817 ();
 sg13g2_fill_1 FILLER_49_1819 ();
 sg13g2_fill_2 FILLER_49_1855 ();
 sg13g2_decap_8 FILLER_49_1872 ();
 sg13g2_fill_2 FILLER_49_1884 ();
 sg13g2_fill_2 FILLER_49_1957 ();
 sg13g2_decap_8 FILLER_49_1990 ();
 sg13g2_decap_8 FILLER_49_1997 ();
 sg13g2_decap_4 FILLER_49_2004 ();
 sg13g2_fill_1 FILLER_49_2008 ();
 sg13g2_fill_2 FILLER_49_2039 ();
 sg13g2_fill_1 FILLER_49_2041 ();
 sg13g2_decap_8 FILLER_49_2097 ();
 sg13g2_fill_1 FILLER_49_2104 ();
 sg13g2_decap_8 FILLER_49_2114 ();
 sg13g2_decap_8 FILLER_49_2121 ();
 sg13g2_decap_8 FILLER_49_2167 ();
 sg13g2_decap_4 FILLER_49_2174 ();
 sg13g2_fill_2 FILLER_49_2221 ();
 sg13g2_fill_2 FILLER_49_2228 ();
 sg13g2_decap_4 FILLER_49_2244 ();
 sg13g2_fill_2 FILLER_49_2285 ();
 sg13g2_fill_1 FILLER_49_2287 ();
 sg13g2_decap_8 FILLER_49_2344 ();
 sg13g2_decap_8 FILLER_49_2351 ();
 sg13g2_decap_8 FILLER_49_2358 ();
 sg13g2_decap_8 FILLER_49_2365 ();
 sg13g2_decap_8 FILLER_49_2372 ();
 sg13g2_decap_8 FILLER_49_2379 ();
 sg13g2_decap_8 FILLER_49_2386 ();
 sg13g2_decap_8 FILLER_49_2393 ();
 sg13g2_fill_2 FILLER_49_2400 ();
 sg13g2_decap_4 FILLER_49_2428 ();
 sg13g2_fill_1 FILLER_49_2432 ();
 sg13g2_decap_8 FILLER_49_2466 ();
 sg13g2_decap_4 FILLER_49_2473 ();
 sg13g2_fill_1 FILLER_49_2477 ();
 sg13g2_decap_8 FILLER_49_2482 ();
 sg13g2_decap_8 FILLER_49_2489 ();
 sg13g2_decap_8 FILLER_49_2503 ();
 sg13g2_fill_1 FILLER_49_2510 ();
 sg13g2_decap_8 FILLER_49_2519 ();
 sg13g2_decap_8 FILLER_49_2526 ();
 sg13g2_decap_8 FILLER_49_2533 ();
 sg13g2_decap_8 FILLER_49_2566 ();
 sg13g2_decap_8 FILLER_49_2573 ();
 sg13g2_decap_8 FILLER_49_2580 ();
 sg13g2_decap_8 FILLER_49_2587 ();
 sg13g2_decap_8 FILLER_49_2594 ();
 sg13g2_decap_8 FILLER_49_2601 ();
 sg13g2_decap_8 FILLER_49_2608 ();
 sg13g2_decap_8 FILLER_49_2615 ();
 sg13g2_decap_8 FILLER_49_2622 ();
 sg13g2_decap_8 FILLER_49_2629 ();
 sg13g2_decap_8 FILLER_49_2636 ();
 sg13g2_decap_8 FILLER_49_2643 ();
 sg13g2_decap_8 FILLER_49_2650 ();
 sg13g2_decap_8 FILLER_49_2657 ();
 sg13g2_decap_4 FILLER_49_2664 ();
 sg13g2_fill_2 FILLER_49_2668 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_37 ();
 sg13g2_fill_1 FILLER_50_65 ();
 sg13g2_fill_2 FILLER_50_70 ();
 sg13g2_fill_1 FILLER_50_72 ();
 sg13g2_fill_1 FILLER_50_78 ();
 sg13g2_decap_8 FILLER_50_83 ();
 sg13g2_decap_4 FILLER_50_90 ();
 sg13g2_fill_2 FILLER_50_94 ();
 sg13g2_fill_2 FILLER_50_118 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_fill_1 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_fill_2 FILLER_50_149 ();
 sg13g2_decap_8 FILLER_50_186 ();
 sg13g2_fill_2 FILLER_50_193 ();
 sg13g2_fill_1 FILLER_50_195 ();
 sg13g2_fill_2 FILLER_50_237 ();
 sg13g2_fill_2 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_246 ();
 sg13g2_fill_2 FILLER_50_252 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_fill_2 FILLER_50_264 ();
 sg13g2_fill_1 FILLER_50_266 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_decap_8 FILLER_50_317 ();
 sg13g2_decap_4 FILLER_50_324 ();
 sg13g2_fill_2 FILLER_50_328 ();
 sg13g2_fill_2 FILLER_50_336 ();
 sg13g2_decap_4 FILLER_50_344 ();
 sg13g2_fill_1 FILLER_50_348 ();
 sg13g2_decap_4 FILLER_50_391 ();
 sg13g2_fill_1 FILLER_50_395 ();
 sg13g2_fill_2 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_413 ();
 sg13g2_fill_2 FILLER_50_422 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_decap_8 FILLER_50_442 ();
 sg13g2_fill_2 FILLER_50_449 ();
 sg13g2_fill_1 FILLER_50_451 ();
 sg13g2_decap_8 FILLER_50_480 ();
 sg13g2_decap_4 FILLER_50_487 ();
 sg13g2_fill_1 FILLER_50_491 ();
 sg13g2_decap_8 FILLER_50_495 ();
 sg13g2_fill_2 FILLER_50_502 ();
 sg13g2_fill_2 FILLER_50_528 ();
 sg13g2_decap_8 FILLER_50_540 ();
 sg13g2_fill_2 FILLER_50_547 ();
 sg13g2_decap_8 FILLER_50_572 ();
 sg13g2_fill_1 FILLER_50_579 ();
 sg13g2_fill_2 FILLER_50_591 ();
 sg13g2_fill_1 FILLER_50_593 ();
 sg13g2_decap_4 FILLER_50_598 ();
 sg13g2_fill_1 FILLER_50_602 ();
 sg13g2_fill_1 FILLER_50_612 ();
 sg13g2_fill_1 FILLER_50_628 ();
 sg13g2_fill_1 FILLER_50_639 ();
 sg13g2_fill_1 FILLER_50_655 ();
 sg13g2_decap_4 FILLER_50_660 ();
 sg13g2_fill_1 FILLER_50_664 ();
 sg13g2_fill_1 FILLER_50_681 ();
 sg13g2_decap_4 FILLER_50_747 ();
 sg13g2_fill_2 FILLER_50_755 ();
 sg13g2_fill_1 FILLER_50_757 ();
 sg13g2_decap_8 FILLER_50_764 ();
 sg13g2_decap_4 FILLER_50_777 ();
 sg13g2_fill_2 FILLER_50_781 ();
 sg13g2_decap_8 FILLER_50_796 ();
 sg13g2_fill_1 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_827 ();
 sg13g2_fill_2 FILLER_50_834 ();
 sg13g2_fill_1 FILLER_50_836 ();
 sg13g2_fill_1 FILLER_50_867 ();
 sg13g2_fill_1 FILLER_50_904 ();
 sg13g2_decap_4 FILLER_50_936 ();
 sg13g2_fill_1 FILLER_50_940 ();
 sg13g2_decap_8 FILLER_50_946 ();
 sg13g2_decap_4 FILLER_50_953 ();
 sg13g2_decap_4 FILLER_50_962 ();
 sg13g2_fill_1 FILLER_50_982 ();
 sg13g2_decap_8 FILLER_50_989 ();
 sg13g2_fill_1 FILLER_50_996 ();
 sg13g2_fill_1 FILLER_50_1009 ();
 sg13g2_fill_2 FILLER_50_1016 ();
 sg13g2_fill_1 FILLER_50_1023 ();
 sg13g2_fill_2 FILLER_50_1031 ();
 sg13g2_decap_8 FILLER_50_1068 ();
 sg13g2_decap_8 FILLER_50_1075 ();
 sg13g2_decap_4 FILLER_50_1082 ();
 sg13g2_fill_2 FILLER_50_1086 ();
 sg13g2_decap_8 FILLER_50_1114 ();
 sg13g2_decap_8 FILLER_50_1136 ();
 sg13g2_decap_4 FILLER_50_1143 ();
 sg13g2_decap_8 FILLER_50_1178 ();
 sg13g2_fill_2 FILLER_50_1185 ();
 sg13g2_fill_2 FILLER_50_1191 ();
 sg13g2_fill_1 FILLER_50_1193 ();
 sg13g2_decap_8 FILLER_50_1251 ();
 sg13g2_decap_8 FILLER_50_1258 ();
 sg13g2_decap_8 FILLER_50_1265 ();
 sg13g2_fill_2 FILLER_50_1272 ();
 sg13g2_decap_8 FILLER_50_1280 ();
 sg13g2_fill_1 FILLER_50_1287 ();
 sg13g2_decap_8 FILLER_50_1293 ();
 sg13g2_fill_2 FILLER_50_1300 ();
 sg13g2_fill_2 FILLER_50_1328 ();
 sg13g2_fill_1 FILLER_50_1336 ();
 sg13g2_decap_4 FILLER_50_1344 ();
 sg13g2_fill_1 FILLER_50_1353 ();
 sg13g2_decap_8 FILLER_50_1380 ();
 sg13g2_decap_4 FILLER_50_1387 ();
 sg13g2_fill_2 FILLER_50_1391 ();
 sg13g2_fill_1 FILLER_50_1397 ();
 sg13g2_fill_2 FILLER_50_1437 ();
 sg13g2_fill_2 FILLER_50_1464 ();
 sg13g2_fill_1 FILLER_50_1466 ();
 sg13g2_fill_1 FILLER_50_1472 ();
 sg13g2_decap_8 FILLER_50_1513 ();
 sg13g2_decap_8 FILLER_50_1520 ();
 sg13g2_decap_8 FILLER_50_1553 ();
 sg13g2_decap_8 FILLER_50_1560 ();
 sg13g2_fill_2 FILLER_50_1567 ();
 sg13g2_fill_1 FILLER_50_1569 ();
 sg13g2_fill_2 FILLER_50_1574 ();
 sg13g2_fill_2 FILLER_50_1581 ();
 sg13g2_decap_8 FILLER_50_1618 ();
 sg13g2_fill_1 FILLER_50_1625 ();
 sg13g2_decap_8 FILLER_50_1644 ();
 sg13g2_decap_8 FILLER_50_1651 ();
 sg13g2_fill_2 FILLER_50_1680 ();
 sg13g2_fill_2 FILLER_50_1714 ();
 sg13g2_decap_8 FILLER_50_1720 ();
 sg13g2_decap_4 FILLER_50_1727 ();
 sg13g2_fill_2 FILLER_50_1731 ();
 sg13g2_decap_8 FILLER_50_1741 ();
 sg13g2_decap_4 FILLER_50_1748 ();
 sg13g2_fill_1 FILLER_50_1752 ();
 sg13g2_decap_8 FILLER_50_1758 ();
 sg13g2_decap_4 FILLER_50_1765 ();
 sg13g2_fill_1 FILLER_50_1769 ();
 sg13g2_decap_4 FILLER_50_1780 ();
 sg13g2_fill_1 FILLER_50_1784 ();
 sg13g2_decap_8 FILLER_50_1799 ();
 sg13g2_fill_1 FILLER_50_1806 ();
 sg13g2_fill_1 FILLER_50_1812 ();
 sg13g2_decap_8 FILLER_50_1818 ();
 sg13g2_decap_4 FILLER_50_1825 ();
 sg13g2_fill_2 FILLER_50_1829 ();
 sg13g2_fill_1 FILLER_50_1856 ();
 sg13g2_decap_8 FILLER_50_1895 ();
 sg13g2_decap_8 FILLER_50_1902 ();
 sg13g2_decap_8 FILLER_50_1909 ();
 sg13g2_fill_2 FILLER_50_1926 ();
 sg13g2_decap_4 FILLER_50_1932 ();
 sg13g2_decap_8 FILLER_50_1942 ();
 sg13g2_fill_1 FILLER_50_1949 ();
 sg13g2_fill_1 FILLER_50_1955 ();
 sg13g2_decap_4 FILLER_50_1988 ();
 sg13g2_fill_2 FILLER_50_1992 ();
 sg13g2_decap_8 FILLER_50_2008 ();
 sg13g2_decap_8 FILLER_50_2025 ();
 sg13g2_fill_2 FILLER_50_2032 ();
 sg13g2_fill_1 FILLER_50_2034 ();
 sg13g2_fill_2 FILLER_50_2047 ();
 sg13g2_fill_2 FILLER_50_2059 ();
 sg13g2_decap_8 FILLER_50_2094 ();
 sg13g2_decap_4 FILLER_50_2101 ();
 sg13g2_decap_8 FILLER_50_2109 ();
 sg13g2_decap_8 FILLER_50_2116 ();
 sg13g2_fill_1 FILLER_50_2123 ();
 sg13g2_decap_8 FILLER_50_2133 ();
 sg13g2_decap_8 FILLER_50_2145 ();
 sg13g2_fill_2 FILLER_50_2197 ();
 sg13g2_decap_8 FILLER_50_2229 ();
 sg13g2_decap_8 FILLER_50_2236 ();
 sg13g2_decap_4 FILLER_50_2243 ();
 sg13g2_fill_1 FILLER_50_2247 ();
 sg13g2_fill_2 FILLER_50_2257 ();
 sg13g2_decap_8 FILLER_50_2342 ();
 sg13g2_decap_8 FILLER_50_2349 ();
 sg13g2_fill_1 FILLER_50_2356 ();
 sg13g2_decap_8 FILLER_50_2387 ();
 sg13g2_decap_8 FILLER_50_2402 ();
 sg13g2_fill_2 FILLER_50_2409 ();
 sg13g2_fill_2 FILLER_50_2415 ();
 sg13g2_fill_1 FILLER_50_2417 ();
 sg13g2_decap_4 FILLER_50_2424 ();
 sg13g2_decap_8 FILLER_50_2470 ();
 sg13g2_decap_8 FILLER_50_2477 ();
 sg13g2_fill_1 FILLER_50_2484 ();
 sg13g2_fill_2 FILLER_50_2545 ();
 sg13g2_decap_8 FILLER_50_2551 ();
 sg13g2_decap_8 FILLER_50_2558 ();
 sg13g2_fill_1 FILLER_50_2565 ();
 sg13g2_decap_8 FILLER_50_2570 ();
 sg13g2_decap_8 FILLER_50_2577 ();
 sg13g2_decap_8 FILLER_50_2584 ();
 sg13g2_decap_8 FILLER_50_2591 ();
 sg13g2_decap_8 FILLER_50_2598 ();
 sg13g2_decap_8 FILLER_50_2605 ();
 sg13g2_decap_8 FILLER_50_2612 ();
 sg13g2_decap_8 FILLER_50_2619 ();
 sg13g2_decap_8 FILLER_50_2626 ();
 sg13g2_decap_8 FILLER_50_2633 ();
 sg13g2_decap_8 FILLER_50_2640 ();
 sg13g2_decap_8 FILLER_50_2647 ();
 sg13g2_decap_8 FILLER_50_2654 ();
 sg13g2_decap_8 FILLER_50_2661 ();
 sg13g2_fill_2 FILLER_50_2668 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_83 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_decap_4 FILLER_51_149 ();
 sg13g2_fill_1 FILLER_51_153 ();
 sg13g2_decap_8 FILLER_51_163 ();
 sg13g2_decap_8 FILLER_51_170 ();
 sg13g2_decap_8 FILLER_51_177 ();
 sg13g2_decap_8 FILLER_51_184 ();
 sg13g2_decap_8 FILLER_51_191 ();
 sg13g2_fill_2 FILLER_51_198 ();
 sg13g2_fill_2 FILLER_51_213 ();
 sg13g2_fill_1 FILLER_51_222 ();
 sg13g2_decap_4 FILLER_51_228 ();
 sg13g2_fill_1 FILLER_51_232 ();
 sg13g2_decap_8 FILLER_51_241 ();
 sg13g2_decap_4 FILLER_51_253 ();
 sg13g2_fill_1 FILLER_51_257 ();
 sg13g2_decap_8 FILLER_51_264 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_1 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_288 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_fill_1 FILLER_51_300 ();
 sg13g2_fill_2 FILLER_51_336 ();
 sg13g2_decap_4 FILLER_51_343 ();
 sg13g2_fill_2 FILLER_51_362 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_fill_2 FILLER_51_399 ();
 sg13g2_fill_1 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_417 ();
 sg13g2_fill_1 FILLER_51_422 ();
 sg13g2_fill_2 FILLER_51_427 ();
 sg13g2_fill_1 FILLER_51_434 ();
 sg13g2_decap_8 FILLER_51_440 ();
 sg13g2_decap_8 FILLER_51_447 ();
 sg13g2_decap_8 FILLER_51_454 ();
 sg13g2_fill_2 FILLER_51_461 ();
 sg13g2_fill_1 FILLER_51_468 ();
 sg13g2_decap_8 FILLER_51_474 ();
 sg13g2_decap_8 FILLER_51_490 ();
 sg13g2_decap_8 FILLER_51_497 ();
 sg13g2_fill_2 FILLER_51_504 ();
 sg13g2_fill_1 FILLER_51_506 ();
 sg13g2_decap_8 FILLER_51_515 ();
 sg13g2_decap_4 FILLER_51_522 ();
 sg13g2_fill_2 FILLER_51_530 ();
 sg13g2_fill_1 FILLER_51_532 ();
 sg13g2_fill_2 FILLER_51_548 ();
 sg13g2_decap_8 FILLER_51_559 ();
 sg13g2_decap_8 FILLER_51_566 ();
 sg13g2_decap_4 FILLER_51_573 ();
 sg13g2_fill_1 FILLER_51_577 ();
 sg13g2_decap_8 FILLER_51_591 ();
 sg13g2_decap_8 FILLER_51_598 ();
 sg13g2_fill_1 FILLER_51_615 ();
 sg13g2_fill_2 FILLER_51_629 ();
 sg13g2_fill_1 FILLER_51_638 ();
 sg13g2_decap_8 FILLER_51_646 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_fill_1 FILLER_51_687 ();
 sg13g2_fill_1 FILLER_51_700 ();
 sg13g2_decap_4 FILLER_51_714 ();
 sg13g2_decap_4 FILLER_51_743 ();
 sg13g2_decap_4 FILLER_51_782 ();
 sg13g2_fill_1 FILLER_51_786 ();
 sg13g2_decap_4 FILLER_51_792 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_4 FILLER_51_850 ();
 sg13g2_fill_1 FILLER_51_854 ();
 sg13g2_fill_1 FILLER_51_859 ();
 sg13g2_fill_2 FILLER_51_864 ();
 sg13g2_decap_8 FILLER_51_877 ();
 sg13g2_decap_8 FILLER_51_884 ();
 sg13g2_fill_2 FILLER_51_891 ();
 sg13g2_fill_1 FILLER_51_893 ();
 sg13g2_decap_4 FILLER_51_904 ();
 sg13g2_decap_8 FILLER_51_915 ();
 sg13g2_fill_1 FILLER_51_922 ();
 sg13g2_decap_8 FILLER_51_983 ();
 sg13g2_decap_4 FILLER_51_990 ();
 sg13g2_fill_1 FILLER_51_994 ();
 sg13g2_decap_8 FILLER_51_1008 ();
 sg13g2_fill_1 FILLER_51_1015 ();
 sg13g2_fill_1 FILLER_51_1038 ();
 sg13g2_decap_8 FILLER_51_1056 ();
 sg13g2_decap_4 FILLER_51_1063 ();
 sg13g2_fill_1 FILLER_51_1067 ();
 sg13g2_decap_4 FILLER_51_1103 ();
 sg13g2_fill_1 FILLER_51_1107 ();
 sg13g2_fill_2 FILLER_51_1112 ();
 sg13g2_fill_2 FILLER_51_1120 ();
 sg13g2_decap_8 FILLER_51_1174 ();
 sg13g2_decap_4 FILLER_51_1181 ();
 sg13g2_fill_2 FILLER_51_1185 ();
 sg13g2_decap_8 FILLER_51_1192 ();
 sg13g2_fill_2 FILLER_51_1199 ();
 sg13g2_fill_2 FILLER_51_1206 ();
 sg13g2_fill_1 FILLER_51_1208 ();
 sg13g2_decap_4 FILLER_51_1219 ();
 sg13g2_decap_8 FILLER_51_1231 ();
 sg13g2_fill_2 FILLER_51_1243 ();
 sg13g2_fill_1 FILLER_51_1245 ();
 sg13g2_fill_2 FILLER_51_1259 ();
 sg13g2_fill_1 FILLER_51_1261 ();
 sg13g2_decap_8 FILLER_51_1268 ();
 sg13g2_decap_8 FILLER_51_1275 ();
 sg13g2_decap_8 FILLER_51_1290 ();
 sg13g2_decap_8 FILLER_51_1297 ();
 sg13g2_fill_2 FILLER_51_1304 ();
 sg13g2_fill_1 FILLER_51_1306 ();
 sg13g2_fill_2 FILLER_51_1317 ();
 sg13g2_decap_8 FILLER_51_1340 ();
 sg13g2_decap_8 FILLER_51_1347 ();
 sg13g2_decap_8 FILLER_51_1354 ();
 sg13g2_fill_2 FILLER_51_1361 ();
 sg13g2_fill_1 FILLER_51_1363 ();
 sg13g2_decap_8 FILLER_51_1369 ();
 sg13g2_decap_8 FILLER_51_1382 ();
 sg13g2_decap_8 FILLER_51_1389 ();
 sg13g2_fill_2 FILLER_51_1396 ();
 sg13g2_decap_8 FILLER_51_1402 ();
 sg13g2_decap_4 FILLER_51_1409 ();
 sg13g2_fill_2 FILLER_51_1413 ();
 sg13g2_fill_1 FILLER_51_1447 ();
 sg13g2_decap_8 FILLER_51_1486 ();
 sg13g2_decap_8 FILLER_51_1493 ();
 sg13g2_decap_8 FILLER_51_1500 ();
 sg13g2_fill_1 FILLER_51_1543 ();
 sg13g2_decap_8 FILLER_51_1557 ();
 sg13g2_fill_2 FILLER_51_1564 ();
 sg13g2_decap_8 FILLER_51_1607 ();
 sg13g2_decap_8 FILLER_51_1614 ();
 sg13g2_decap_8 FILLER_51_1621 ();
 sg13g2_decap_8 FILLER_51_1628 ();
 sg13g2_fill_2 FILLER_51_1635 ();
 sg13g2_decap_8 FILLER_51_1652 ();
 sg13g2_fill_1 FILLER_51_1664 ();
 sg13g2_fill_2 FILLER_51_1694 ();
 sg13g2_fill_1 FILLER_51_1696 ();
 sg13g2_fill_2 FILLER_51_1703 ();
 sg13g2_fill_1 FILLER_51_1705 ();
 sg13g2_decap_4 FILLER_51_1725 ();
 sg13g2_fill_1 FILLER_51_1729 ();
 sg13g2_decap_8 FILLER_51_1735 ();
 sg13g2_decap_8 FILLER_51_1742 ();
 sg13g2_decap_8 FILLER_51_1749 ();
 sg13g2_decap_8 FILLER_51_1756 ();
 sg13g2_decap_8 FILLER_51_1763 ();
 sg13g2_decap_8 FILLER_51_1770 ();
 sg13g2_decap_8 FILLER_51_1777 ();
 sg13g2_fill_2 FILLER_51_1784 ();
 sg13g2_fill_1 FILLER_51_1786 ();
 sg13g2_decap_8 FILLER_51_1791 ();
 sg13g2_decap_8 FILLER_51_1798 ();
 sg13g2_decap_8 FILLER_51_1818 ();
 sg13g2_decap_8 FILLER_51_1825 ();
 sg13g2_decap_8 FILLER_51_1832 ();
 sg13g2_fill_1 FILLER_51_1839 ();
 sg13g2_decap_8 FILLER_51_1845 ();
 sg13g2_fill_2 FILLER_51_1852 ();
 sg13g2_decap_8 FILLER_51_1870 ();
 sg13g2_decap_4 FILLER_51_1877 ();
 sg13g2_fill_2 FILLER_51_1881 ();
 sg13g2_decap_8 FILLER_51_1889 ();
 sg13g2_decap_8 FILLER_51_1896 ();
 sg13g2_decap_8 FILLER_51_1903 ();
 sg13g2_decap_8 FILLER_51_1910 ();
 sg13g2_fill_2 FILLER_51_1917 ();
 sg13g2_decap_8 FILLER_51_1924 ();
 sg13g2_fill_1 FILLER_51_1931 ();
 sg13g2_fill_1 FILLER_51_1938 ();
 sg13g2_fill_1 FILLER_51_1944 ();
 sg13g2_decap_8 FILLER_51_1949 ();
 sg13g2_decap_4 FILLER_51_1956 ();
 sg13g2_fill_1 FILLER_51_1960 ();
 sg13g2_decap_4 FILLER_51_1966 ();
 sg13g2_fill_1 FILLER_51_1970 ();
 sg13g2_fill_2 FILLER_51_1988 ();
 sg13g2_decap_8 FILLER_51_2020 ();
 sg13g2_decap_8 FILLER_51_2027 ();
 sg13g2_decap_4 FILLER_51_2034 ();
 sg13g2_fill_2 FILLER_51_2042 ();
 sg13g2_decap_8 FILLER_51_2053 ();
 sg13g2_fill_2 FILLER_51_2068 ();
 sg13g2_decap_4 FILLER_51_2075 ();
 sg13g2_fill_1 FILLER_51_2079 ();
 sg13g2_decap_8 FILLER_51_2111 ();
 sg13g2_decap_8 FILLER_51_2118 ();
 sg13g2_fill_1 FILLER_51_2125 ();
 sg13g2_decap_8 FILLER_51_2187 ();
 sg13g2_decap_4 FILLER_51_2194 ();
 sg13g2_fill_1 FILLER_51_2198 ();
 sg13g2_decap_4 FILLER_51_2204 ();
 sg13g2_fill_1 FILLER_51_2208 ();
 sg13g2_decap_8 FILLER_51_2235 ();
 sg13g2_decap_8 FILLER_51_2242 ();
 sg13g2_decap_8 FILLER_51_2249 ();
 sg13g2_decap_8 FILLER_51_2256 ();
 sg13g2_decap_8 FILLER_51_2263 ();
 sg13g2_decap_8 FILLER_51_2270 ();
 sg13g2_fill_1 FILLER_51_2277 ();
 sg13g2_fill_1 FILLER_51_2310 ();
 sg13g2_fill_1 FILLER_51_2328 ();
 sg13g2_fill_2 FILLER_51_2355 ();
 sg13g2_decap_8 FILLER_51_2362 ();
 sg13g2_decap_8 FILLER_51_2369 ();
 sg13g2_decap_4 FILLER_51_2376 ();
 sg13g2_fill_1 FILLER_51_2463 ();
 sg13g2_fill_2 FILLER_51_2532 ();
 sg13g2_fill_2 FILLER_51_2538 ();
 sg13g2_fill_1 FILLER_51_2540 ();
 sg13g2_decap_4 FILLER_51_2551 ();
 sg13g2_decap_8 FILLER_51_2585 ();
 sg13g2_decap_8 FILLER_51_2592 ();
 sg13g2_decap_8 FILLER_51_2599 ();
 sg13g2_decap_8 FILLER_51_2606 ();
 sg13g2_decap_8 FILLER_51_2613 ();
 sg13g2_decap_8 FILLER_51_2620 ();
 sg13g2_decap_8 FILLER_51_2627 ();
 sg13g2_decap_8 FILLER_51_2634 ();
 sg13g2_decap_8 FILLER_51_2641 ();
 sg13g2_decap_8 FILLER_51_2648 ();
 sg13g2_decap_8 FILLER_51_2655 ();
 sg13g2_decap_8 FILLER_51_2662 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_76 ();
 sg13g2_decap_8 FILLER_52_82 ();
 sg13g2_decap_4 FILLER_52_89 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_decap_4 FILLER_52_98 ();
 sg13g2_decap_4 FILLER_52_116 ();
 sg13g2_fill_1 FILLER_52_120 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_157 ();
 sg13g2_decap_8 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_171 ();
 sg13g2_fill_2 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_235 ();
 sg13g2_decap_4 FILLER_52_241 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_274 ();
 sg13g2_fill_2 FILLER_52_336 ();
 sg13g2_fill_1 FILLER_52_354 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_decap_4 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_fill_2 FILLER_52_402 ();
 sg13g2_fill_1 FILLER_52_404 ();
 sg13g2_fill_2 FILLER_52_426 ();
 sg13g2_fill_1 FILLER_52_428 ();
 sg13g2_decap_4 FILLER_52_443 ();
 sg13g2_fill_1 FILLER_52_447 ();
 sg13g2_decap_8 FILLER_52_459 ();
 sg13g2_decap_8 FILLER_52_466 ();
 sg13g2_decap_8 FILLER_52_478 ();
 sg13g2_decap_8 FILLER_52_485 ();
 sg13g2_decap_4 FILLER_52_492 ();
 sg13g2_fill_2 FILLER_52_496 ();
 sg13g2_fill_2 FILLER_52_508 ();
 sg13g2_decap_4 FILLER_52_515 ();
 sg13g2_fill_1 FILLER_52_519 ();
 sg13g2_fill_2 FILLER_52_526 ();
 sg13g2_decap_8 FILLER_52_548 ();
 sg13g2_fill_1 FILLER_52_555 ();
 sg13g2_fill_2 FILLER_52_561 ();
 sg13g2_fill_1 FILLER_52_563 ();
 sg13g2_decap_4 FILLER_52_586 ();
 sg13g2_decap_8 FILLER_52_595 ();
 sg13g2_fill_1 FILLER_52_602 ();
 sg13g2_fill_2 FILLER_52_608 ();
 sg13g2_decap_4 FILLER_52_614 ();
 sg13g2_fill_1 FILLER_52_623 ();
 sg13g2_fill_2 FILLER_52_638 ();
 sg13g2_decap_4 FILLER_52_648 ();
 sg13g2_decap_8 FILLER_52_657 ();
 sg13g2_fill_2 FILLER_52_690 ();
 sg13g2_fill_2 FILLER_52_713 ();
 sg13g2_fill_1 FILLER_52_715 ();
 sg13g2_decap_8 FILLER_52_721 ();
 sg13g2_fill_1 FILLER_52_728 ();
 sg13g2_fill_1 FILLER_52_733 ();
 sg13g2_decap_8 FILLER_52_746 ();
 sg13g2_decap_8 FILLER_52_753 ();
 sg13g2_decap_8 FILLER_52_760 ();
 sg13g2_decap_8 FILLER_52_767 ();
 sg13g2_fill_2 FILLER_52_779 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_decap_4 FILLER_52_800 ();
 sg13g2_fill_1 FILLER_52_804 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_fill_2 FILLER_52_836 ();
 sg13g2_fill_1 FILLER_52_838 ();
 sg13g2_decap_8 FILLER_52_843 ();
 sg13g2_decap_4 FILLER_52_850 ();
 sg13g2_fill_2 FILLER_52_854 ();
 sg13g2_decap_8 FILLER_52_866 ();
 sg13g2_decap_8 FILLER_52_873 ();
 sg13g2_decap_8 FILLER_52_880 ();
 sg13g2_decap_8 FILLER_52_887 ();
 sg13g2_fill_2 FILLER_52_894 ();
 sg13g2_fill_1 FILLER_52_904 ();
 sg13g2_decap_4 FILLER_52_910 ();
 sg13g2_fill_2 FILLER_52_914 ();
 sg13g2_decap_8 FILLER_52_925 ();
 sg13g2_decap_4 FILLER_52_936 ();
 sg13g2_fill_2 FILLER_52_940 ();
 sg13g2_decap_8 FILLER_52_947 ();
 sg13g2_decap_4 FILLER_52_954 ();
 sg13g2_fill_2 FILLER_52_958 ();
 sg13g2_decap_8 FILLER_52_964 ();
 sg13g2_fill_2 FILLER_52_971 ();
 sg13g2_fill_1 FILLER_52_973 ();
 sg13g2_decap_8 FILLER_52_1004 ();
 sg13g2_decap_4 FILLER_52_1011 ();
 sg13g2_decap_8 FILLER_52_1019 ();
 sg13g2_fill_2 FILLER_52_1026 ();
 sg13g2_decap_4 FILLER_52_1031 ();
 sg13g2_fill_2 FILLER_52_1107 ();
 sg13g2_fill_1 FILLER_52_1109 ();
 sg13g2_fill_1 FILLER_52_1118 ();
 sg13g2_fill_2 FILLER_52_1151 ();
 sg13g2_fill_1 FILLER_52_1153 ();
 sg13g2_decap_8 FILLER_52_1164 ();
 sg13g2_decap_8 FILLER_52_1171 ();
 sg13g2_fill_1 FILLER_52_1178 ();
 sg13g2_fill_1 FILLER_52_1188 ();
 sg13g2_fill_2 FILLER_52_1251 ();
 sg13g2_fill_1 FILLER_52_1253 ();
 sg13g2_decap_4 FILLER_52_1312 ();
 sg13g2_decap_4 FILLER_52_1350 ();
 sg13g2_decap_4 FILLER_52_1360 ();
 sg13g2_fill_1 FILLER_52_1364 ();
 sg13g2_fill_1 FILLER_52_1385 ();
 sg13g2_decap_8 FILLER_52_1390 ();
 sg13g2_decap_8 FILLER_52_1397 ();
 sg13g2_decap_8 FILLER_52_1404 ();
 sg13g2_fill_2 FILLER_52_1411 ();
 sg13g2_fill_1 FILLER_52_1413 ();
 sg13g2_fill_2 FILLER_52_1429 ();
 sg13g2_fill_2 FILLER_52_1446 ();
 sg13g2_decap_8 FILLER_52_1459 ();
 sg13g2_decap_8 FILLER_52_1466 ();
 sg13g2_decap_8 FILLER_52_1473 ();
 sg13g2_decap_8 FILLER_52_1480 ();
 sg13g2_fill_1 FILLER_52_1487 ();
 sg13g2_fill_2 FILLER_52_1492 ();
 sg13g2_decap_8 FILLER_52_1528 ();
 sg13g2_fill_2 FILLER_52_1535 ();
 sg13g2_decap_4 FILLER_52_1546 ();
 sg13g2_fill_2 FILLER_52_1563 ();
 sg13g2_fill_1 FILLER_52_1608 ();
 sg13g2_decap_8 FILLER_52_1621 ();
 sg13g2_decap_8 FILLER_52_1628 ();
 sg13g2_decap_4 FILLER_52_1635 ();
 sg13g2_fill_1 FILLER_52_1639 ();
 sg13g2_decap_8 FILLER_52_1670 ();
 sg13g2_fill_1 FILLER_52_1681 ();
 sg13g2_fill_1 FILLER_52_1688 ();
 sg13g2_fill_1 FILLER_52_1720 ();
 sg13g2_decap_8 FILLER_52_1760 ();
 sg13g2_decap_8 FILLER_52_1767 ();
 sg13g2_decap_4 FILLER_52_1774 ();
 sg13g2_fill_2 FILLER_52_1778 ();
 sg13g2_decap_8 FILLER_52_1786 ();
 sg13g2_decap_8 FILLER_52_1793 ();
 sg13g2_decap_8 FILLER_52_1800 ();
 sg13g2_decap_4 FILLER_52_1812 ();
 sg13g2_fill_1 FILLER_52_1816 ();
 sg13g2_decap_4 FILLER_52_1830 ();
 sg13g2_fill_1 FILLER_52_1834 ();
 sg13g2_fill_2 FILLER_52_1839 ();
 sg13g2_decap_4 FILLER_52_1872 ();
 sg13g2_fill_2 FILLER_52_1876 ();
 sg13g2_decap_8 FILLER_52_1888 ();
 sg13g2_decap_8 FILLER_52_1895 ();
 sg13g2_decap_8 FILLER_52_1902 ();
 sg13g2_decap_4 FILLER_52_1909 ();
 sg13g2_fill_2 FILLER_52_1913 ();
 sg13g2_decap_8 FILLER_52_1967 ();
 sg13g2_fill_2 FILLER_52_1979 ();
 sg13g2_fill_2 FILLER_52_2011 ();
 sg13g2_fill_1 FILLER_52_2013 ();
 sg13g2_decap_8 FILLER_52_2086 ();
 sg13g2_decap_8 FILLER_52_2093 ();
 sg13g2_decap_4 FILLER_52_2100 ();
 sg13g2_fill_2 FILLER_52_2104 ();
 sg13g2_decap_8 FILLER_52_2142 ();
 sg13g2_fill_2 FILLER_52_2149 ();
 sg13g2_fill_1 FILLER_52_2151 ();
 sg13g2_decap_8 FILLER_52_2156 ();
 sg13g2_decap_8 FILLER_52_2163 ();
 sg13g2_decap_8 FILLER_52_2170 ();
 sg13g2_decap_8 FILLER_52_2177 ();
 sg13g2_decap_8 FILLER_52_2184 ();
 sg13g2_decap_8 FILLER_52_2191 ();
 sg13g2_fill_2 FILLER_52_2211 ();
 sg13g2_fill_1 FILLER_52_2213 ();
 sg13g2_decap_4 FILLER_52_2240 ();
 sg13g2_fill_1 FILLER_52_2244 ();
 sg13g2_fill_2 FILLER_52_2258 ();
 sg13g2_fill_1 FILLER_52_2260 ();
 sg13g2_decap_8 FILLER_52_2292 ();
 sg13g2_fill_2 FILLER_52_2299 ();
 sg13g2_fill_2 FILLER_52_2314 ();
 sg13g2_decap_4 FILLER_52_2327 ();
 sg13g2_fill_2 FILLER_52_2336 ();
 sg13g2_decap_4 FILLER_52_2370 ();
 sg13g2_decap_4 FILLER_52_2383 ();
 sg13g2_fill_1 FILLER_52_2387 ();
 sg13g2_decap_4 FILLER_52_2414 ();
 sg13g2_fill_2 FILLER_52_2423 ();
 sg13g2_fill_1 FILLER_52_2425 ();
 sg13g2_fill_2 FILLER_52_2430 ();
 sg13g2_fill_1 FILLER_52_2432 ();
 sg13g2_decap_4 FILLER_52_2437 ();
 sg13g2_fill_2 FILLER_52_2441 ();
 sg13g2_decap_8 FILLER_52_2460 ();
 sg13g2_decap_4 FILLER_52_2467 ();
 sg13g2_fill_2 FILLER_52_2508 ();
 sg13g2_decap_8 FILLER_52_2540 ();
 sg13g2_decap_8 FILLER_52_2547 ();
 sg13g2_decap_8 FILLER_52_2554 ();
 sg13g2_decap_8 FILLER_52_2561 ();
 sg13g2_decap_8 FILLER_52_2568 ();
 sg13g2_decap_8 FILLER_52_2575 ();
 sg13g2_decap_8 FILLER_52_2582 ();
 sg13g2_decap_8 FILLER_52_2589 ();
 sg13g2_decap_8 FILLER_52_2596 ();
 sg13g2_decap_8 FILLER_52_2603 ();
 sg13g2_decap_8 FILLER_52_2610 ();
 sg13g2_decap_8 FILLER_52_2617 ();
 sg13g2_decap_8 FILLER_52_2624 ();
 sg13g2_decap_8 FILLER_52_2631 ();
 sg13g2_decap_8 FILLER_52_2638 ();
 sg13g2_decap_8 FILLER_52_2645 ();
 sg13g2_decap_8 FILLER_52_2652 ();
 sg13g2_decap_8 FILLER_52_2659 ();
 sg13g2_decap_4 FILLER_52_2666 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_40 ();
 sg13g2_fill_1 FILLER_53_57 ();
 sg13g2_fill_1 FILLER_53_62 ();
 sg13g2_fill_1 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_76 ();
 sg13g2_fill_2 FILLER_53_82 ();
 sg13g2_decap_8 FILLER_53_97 ();
 sg13g2_decap_8 FILLER_53_104 ();
 sg13g2_decap_8 FILLER_53_137 ();
 sg13g2_decap_4 FILLER_53_144 ();
 sg13g2_decap_4 FILLER_53_174 ();
 sg13g2_decap_8 FILLER_53_183 ();
 sg13g2_decap_4 FILLER_53_190 ();
 sg13g2_fill_1 FILLER_53_194 ();
 sg13g2_decap_8 FILLER_53_206 ();
 sg13g2_decap_8 FILLER_53_213 ();
 sg13g2_decap_4 FILLER_53_220 ();
 sg13g2_fill_2 FILLER_53_224 ();
 sg13g2_decap_4 FILLER_53_229 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_decap_8 FILLER_53_237 ();
 sg13g2_fill_2 FILLER_53_244 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_decap_4 FILLER_53_252 ();
 sg13g2_fill_2 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_267 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_fill_1 FILLER_53_297 ();
 sg13g2_fill_1 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_307 ();
 sg13g2_fill_2 FILLER_53_313 ();
 sg13g2_fill_2 FILLER_53_318 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_340 ();
 sg13g2_decap_8 FILLER_53_347 ();
 sg13g2_decap_8 FILLER_53_373 ();
 sg13g2_fill_2 FILLER_53_380 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_fill_2 FILLER_53_387 ();
 sg13g2_fill_1 FILLER_53_389 ();
 sg13g2_decap_4 FILLER_53_394 ();
 sg13g2_fill_1 FILLER_53_398 ();
 sg13g2_fill_2 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_53_405 ();
 sg13g2_decap_4 FILLER_53_411 ();
 sg13g2_fill_1 FILLER_53_415 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_fill_1 FILLER_53_428 ();
 sg13g2_fill_2 FILLER_53_433 ();
 sg13g2_fill_1 FILLER_53_435 ();
 sg13g2_decap_8 FILLER_53_459 ();
 sg13g2_decap_8 FILLER_53_466 ();
 sg13g2_decap_8 FILLER_53_473 ();
 sg13g2_decap_8 FILLER_53_480 ();
 sg13g2_decap_4 FILLER_53_487 ();
 sg13g2_fill_2 FILLER_53_491 ();
 sg13g2_fill_1 FILLER_53_516 ();
 sg13g2_fill_1 FILLER_53_521 ();
 sg13g2_fill_2 FILLER_53_527 ();
 sg13g2_fill_2 FILLER_53_533 ();
 sg13g2_fill_2 FILLER_53_539 ();
 sg13g2_fill_1 FILLER_53_541 ();
 sg13g2_decap_8 FILLER_53_547 ();
 sg13g2_decap_8 FILLER_53_554 ();
 sg13g2_decap_4 FILLER_53_561 ();
 sg13g2_decap_8 FILLER_53_573 ();
 sg13g2_fill_2 FILLER_53_584 ();
 sg13g2_decap_8 FILLER_53_619 ();
 sg13g2_fill_2 FILLER_53_626 ();
 sg13g2_fill_1 FILLER_53_638 ();
 sg13g2_fill_1 FILLER_53_674 ();
 sg13g2_fill_2 FILLER_53_679 ();
 sg13g2_fill_2 FILLER_53_686 ();
 sg13g2_fill_1 FILLER_53_706 ();
 sg13g2_fill_2 FILLER_53_737 ();
 sg13g2_fill_1 FILLER_53_739 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_fill_2 FILLER_53_779 ();
 sg13g2_decap_8 FILLER_53_810 ();
 sg13g2_decap_8 FILLER_53_835 ();
 sg13g2_fill_1 FILLER_53_842 ();
 sg13g2_fill_2 FILLER_53_851 ();
 sg13g2_decap_4 FILLER_53_862 ();
 sg13g2_fill_2 FILLER_53_866 ();
 sg13g2_decap_4 FILLER_53_872 ();
 sg13g2_decap_8 FILLER_53_907 ();
 sg13g2_fill_2 FILLER_53_914 ();
 sg13g2_decap_8 FILLER_53_942 ();
 sg13g2_decap_8 FILLER_53_949 ();
 sg13g2_decap_4 FILLER_53_960 ();
 sg13g2_fill_1 FILLER_53_964 ();
 sg13g2_decap_8 FILLER_53_971 ();
 sg13g2_decap_8 FILLER_53_978 ();
 sg13g2_decap_8 FILLER_53_985 ();
 sg13g2_fill_2 FILLER_53_992 ();
 sg13g2_fill_1 FILLER_53_994 ();
 sg13g2_decap_8 FILLER_53_1033 ();
 sg13g2_fill_2 FILLER_53_1040 ();
 sg13g2_fill_1 FILLER_53_1042 ();
 sg13g2_decap_8 FILLER_53_1049 ();
 sg13g2_decap_8 FILLER_53_1056 ();
 sg13g2_fill_2 FILLER_53_1086 ();
 sg13g2_fill_1 FILLER_53_1098 ();
 sg13g2_fill_2 FILLER_53_1111 ();
 sg13g2_fill_2 FILLER_53_1127 ();
 sg13g2_decap_4 FILLER_53_1136 ();
 sg13g2_fill_2 FILLER_53_1146 ();
 sg13g2_fill_1 FILLER_53_1148 ();
 sg13g2_fill_2 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1163 ();
 sg13g2_fill_1 FILLER_53_1170 ();
 sg13g2_fill_1 FILLER_53_1179 ();
 sg13g2_fill_2 FILLER_53_1222 ();
 sg13g2_fill_1 FILLER_53_1224 ();
 sg13g2_fill_1 FILLER_53_1236 ();
 sg13g2_fill_1 FILLER_53_1243 ();
 sg13g2_decap_4 FILLER_53_1250 ();
 sg13g2_fill_1 FILLER_53_1267 ();
 sg13g2_fill_2 FILLER_53_1274 ();
 sg13g2_fill_2 FILLER_53_1282 ();
 sg13g2_fill_1 FILLER_53_1284 ();
 sg13g2_fill_2 FILLER_53_1316 ();
 sg13g2_decap_8 FILLER_53_1334 ();
 sg13g2_fill_1 FILLER_53_1341 ();
 sg13g2_fill_2 FILLER_53_1377 ();
 sg13g2_fill_1 FILLER_53_1422 ();
 sg13g2_fill_1 FILLER_53_1487 ();
 sg13g2_fill_2 FILLER_53_1493 ();
 sg13g2_fill_1 FILLER_53_1499 ();
 sg13g2_fill_2 FILLER_53_1505 ();
 sg13g2_fill_1 FILLER_53_1507 ();
 sg13g2_decap_8 FILLER_53_1521 ();
 sg13g2_decap_8 FILLER_53_1528 ();
 sg13g2_decap_4 FILLER_53_1548 ();
 sg13g2_fill_1 FILLER_53_1593 ();
 sg13g2_decap_8 FILLER_53_1620 ();
 sg13g2_fill_1 FILLER_53_1627 ();
 sg13g2_fill_2 FILLER_53_1634 ();
 sg13g2_fill_1 FILLER_53_1636 ();
 sg13g2_fill_2 FILLER_53_1641 ();
 sg13g2_fill_1 FILLER_53_1643 ();
 sg13g2_decap_4 FILLER_53_1650 ();
 sg13g2_fill_2 FILLER_53_1654 ();
 sg13g2_decap_4 FILLER_53_1661 ();
 sg13g2_decap_8 FILLER_53_1671 ();
 sg13g2_decap_4 FILLER_53_1678 ();
 sg13g2_fill_1 FILLER_53_1682 ();
 sg13g2_decap_8 FILLER_53_1709 ();
 sg13g2_decap_8 FILLER_53_1716 ();
 sg13g2_fill_2 FILLER_53_1760 ();
 sg13g2_fill_1 FILLER_53_1762 ();
 sg13g2_decap_4 FILLER_53_1768 ();
 sg13g2_decap_8 FILLER_53_1776 ();
 sg13g2_decap_8 FILLER_53_1783 ();
 sg13g2_decap_4 FILLER_53_1822 ();
 sg13g2_fill_2 FILLER_53_1866 ();
 sg13g2_fill_1 FILLER_53_1868 ();
 sg13g2_fill_1 FILLER_53_1905 ();
 sg13g2_fill_1 FILLER_53_1932 ();
 sg13g2_fill_1 FILLER_53_1937 ();
 sg13g2_fill_1 FILLER_53_1969 ();
 sg13g2_decap_8 FILLER_53_1996 ();
 sg13g2_decap_8 FILLER_53_2003 ();
 sg13g2_decap_4 FILLER_53_2010 ();
 sg13g2_fill_1 FILLER_53_2014 ();
 sg13g2_fill_2 FILLER_53_2060 ();
 sg13g2_fill_1 FILLER_53_2062 ();
 sg13g2_fill_1 FILLER_53_2089 ();
 sg13g2_fill_2 FILLER_53_2095 ();
 sg13g2_fill_2 FILLER_53_2101 ();
 sg13g2_fill_1 FILLER_53_2103 ();
 sg13g2_fill_2 FILLER_53_2130 ();
 sg13g2_fill_1 FILLER_53_2132 ();
 sg13g2_fill_2 FILLER_53_2137 ();
 sg13g2_fill_2 FILLER_53_2148 ();
 sg13g2_fill_1 FILLER_53_2153 ();
 sg13g2_decap_8 FILLER_53_2180 ();
 sg13g2_decap_4 FILLER_53_2187 ();
 sg13g2_fill_2 FILLER_53_2191 ();
 sg13g2_fill_1 FILLER_53_2228 ();
 sg13g2_fill_1 FILLER_53_2233 ();
 sg13g2_fill_2 FILLER_53_2240 ();
 sg13g2_fill_1 FILLER_53_2268 ();
 sg13g2_decap_8 FILLER_53_2297 ();
 sg13g2_decap_8 FILLER_53_2304 ();
 sg13g2_decap_8 FILLER_53_2311 ();
 sg13g2_decap_8 FILLER_53_2318 ();
 sg13g2_decap_8 FILLER_53_2325 ();
 sg13g2_fill_1 FILLER_53_2332 ();
 sg13g2_decap_4 FILLER_53_2337 ();
 sg13g2_fill_1 FILLER_53_2341 ();
 sg13g2_decap_8 FILLER_53_2348 ();
 sg13g2_decap_8 FILLER_53_2355 ();
 sg13g2_decap_4 FILLER_53_2362 ();
 sg13g2_fill_1 FILLER_53_2366 ();
 sg13g2_decap_8 FILLER_53_2376 ();
 sg13g2_decap_8 FILLER_53_2383 ();
 sg13g2_decap_8 FILLER_53_2390 ();
 sg13g2_decap_8 FILLER_53_2397 ();
 sg13g2_decap_8 FILLER_53_2404 ();
 sg13g2_decap_8 FILLER_53_2411 ();
 sg13g2_decap_8 FILLER_53_2418 ();
 sg13g2_decap_8 FILLER_53_2425 ();
 sg13g2_decap_8 FILLER_53_2432 ();
 sg13g2_decap_8 FILLER_53_2439 ();
 sg13g2_decap_8 FILLER_53_2446 ();
 sg13g2_decap_8 FILLER_53_2453 ();
 sg13g2_fill_1 FILLER_53_2460 ();
 sg13g2_fill_2 FILLER_53_2466 ();
 sg13g2_fill_2 FILLER_53_2472 ();
 sg13g2_fill_2 FILLER_53_2479 ();
 sg13g2_fill_2 FILLER_53_2507 ();
 sg13g2_decap_4 FILLER_53_2519 ();
 sg13g2_fill_2 FILLER_53_2527 ();
 sg13g2_decap_8 FILLER_53_2565 ();
 sg13g2_decap_8 FILLER_53_2572 ();
 sg13g2_decap_8 FILLER_53_2579 ();
 sg13g2_decap_8 FILLER_53_2586 ();
 sg13g2_decap_8 FILLER_53_2593 ();
 sg13g2_decap_8 FILLER_53_2600 ();
 sg13g2_decap_8 FILLER_53_2607 ();
 sg13g2_decap_8 FILLER_53_2614 ();
 sg13g2_decap_8 FILLER_53_2621 ();
 sg13g2_decap_8 FILLER_53_2628 ();
 sg13g2_decap_8 FILLER_53_2635 ();
 sg13g2_decap_8 FILLER_53_2642 ();
 sg13g2_decap_8 FILLER_53_2649 ();
 sg13g2_decap_8 FILLER_53_2656 ();
 sg13g2_decap_8 FILLER_53_2663 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_37 ();
 sg13g2_fill_1 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_59 ();
 sg13g2_fill_2 FILLER_54_64 ();
 sg13g2_fill_1 FILLER_54_66 ();
 sg13g2_decap_8 FILLER_54_97 ();
 sg13g2_decap_8 FILLER_54_104 ();
 sg13g2_decap_8 FILLER_54_111 ();
 sg13g2_decap_8 FILLER_54_118 ();
 sg13g2_decap_8 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_150 ();
 sg13g2_fill_2 FILLER_54_177 ();
 sg13g2_fill_1 FILLER_54_216 ();
 sg13g2_decap_8 FILLER_54_221 ();
 sg13g2_fill_1 FILLER_54_228 ();
 sg13g2_decap_8 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_267 ();
 sg13g2_decap_8 FILLER_54_272 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_decap_8 FILLER_54_289 ();
 sg13g2_fill_2 FILLER_54_296 ();
 sg13g2_fill_1 FILLER_54_298 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_decap_8 FILLER_54_342 ();
 sg13g2_decap_4 FILLER_54_349 ();
 sg13g2_fill_1 FILLER_54_353 ();
 sg13g2_decap_8 FILLER_54_358 ();
 sg13g2_decap_4 FILLER_54_365 ();
 sg13g2_fill_2 FILLER_54_409 ();
 sg13g2_fill_1 FILLER_54_411 ();
 sg13g2_fill_2 FILLER_54_422 ();
 sg13g2_fill_1 FILLER_54_433 ();
 sg13g2_fill_1 FILLER_54_438 ();
 sg13g2_fill_1 FILLER_54_445 ();
 sg13g2_fill_1 FILLER_54_451 ();
 sg13g2_fill_2 FILLER_54_463 ();
 sg13g2_fill_1 FILLER_54_465 ();
 sg13g2_decap_4 FILLER_54_470 ();
 sg13g2_fill_2 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_fill_1 FILLER_54_509 ();
 sg13g2_fill_1 FILLER_54_515 ();
 sg13g2_fill_1 FILLER_54_526 ();
 sg13g2_decap_8 FILLER_54_546 ();
 sg13g2_decap_8 FILLER_54_553 ();
 sg13g2_decap_8 FILLER_54_560 ();
 sg13g2_fill_2 FILLER_54_567 ();
 sg13g2_fill_1 FILLER_54_589 ();
 sg13g2_decap_4 FILLER_54_633 ();
 sg13g2_fill_1 FILLER_54_641 ();
 sg13g2_fill_1 FILLER_54_655 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_fill_2 FILLER_54_713 ();
 sg13g2_fill_1 FILLER_54_741 ();
 sg13g2_fill_1 FILLER_54_748 ();
 sg13g2_fill_1 FILLER_54_781 ();
 sg13g2_decap_8 FILLER_54_818 ();
 sg13g2_decap_4 FILLER_54_851 ();
 sg13g2_fill_1 FILLER_54_855 ();
 sg13g2_fill_2 FILLER_54_861 ();
 sg13g2_fill_1 FILLER_54_863 ();
 sg13g2_fill_2 FILLER_54_890 ();
 sg13g2_fill_2 FILLER_54_897 ();
 sg13g2_fill_1 FILLER_54_899 ();
 sg13g2_fill_2 FILLER_54_905 ();
 sg13g2_fill_1 FILLER_54_907 ();
 sg13g2_fill_2 FILLER_54_934 ();
 sg13g2_decap_8 FILLER_54_966 ();
 sg13g2_decap_4 FILLER_54_973 ();
 sg13g2_fill_1 FILLER_54_977 ();
 sg13g2_decap_8 FILLER_54_984 ();
 sg13g2_decap_4 FILLER_54_991 ();
 sg13g2_fill_2 FILLER_54_995 ();
 sg13g2_decap_8 FILLER_54_1018 ();
 sg13g2_decap_8 FILLER_54_1025 ();
 sg13g2_fill_2 FILLER_54_1032 ();
 sg13g2_fill_1 FILLER_54_1034 ();
 sg13g2_fill_2 FILLER_54_1090 ();
 sg13g2_fill_1 FILLER_54_1098 ();
 sg13g2_fill_2 FILLER_54_1163 ();
 sg13g2_fill_2 FILLER_54_1169 ();
 sg13g2_fill_2 FILLER_54_1177 ();
 sg13g2_fill_1 FILLER_54_1179 ();
 sg13g2_fill_2 FILLER_54_1186 ();
 sg13g2_fill_1 FILLER_54_1188 ();
 sg13g2_fill_2 FILLER_54_1195 ();
 sg13g2_fill_1 FILLER_54_1197 ();
 sg13g2_decap_4 FILLER_54_1202 ();
 sg13g2_fill_2 FILLER_54_1206 ();
 sg13g2_decap_8 FILLER_54_1222 ();
 sg13g2_fill_1 FILLER_54_1229 ();
 sg13g2_decap_4 FILLER_54_1236 ();
 sg13g2_fill_2 FILLER_54_1240 ();
 sg13g2_decap_4 FILLER_54_1275 ();
 sg13g2_fill_1 FILLER_54_1279 ();
 sg13g2_fill_1 FILLER_54_1291 ();
 sg13g2_fill_1 FILLER_54_1302 ();
 sg13g2_decap_4 FILLER_54_1312 ();
 sg13g2_fill_2 FILLER_54_1316 ();
 sg13g2_fill_2 FILLER_54_1323 ();
 sg13g2_fill_1 FILLER_54_1325 ();
 sg13g2_fill_2 FILLER_54_1352 ();
 sg13g2_fill_1 FILLER_54_1357 ();
 sg13g2_fill_1 FILLER_54_1361 ();
 sg13g2_fill_2 FILLER_54_1379 ();
 sg13g2_fill_1 FILLER_54_1419 ();
 sg13g2_fill_1 FILLER_54_1427 ();
 sg13g2_fill_2 FILLER_54_1448 ();
 sg13g2_fill_2 FILLER_54_1462 ();
 sg13g2_fill_2 FILLER_54_1469 ();
 sg13g2_fill_2 FILLER_54_1497 ();
 sg13g2_decap_8 FILLER_54_1535 ();
 sg13g2_decap_4 FILLER_54_1542 ();
 sg13g2_fill_1 FILLER_54_1546 ();
 sg13g2_decap_8 FILLER_54_1552 ();
 sg13g2_decap_8 FILLER_54_1559 ();
 sg13g2_decap_4 FILLER_54_1626 ();
 sg13g2_fill_2 FILLER_54_1630 ();
 sg13g2_fill_1 FILLER_54_1637 ();
 sg13g2_decap_4 FILLER_54_1662 ();
 sg13g2_fill_2 FILLER_54_1666 ();
 sg13g2_decap_4 FILLER_54_1672 ();
 sg13g2_fill_1 FILLER_54_1676 ();
 sg13g2_fill_2 FILLER_54_1683 ();
 sg13g2_fill_1 FILLER_54_1685 ();
 sg13g2_fill_2 FILLER_54_1691 ();
 sg13g2_decap_4 FILLER_54_1702 ();
 sg13g2_fill_2 FILLER_54_1710 ();
 sg13g2_fill_2 FILLER_54_1743 ();
 sg13g2_decap_8 FILLER_54_1749 ();
 sg13g2_fill_1 FILLER_54_1756 ();
 sg13g2_decap_8 FILLER_54_1786 ();
 sg13g2_decap_8 FILLER_54_1793 ();
 sg13g2_decap_4 FILLER_54_1800 ();
 sg13g2_fill_2 FILLER_54_1804 ();
 sg13g2_fill_1 FILLER_54_1815 ();
 sg13g2_fill_2 FILLER_54_1842 ();
 sg13g2_fill_1 FILLER_54_1889 ();
 sg13g2_fill_1 FILLER_54_1895 ();
 sg13g2_decap_8 FILLER_54_1902 ();
 sg13g2_fill_2 FILLER_54_1909 ();
 sg13g2_fill_1 FILLER_54_1911 ();
 sg13g2_fill_1 FILLER_54_1917 ();
 sg13g2_fill_2 FILLER_54_1927 ();
 sg13g2_fill_1 FILLER_54_1934 ();
 sg13g2_fill_2 FILLER_54_1939 ();
 sg13g2_fill_2 FILLER_54_2010 ();
 sg13g2_fill_1 FILLER_54_2012 ();
 sg13g2_fill_2 FILLER_54_2039 ();
 sg13g2_fill_1 FILLER_54_2041 ();
 sg13g2_fill_2 FILLER_54_2085 ();
 sg13g2_decap_8 FILLER_54_2123 ();
 sg13g2_decap_4 FILLER_54_2130 ();
 sg13g2_fill_2 FILLER_54_2147 ();
 sg13g2_fill_1 FILLER_54_2149 ();
 sg13g2_decap_4 FILLER_54_2159 ();
 sg13g2_fill_1 FILLER_54_2163 ();
 sg13g2_decap_4 FILLER_54_2170 ();
 sg13g2_fill_2 FILLER_54_2174 ();
 sg13g2_fill_2 FILLER_54_2282 ();
 sg13g2_fill_1 FILLER_54_2284 ();
 sg13g2_decap_4 FILLER_54_2298 ();
 sg13g2_fill_1 FILLER_54_2302 ();
 sg13g2_fill_1 FILLER_54_2309 ();
 sg13g2_fill_2 FILLER_54_2336 ();
 sg13g2_fill_2 FILLER_54_2344 ();
 sg13g2_fill_2 FILLER_54_2372 ();
 sg13g2_decap_8 FILLER_54_2400 ();
 sg13g2_decap_4 FILLER_54_2407 ();
 sg13g2_decap_4 FILLER_54_2419 ();
 sg13g2_decap_4 FILLER_54_2435 ();
 sg13g2_fill_2 FILLER_54_2469 ();
 sg13g2_decap_8 FILLER_54_2518 ();
 sg13g2_decap_8 FILLER_54_2525 ();
 sg13g2_decap_8 FILLER_54_2532 ();
 sg13g2_decap_4 FILLER_54_2539 ();
 sg13g2_fill_1 FILLER_54_2543 ();
 sg13g2_decap_8 FILLER_54_2548 ();
 sg13g2_decap_8 FILLER_54_2555 ();
 sg13g2_decap_8 FILLER_54_2562 ();
 sg13g2_decap_8 FILLER_54_2569 ();
 sg13g2_decap_8 FILLER_54_2576 ();
 sg13g2_decap_8 FILLER_54_2583 ();
 sg13g2_decap_8 FILLER_54_2590 ();
 sg13g2_decap_8 FILLER_54_2597 ();
 sg13g2_decap_8 FILLER_54_2604 ();
 sg13g2_decap_8 FILLER_54_2611 ();
 sg13g2_decap_8 FILLER_54_2618 ();
 sg13g2_decap_8 FILLER_54_2625 ();
 sg13g2_decap_8 FILLER_54_2632 ();
 sg13g2_decap_8 FILLER_54_2639 ();
 sg13g2_decap_8 FILLER_54_2646 ();
 sg13g2_decap_8 FILLER_54_2653 ();
 sg13g2_decap_8 FILLER_54_2660 ();
 sg13g2_fill_2 FILLER_54_2667 ();
 sg13g2_fill_1 FILLER_54_2669 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_4 FILLER_55_56 ();
 sg13g2_fill_1 FILLER_55_60 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_fill_1 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_159 ();
 sg13g2_decap_4 FILLER_55_166 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_187 ();
 sg13g2_decap_8 FILLER_55_204 ();
 sg13g2_fill_1 FILLER_55_211 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_4 FILLER_55_224 ();
 sg13g2_fill_1 FILLER_55_254 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_289 ();
 sg13g2_fill_2 FILLER_55_295 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_2 FILLER_55_321 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_fill_1 FILLER_55_347 ();
 sg13g2_fill_1 FILLER_55_371 ();
 sg13g2_fill_1 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_398 ();
 sg13g2_fill_1 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_411 ();
 sg13g2_fill_1 FILLER_55_417 ();
 sg13g2_fill_1 FILLER_55_422 ();
 sg13g2_fill_1 FILLER_55_437 ();
 sg13g2_fill_2 FILLER_55_461 ();
 sg13g2_fill_2 FILLER_55_486 ();
 sg13g2_fill_1 FILLER_55_493 ();
 sg13g2_fill_2 FILLER_55_502 ();
 sg13g2_fill_2 FILLER_55_512 ();
 sg13g2_fill_1 FILLER_55_514 ();
 sg13g2_fill_2 FILLER_55_525 ();
 sg13g2_decap_8 FILLER_55_531 ();
 sg13g2_fill_1 FILLER_55_538 ();
 sg13g2_decap_4 FILLER_55_544 ();
 sg13g2_fill_1 FILLER_55_548 ();
 sg13g2_decap_8 FILLER_55_564 ();
 sg13g2_fill_1 FILLER_55_575 ();
 sg13g2_fill_1 FILLER_55_581 ();
 sg13g2_fill_1 FILLER_55_587 ();
 sg13g2_decap_4 FILLER_55_593 ();
 sg13g2_fill_2 FILLER_55_597 ();
 sg13g2_fill_2 FILLER_55_607 ();
 sg13g2_fill_1 FILLER_55_623 ();
 sg13g2_fill_2 FILLER_55_637 ();
 sg13g2_fill_1 FILLER_55_651 ();
 sg13g2_decap_8 FILLER_55_662 ();
 sg13g2_decap_4 FILLER_55_669 ();
 sg13g2_fill_1 FILLER_55_673 ();
 sg13g2_fill_2 FILLER_55_686 ();
 sg13g2_fill_2 FILLER_55_702 ();
 sg13g2_fill_1 FILLER_55_744 ();
 sg13g2_decap_8 FILLER_55_782 ();
 sg13g2_decap_8 FILLER_55_789 ();
 sg13g2_decap_8 FILLER_55_796 ();
 sg13g2_decap_8 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_810 ();
 sg13g2_fill_1 FILLER_55_817 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_decap_4 FILLER_55_835 ();
 sg13g2_fill_1 FILLER_55_839 ();
 sg13g2_decap_8 FILLER_55_866 ();
 sg13g2_decap_8 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_55_884 ();
 sg13g2_decap_8 FILLER_55_891 ();
 sg13g2_fill_1 FILLER_55_898 ();
 sg13g2_decap_8 FILLER_55_934 ();
 sg13g2_decap_8 FILLER_55_941 ();
 sg13g2_fill_2 FILLER_55_948 ();
 sg13g2_fill_1 FILLER_55_950 ();
 sg13g2_fill_2 FILLER_55_1018 ();
 sg13g2_fill_1 FILLER_55_1020 ();
 sg13g2_fill_2 FILLER_55_1026 ();
 sg13g2_fill_1 FILLER_55_1028 ();
 sg13g2_decap_4 FILLER_55_1033 ();
 sg13g2_decap_8 FILLER_55_1041 ();
 sg13g2_decap_8 FILLER_55_1053 ();
 sg13g2_decap_8 FILLER_55_1060 ();
 sg13g2_fill_2 FILLER_55_1067 ();
 sg13g2_fill_1 FILLER_55_1085 ();
 sg13g2_fill_1 FILLER_55_1091 ();
 sg13g2_fill_2 FILLER_55_1100 ();
 sg13g2_fill_1 FILLER_55_1108 ();
 sg13g2_fill_2 FILLER_55_1113 ();
 sg13g2_fill_2 FILLER_55_1131 ();
 sg13g2_decap_4 FILLER_55_1139 ();
 sg13g2_fill_1 FILLER_55_1143 ();
 sg13g2_fill_2 FILLER_55_1183 ();
 sg13g2_fill_1 FILLER_55_1191 ();
 sg13g2_fill_1 FILLER_55_1229 ();
 sg13g2_fill_2 FILLER_55_1245 ();
 sg13g2_fill_1 FILLER_55_1247 ();
 sg13g2_decap_8 FILLER_55_1273 ();
 sg13g2_fill_2 FILLER_55_1280 ();
 sg13g2_decap_8 FILLER_55_1321 ();
 sg13g2_decap_8 FILLER_55_1328 ();
 sg13g2_decap_4 FILLER_55_1335 ();
 sg13g2_fill_2 FILLER_55_1343 ();
 sg13g2_fill_2 FILLER_55_1362 ();
 sg13g2_fill_2 FILLER_55_1405 ();
 sg13g2_fill_2 FILLER_55_1411 ();
 sg13g2_decap_8 FILLER_55_1484 ();
 sg13g2_decap_8 FILLER_55_1491 ();
 sg13g2_fill_1 FILLER_55_1498 ();
 sg13g2_decap_8 FILLER_55_1504 ();
 sg13g2_decap_8 FILLER_55_1511 ();
 sg13g2_fill_2 FILLER_55_1518 ();
 sg13g2_fill_2 FILLER_55_1535 ();
 sg13g2_decap_8 FILLER_55_1541 ();
 sg13g2_decap_8 FILLER_55_1553 ();
 sg13g2_decap_4 FILLER_55_1560 ();
 sg13g2_fill_2 FILLER_55_1587 ();
 sg13g2_fill_2 FILLER_55_1615 ();
 sg13g2_fill_1 FILLER_55_1617 ();
 sg13g2_fill_2 FILLER_55_1650 ();
 sg13g2_decap_8 FILLER_55_1678 ();
 sg13g2_fill_2 FILLER_55_1685 ();
 sg13g2_fill_1 FILLER_55_1693 ();
 sg13g2_decap_4 FILLER_55_1720 ();
 sg13g2_fill_1 FILLER_55_1724 ();
 sg13g2_fill_2 FILLER_55_1743 ();
 sg13g2_fill_2 FILLER_55_1791 ();
 sg13g2_decap_4 FILLER_55_1801 ();
 sg13g2_fill_1 FILLER_55_1805 ();
 sg13g2_fill_2 FILLER_55_1810 ();
 sg13g2_decap_4 FILLER_55_1818 ();
 sg13g2_decap_4 FILLER_55_1827 ();
 sg13g2_fill_1 FILLER_55_1864 ();
 sg13g2_decap_8 FILLER_55_1913 ();
 sg13g2_decap_8 FILLER_55_1920 ();
 sg13g2_decap_4 FILLER_55_1932 ();
 sg13g2_fill_2 FILLER_55_1936 ();
 sg13g2_fill_1 FILLER_55_1950 ();
 sg13g2_decap_8 FILLER_55_1959 ();
 sg13g2_fill_1 FILLER_55_1966 ();
 sg13g2_fill_2 FILLER_55_1973 ();
 sg13g2_fill_1 FILLER_55_1987 ();
 sg13g2_decap_4 FILLER_55_1993 ();
 sg13g2_fill_2 FILLER_55_1997 ();
 sg13g2_fill_2 FILLER_55_2005 ();
 sg13g2_fill_1 FILLER_55_2007 ();
 sg13g2_fill_1 FILLER_55_2014 ();
 sg13g2_fill_2 FILLER_55_2020 ();
 sg13g2_fill_1 FILLER_55_2022 ();
 sg13g2_decap_8 FILLER_55_2027 ();
 sg13g2_decap_4 FILLER_55_2034 ();
 sg13g2_decap_8 FILLER_55_2071 ();
 sg13g2_decap_8 FILLER_55_2078 ();
 sg13g2_decap_8 FILLER_55_2085 ();
 sg13g2_decap_4 FILLER_55_2102 ();
 sg13g2_decap_4 FILLER_55_2132 ();
 sg13g2_decap_4 FILLER_55_2162 ();
 sg13g2_decap_8 FILLER_55_2179 ();
 sg13g2_fill_2 FILLER_55_2194 ();
 sg13g2_fill_2 FILLER_55_2237 ();
 sg13g2_fill_2 FILLER_55_2244 ();
 sg13g2_fill_2 FILLER_55_2250 ();
 sg13g2_fill_1 FILLER_55_2252 ();
 sg13g2_decap_8 FILLER_55_2262 ();
 sg13g2_decap_8 FILLER_55_2269 ();
 sg13g2_fill_2 FILLER_55_2276 ();
 sg13g2_fill_1 FILLER_55_2278 ();
 sg13g2_fill_1 FILLER_55_2284 ();
 sg13g2_decap_8 FILLER_55_2290 ();
 sg13g2_decap_8 FILLER_55_2310 ();
 sg13g2_decap_4 FILLER_55_2317 ();
 sg13g2_fill_2 FILLER_55_2321 ();
 sg13g2_fill_1 FILLER_55_2360 ();
 sg13g2_decap_4 FILLER_55_2365 ();
 sg13g2_decap_4 FILLER_55_2374 ();
 sg13g2_fill_2 FILLER_55_2378 ();
 sg13g2_fill_2 FILLER_55_2406 ();
 sg13g2_fill_2 FILLER_55_2412 ();
 sg13g2_fill_2 FILLER_55_2469 ();
 sg13g2_fill_1 FILLER_55_2481 ();
 sg13g2_decap_8 FILLER_55_2513 ();
 sg13g2_decap_8 FILLER_55_2520 ();
 sg13g2_decap_8 FILLER_55_2527 ();
 sg13g2_fill_1 FILLER_55_2534 ();
 sg13g2_decap_8 FILLER_55_2565 ();
 sg13g2_decap_8 FILLER_55_2572 ();
 sg13g2_decap_8 FILLER_55_2579 ();
 sg13g2_decap_8 FILLER_55_2586 ();
 sg13g2_decap_8 FILLER_55_2593 ();
 sg13g2_decap_8 FILLER_55_2600 ();
 sg13g2_decap_8 FILLER_55_2607 ();
 sg13g2_decap_8 FILLER_55_2614 ();
 sg13g2_decap_8 FILLER_55_2621 ();
 sg13g2_decap_8 FILLER_55_2628 ();
 sg13g2_decap_8 FILLER_55_2635 ();
 sg13g2_decap_8 FILLER_55_2642 ();
 sg13g2_decap_8 FILLER_55_2649 ();
 sg13g2_decap_8 FILLER_55_2656 ();
 sg13g2_decap_8 FILLER_55_2663 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_4 FILLER_56_84 ();
 sg13g2_fill_2 FILLER_56_88 ();
 sg13g2_decap_8 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_101 ();
 sg13g2_decap_8 FILLER_56_108 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_decap_8 FILLER_56_122 ();
 sg13g2_decap_8 FILLER_56_129 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_150 ();
 sg13g2_decap_8 FILLER_56_157 ();
 sg13g2_decap_8 FILLER_56_164 ();
 sg13g2_decap_8 FILLER_56_171 ();
 sg13g2_decap_8 FILLER_56_178 ();
 sg13g2_decap_8 FILLER_56_185 ();
 sg13g2_decap_8 FILLER_56_192 ();
 sg13g2_decap_8 FILLER_56_199 ();
 sg13g2_decap_8 FILLER_56_206 ();
 sg13g2_decap_8 FILLER_56_213 ();
 sg13g2_decap_8 FILLER_56_220 ();
 sg13g2_decap_4 FILLER_56_227 ();
 sg13g2_fill_2 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_236 ();
 sg13g2_decap_8 FILLER_56_243 ();
 sg13g2_decap_4 FILLER_56_250 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_fill_1 FILLER_56_350 ();
 sg13g2_fill_2 FILLER_56_355 ();
 sg13g2_fill_1 FILLER_56_365 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_4 FILLER_56_424 ();
 sg13g2_fill_1 FILLER_56_428 ();
 sg13g2_fill_1 FILLER_56_441 ();
 sg13g2_fill_2 FILLER_56_446 ();
 sg13g2_fill_2 FILLER_56_457 ();
 sg13g2_fill_1 FILLER_56_463 ();
 sg13g2_fill_1 FILLER_56_469 ();
 sg13g2_fill_1 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_485 ();
 sg13g2_fill_2 FILLER_56_490 ();
 sg13g2_decap_8 FILLER_56_513 ();
 sg13g2_fill_2 FILLER_56_520 ();
 sg13g2_fill_2 FILLER_56_527 ();
 sg13g2_fill_2 FILLER_56_534 ();
 sg13g2_fill_1 FILLER_56_536 ();
 sg13g2_fill_1 FILLER_56_554 ();
 sg13g2_fill_1 FILLER_56_560 ();
 sg13g2_fill_2 FILLER_56_569 ();
 sg13g2_fill_2 FILLER_56_576 ();
 sg13g2_fill_2 FILLER_56_584 ();
 sg13g2_fill_1 FILLER_56_606 ();
 sg13g2_decap_8 FILLER_56_617 ();
 sg13g2_fill_2 FILLER_56_634 ();
 sg13g2_fill_2 FILLER_56_672 ();
 sg13g2_fill_1 FILLER_56_685 ();
 sg13g2_fill_2 FILLER_56_728 ();
 sg13g2_fill_2 FILLER_56_759 ();
 sg13g2_decap_8 FILLER_56_776 ();
 sg13g2_decap_8 FILLER_56_783 ();
 sg13g2_decap_8 FILLER_56_790 ();
 sg13g2_decap_8 FILLER_56_797 ();
 sg13g2_decap_4 FILLER_56_822 ();
 sg13g2_fill_2 FILLER_56_826 ();
 sg13g2_fill_1 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_864 ();
 sg13g2_decap_4 FILLER_56_913 ();
 sg13g2_decap_8 FILLER_56_921 ();
 sg13g2_decap_8 FILLER_56_928 ();
 sg13g2_decap_8 FILLER_56_935 ();
 sg13g2_fill_1 FILLER_56_942 ();
 sg13g2_decap_8 FILLER_56_956 ();
 sg13g2_decap_8 FILLER_56_963 ();
 sg13g2_fill_1 FILLER_56_970 ();
 sg13g2_decap_8 FILLER_56_976 ();
 sg13g2_decap_4 FILLER_56_997 ();
 sg13g2_fill_1 FILLER_56_1001 ();
 sg13g2_decap_8 FILLER_56_1006 ();
 sg13g2_fill_1 FILLER_56_1048 ();
 sg13g2_fill_2 FILLER_56_1059 ();
 sg13g2_decap_4 FILLER_56_1067 ();
 sg13g2_decap_4 FILLER_56_1079 ();
 sg13g2_fill_2 FILLER_56_1089 ();
 sg13g2_fill_1 FILLER_56_1091 ();
 sg13g2_fill_2 FILLER_56_1112 ();
 sg13g2_fill_1 FILLER_56_1114 ();
 sg13g2_decap_4 FILLER_56_1126 ();
 sg13g2_fill_2 FILLER_56_1182 ();
 sg13g2_fill_1 FILLER_56_1190 ();
 sg13g2_fill_1 FILLER_56_1196 ();
 sg13g2_decap_8 FILLER_56_1208 ();
 sg13g2_fill_1 FILLER_56_1215 ();
 sg13g2_fill_1 FILLER_56_1220 ();
 sg13g2_decap_4 FILLER_56_1238 ();
 sg13g2_fill_1 FILLER_56_1242 ();
 sg13g2_fill_1 FILLER_56_1252 ();
 sg13g2_fill_2 FILLER_56_1279 ();
 sg13g2_fill_1 FILLER_56_1281 ();
 sg13g2_fill_2 FILLER_56_1288 ();
 sg13g2_fill_1 FILLER_56_1290 ();
 sg13g2_fill_1 FILLER_56_1317 ();
 sg13g2_fill_2 FILLER_56_1324 ();
 sg13g2_fill_2 FILLER_56_1383 ();
 sg13g2_fill_1 FILLER_56_1397 ();
 sg13g2_decap_8 FILLER_56_1458 ();
 sg13g2_decap_8 FILLER_56_1465 ();
 sg13g2_decap_4 FILLER_56_1472 ();
 sg13g2_fill_2 FILLER_56_1476 ();
 sg13g2_decap_8 FILLER_56_1489 ();
 sg13g2_decap_8 FILLER_56_1496 ();
 sg13g2_decap_8 FILLER_56_1503 ();
 sg13g2_decap_8 FILLER_56_1510 ();
 sg13g2_decap_4 FILLER_56_1517 ();
 sg13g2_decap_8 FILLER_56_1545 ();
 sg13g2_decap_8 FILLER_56_1552 ();
 sg13g2_decap_8 FILLER_56_1559 ();
 sg13g2_decap_4 FILLER_56_1566 ();
 sg13g2_fill_2 FILLER_56_1570 ();
 sg13g2_decap_8 FILLER_56_1575 ();
 sg13g2_decap_4 FILLER_56_1582 ();
 sg13g2_fill_2 FILLER_56_1586 ();
 sg13g2_fill_1 FILLER_56_1614 ();
 sg13g2_decap_4 FILLER_56_1618 ();
 sg13g2_decap_8 FILLER_56_1648 ();
 sg13g2_decap_4 FILLER_56_1655 ();
 sg13g2_fill_2 FILLER_56_1659 ();
 sg13g2_decap_4 FILLER_56_1713 ();
 sg13g2_fill_1 FILLER_56_1717 ();
 sg13g2_fill_1 FILLER_56_1722 ();
 sg13g2_decap_8 FILLER_56_1726 ();
 sg13g2_fill_2 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1748 ();
 sg13g2_fill_2 FILLER_56_1755 ();
 sg13g2_fill_2 FILLER_56_1766 ();
 sg13g2_decap_4 FILLER_56_1773 ();
 sg13g2_fill_1 FILLER_56_1777 ();
 sg13g2_fill_1 FILLER_56_1783 ();
 sg13g2_decap_4 FILLER_56_1819 ();
 sg13g2_fill_2 FILLER_56_1823 ();
 sg13g2_fill_2 FILLER_56_1849 ();
 sg13g2_fill_2 FILLER_56_1882 ();
 sg13g2_fill_1 FILLER_56_1884 ();
 sg13g2_decap_4 FILLER_56_1895 ();
 sg13g2_fill_1 FILLER_56_1899 ();
 sg13g2_decap_8 FILLER_56_1917 ();
 sg13g2_decap_8 FILLER_56_1924 ();
 sg13g2_fill_2 FILLER_56_1931 ();
 sg13g2_decap_8 FILLER_56_1950 ();
 sg13g2_decap_8 FILLER_56_1957 ();
 sg13g2_decap_8 FILLER_56_1964 ();
 sg13g2_decap_4 FILLER_56_1971 ();
 sg13g2_fill_2 FILLER_56_1980 ();
 sg13g2_decap_4 FILLER_56_1996 ();
 sg13g2_fill_1 FILLER_56_2000 ();
 sg13g2_decap_8 FILLER_56_2007 ();
 sg13g2_decap_8 FILLER_56_2014 ();
 sg13g2_decap_4 FILLER_56_2021 ();
 sg13g2_fill_1 FILLER_56_2025 ();
 sg13g2_decap_4 FILLER_56_2031 ();
 sg13g2_fill_1 FILLER_56_2035 ();
 sg13g2_decap_8 FILLER_56_2040 ();
 sg13g2_fill_2 FILLER_56_2047 ();
 sg13g2_fill_1 FILLER_56_2049 ();
 sg13g2_decap_8 FILLER_56_2055 ();
 sg13g2_decap_4 FILLER_56_2062 ();
 sg13g2_fill_2 FILLER_56_2066 ();
 sg13g2_fill_1 FILLER_56_2082 ();
 sg13g2_decap_4 FILLER_56_2093 ();
 sg13g2_fill_1 FILLER_56_2097 ();
 sg13g2_fill_1 FILLER_56_2108 ();
 sg13g2_decap_8 FILLER_56_2113 ();
 sg13g2_fill_2 FILLER_56_2120 ();
 sg13g2_fill_1 FILLER_56_2122 ();
 sg13g2_fill_2 FILLER_56_2131 ();
 sg13g2_fill_2 FILLER_56_2138 ();
 sg13g2_fill_1 FILLER_56_2140 ();
 sg13g2_fill_2 FILLER_56_2172 ();
 sg13g2_decap_4 FILLER_56_2187 ();
 sg13g2_decap_8 FILLER_56_2207 ();
 sg13g2_decap_8 FILLER_56_2214 ();
 sg13g2_decap_4 FILLER_56_2221 ();
 sg13g2_fill_1 FILLER_56_2225 ();
 sg13g2_fill_2 FILLER_56_2229 ();
 sg13g2_fill_1 FILLER_56_2231 ();
 sg13g2_decap_8 FILLER_56_2237 ();
 sg13g2_decap_8 FILLER_56_2244 ();
 sg13g2_decap_8 FILLER_56_2251 ();
 sg13g2_decap_4 FILLER_56_2258 ();
 sg13g2_fill_2 FILLER_56_2262 ();
 sg13g2_decap_4 FILLER_56_2277 ();
 sg13g2_fill_1 FILLER_56_2281 ();
 sg13g2_decap_8 FILLER_56_2308 ();
 sg13g2_fill_2 FILLER_56_2315 ();
 sg13g2_fill_1 FILLER_56_2322 ();
 sg13g2_decap_8 FILLER_56_2329 ();
 sg13g2_decap_4 FILLER_56_2350 ();
 sg13g2_decap_8 FILLER_56_2362 ();
 sg13g2_decap_8 FILLER_56_2369 ();
 sg13g2_fill_1 FILLER_56_2376 ();
 sg13g2_decap_8 FILLER_56_2381 ();
 sg13g2_decap_8 FILLER_56_2388 ();
 sg13g2_fill_2 FILLER_56_2405 ();
 sg13g2_fill_1 FILLER_56_2407 ();
 sg13g2_fill_2 FILLER_56_2412 ();
 sg13g2_fill_1 FILLER_56_2440 ();
 sg13g2_fill_1 FILLER_56_2491 ();
 sg13g2_fill_1 FILLER_56_2496 ();
 sg13g2_decap_4 FILLER_56_2505 ();
 sg13g2_fill_1 FILLER_56_2509 ();
 sg13g2_decap_8 FILLER_56_2514 ();
 sg13g2_fill_1 FILLER_56_2521 ();
 sg13g2_decap_4 FILLER_56_2532 ();
 sg13g2_decap_4 FILLER_56_2540 ();
 sg13g2_fill_2 FILLER_56_2544 ();
 sg13g2_decap_8 FILLER_56_2550 ();
 sg13g2_decap_8 FILLER_56_2557 ();
 sg13g2_decap_8 FILLER_56_2564 ();
 sg13g2_decap_8 FILLER_56_2571 ();
 sg13g2_decap_8 FILLER_56_2578 ();
 sg13g2_decap_8 FILLER_56_2585 ();
 sg13g2_decap_8 FILLER_56_2592 ();
 sg13g2_decap_8 FILLER_56_2599 ();
 sg13g2_decap_8 FILLER_56_2606 ();
 sg13g2_decap_8 FILLER_56_2613 ();
 sg13g2_decap_8 FILLER_56_2620 ();
 sg13g2_decap_8 FILLER_56_2627 ();
 sg13g2_decap_8 FILLER_56_2634 ();
 sg13g2_decap_8 FILLER_56_2641 ();
 sg13g2_decap_8 FILLER_56_2648 ();
 sg13g2_decap_8 FILLER_56_2655 ();
 sg13g2_decap_8 FILLER_56_2662 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_21 ();
 sg13g2_decap_4 FILLER_57_26 ();
 sg13g2_decap_4 FILLER_57_34 ();
 sg13g2_fill_2 FILLER_57_45 ();
 sg13g2_fill_1 FILLER_57_47 ();
 sg13g2_decap_4 FILLER_57_52 ();
 sg13g2_fill_2 FILLER_57_56 ();
 sg13g2_decap_4 FILLER_57_62 ();
 sg13g2_decap_4 FILLER_57_74 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_130 ();
 sg13g2_decap_8 FILLER_57_136 ();
 sg13g2_decap_8 FILLER_57_143 ();
 sg13g2_decap_8 FILLER_57_150 ();
 sg13g2_decap_8 FILLER_57_157 ();
 sg13g2_decap_8 FILLER_57_164 ();
 sg13g2_decap_8 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_178 ();
 sg13g2_fill_2 FILLER_57_185 ();
 sg13g2_fill_1 FILLER_57_187 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_decap_8 FILLER_57_225 ();
 sg13g2_fill_2 FILLER_57_232 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_decap_8 FILLER_57_239 ();
 sg13g2_decap_8 FILLER_57_246 ();
 sg13g2_decap_8 FILLER_57_253 ();
 sg13g2_decap_8 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_311 ();
 sg13g2_decap_8 FILLER_57_318 ();
 sg13g2_decap_8 FILLER_57_325 ();
 sg13g2_decap_8 FILLER_57_332 ();
 sg13g2_decap_4 FILLER_57_339 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_decap_8 FILLER_57_363 ();
 sg13g2_fill_2 FILLER_57_370 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_decap_4 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_decap_8 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_57_414 ();
 sg13g2_decap_4 FILLER_57_421 ();
 sg13g2_fill_1 FILLER_57_425 ();
 sg13g2_decap_8 FILLER_57_436 ();
 sg13g2_fill_1 FILLER_57_443 ();
 sg13g2_decap_4 FILLER_57_448 ();
 sg13g2_decap_4 FILLER_57_456 ();
 sg13g2_fill_2 FILLER_57_460 ();
 sg13g2_fill_2 FILLER_57_467 ();
 sg13g2_decap_4 FILLER_57_473 ();
 sg13g2_fill_2 FILLER_57_477 ();
 sg13g2_fill_2 FILLER_57_484 ();
 sg13g2_fill_1 FILLER_57_486 ();
 sg13g2_fill_2 FILLER_57_492 ();
 sg13g2_fill_1 FILLER_57_494 ();
 sg13g2_fill_2 FILLER_57_499 ();
 sg13g2_fill_1 FILLER_57_501 ();
 sg13g2_decap_8 FILLER_57_507 ();
 sg13g2_decap_8 FILLER_57_514 ();
 sg13g2_decap_8 FILLER_57_521 ();
 sg13g2_decap_8 FILLER_57_528 ();
 sg13g2_fill_1 FILLER_57_535 ();
 sg13g2_fill_1 FILLER_57_551 ();
 sg13g2_decap_8 FILLER_57_564 ();
 sg13g2_fill_2 FILLER_57_571 ();
 sg13g2_decap_8 FILLER_57_580 ();
 sg13g2_fill_1 FILLER_57_606 ();
 sg13g2_fill_2 FILLER_57_618 ();
 sg13g2_fill_1 FILLER_57_620 ();
 sg13g2_fill_2 FILLER_57_640 ();
 sg13g2_fill_1 FILLER_57_642 ();
 sg13g2_fill_2 FILLER_57_646 ();
 sg13g2_decap_8 FILLER_57_652 ();
 sg13g2_fill_2 FILLER_57_659 ();
 sg13g2_decap_8 FILLER_57_666 ();
 sg13g2_decap_8 FILLER_57_673 ();
 sg13g2_fill_1 FILLER_57_680 ();
 sg13g2_decap_4 FILLER_57_686 ();
 sg13g2_fill_2 FILLER_57_698 ();
 sg13g2_fill_1 FILLER_57_700 ();
 sg13g2_decap_4 FILLER_57_709 ();
 sg13g2_fill_2 FILLER_57_717 ();
 sg13g2_fill_1 FILLER_57_723 ();
 sg13g2_decap_8 FILLER_57_732 ();
 sg13g2_decap_4 FILLER_57_739 ();
 sg13g2_fill_1 FILLER_57_743 ();
 sg13g2_decap_8 FILLER_57_771 ();
 sg13g2_decap_8 FILLER_57_778 ();
 sg13g2_decap_4 FILLER_57_785 ();
 sg13g2_fill_1 FILLER_57_789 ();
 sg13g2_decap_8 FILLER_57_816 ();
 sg13g2_decap_8 FILLER_57_823 ();
 sg13g2_fill_2 FILLER_57_830 ();
 sg13g2_fill_1 FILLER_57_832 ();
 sg13g2_fill_2 FILLER_57_838 ();
 sg13g2_fill_1 FILLER_57_840 ();
 sg13g2_decap_8 FILLER_57_876 ();
 sg13g2_decap_4 FILLER_57_883 ();
 sg13g2_decap_8 FILLER_57_913 ();
 sg13g2_decap_8 FILLER_57_920 ();
 sg13g2_fill_1 FILLER_57_927 ();
 sg13g2_fill_2 FILLER_57_962 ();
 sg13g2_fill_1 FILLER_57_968 ();
 sg13g2_decap_8 FILLER_57_973 ();
 sg13g2_decap_8 FILLER_57_980 ();
 sg13g2_decap_8 FILLER_57_987 ();
 sg13g2_fill_1 FILLER_57_994 ();
 sg13g2_fill_2 FILLER_57_1025 ();
 sg13g2_fill_1 FILLER_57_1065 ();
 sg13g2_fill_2 FILLER_57_1071 ();
 sg13g2_fill_1 FILLER_57_1073 ();
 sg13g2_fill_2 FILLER_57_1105 ();
 sg13g2_fill_1 FILLER_57_1107 ();
 sg13g2_fill_1 FILLER_57_1142 ();
 sg13g2_decap_4 FILLER_57_1147 ();
 sg13g2_fill_2 FILLER_57_1151 ();
 sg13g2_fill_1 FILLER_57_1182 ();
 sg13g2_decap_4 FILLER_57_1203 ();
 sg13g2_fill_2 FILLER_57_1207 ();
 sg13g2_decap_4 FILLER_57_1235 ();
 sg13g2_fill_1 FILLER_57_1239 ();
 sg13g2_fill_1 FILLER_57_1255 ();
 sg13g2_fill_2 FILLER_57_1282 ();
 sg13g2_fill_1 FILLER_57_1284 ();
 sg13g2_fill_1 FILLER_57_1317 ();
 sg13g2_decap_8 FILLER_57_1364 ();
 sg13g2_decap_4 FILLER_57_1371 ();
 sg13g2_fill_1 FILLER_57_1375 ();
 sg13g2_fill_1 FILLER_57_1411 ();
 sg13g2_fill_1 FILLER_57_1470 ();
 sg13g2_fill_2 FILLER_57_1475 ();
 sg13g2_fill_1 FILLER_57_1477 ();
 sg13g2_decap_4 FILLER_57_1483 ();
 sg13g2_fill_1 FILLER_57_1487 ();
 sg13g2_decap_8 FILLER_57_1492 ();
 sg13g2_decap_8 FILLER_57_1499 ();
 sg13g2_decap_8 FILLER_57_1506 ();
 sg13g2_decap_8 FILLER_57_1526 ();
 sg13g2_fill_2 FILLER_57_1551 ();
 sg13g2_fill_1 FILLER_57_1553 ();
 sg13g2_decap_4 FILLER_57_1567 ();
 sg13g2_fill_1 FILLER_57_1571 ();
 sg13g2_decap_8 FILLER_57_1579 ();
 sg13g2_decap_8 FILLER_57_1586 ();
 sg13g2_decap_8 FILLER_57_1593 ();
 sg13g2_decap_4 FILLER_57_1600 ();
 sg13g2_fill_2 FILLER_57_1604 ();
 sg13g2_fill_2 FILLER_57_1618 ();
 sg13g2_decap_8 FILLER_57_1659 ();
 sg13g2_decap_8 FILLER_57_1666 ();
 sg13g2_decap_8 FILLER_57_1682 ();
 sg13g2_decap_8 FILLER_57_1689 ();
 sg13g2_decap_8 FILLER_57_1696 ();
 sg13g2_fill_2 FILLER_57_1709 ();
 sg13g2_fill_1 FILLER_57_1711 ();
 sg13g2_fill_2 FILLER_57_1717 ();
 sg13g2_fill_1 FILLER_57_1719 ();
 sg13g2_decap_4 FILLER_57_1731 ();
 sg13g2_fill_2 FILLER_57_1785 ();
 sg13g2_fill_1 FILLER_57_1829 ();
 sg13g2_fill_2 FILLER_57_1887 ();
 sg13g2_fill_1 FILLER_57_1889 ();
 sg13g2_decap_8 FILLER_57_1896 ();
 sg13g2_fill_2 FILLER_57_1903 ();
 sg13g2_fill_1 FILLER_57_1905 ();
 sg13g2_fill_2 FILLER_57_1932 ();
 sg13g2_decap_8 FILLER_57_1964 ();
 sg13g2_decap_8 FILLER_57_1971 ();
 sg13g2_decap_8 FILLER_57_1978 ();
 sg13g2_decap_4 FILLER_57_2015 ();
 sg13g2_fill_1 FILLER_57_2027 ();
 sg13g2_decap_8 FILLER_57_2058 ();
 sg13g2_decap_8 FILLER_57_2098 ();
 sg13g2_decap_4 FILLER_57_2105 ();
 sg13g2_decap_8 FILLER_57_2113 ();
 sg13g2_fill_2 FILLER_57_2120 ();
 sg13g2_fill_2 FILLER_57_2126 ();
 sg13g2_fill_1 FILLER_57_2128 ();
 sg13g2_fill_2 FILLER_57_2163 ();
 sg13g2_decap_8 FILLER_57_2171 ();
 sg13g2_decap_8 FILLER_57_2178 ();
 sg13g2_decap_8 FILLER_57_2185 ();
 sg13g2_decap_8 FILLER_57_2192 ();
 sg13g2_decap_8 FILLER_57_2199 ();
 sg13g2_fill_2 FILLER_57_2206 ();
 sg13g2_fill_1 FILLER_57_2208 ();
 sg13g2_decap_8 FILLER_57_2218 ();
 sg13g2_fill_1 FILLER_57_2225 ();
 sg13g2_fill_1 FILLER_57_2231 ();
 sg13g2_fill_2 FILLER_57_2267 ();
 sg13g2_fill_1 FILLER_57_2269 ();
 sg13g2_fill_1 FILLER_57_2296 ();
 sg13g2_fill_2 FILLER_57_2305 ();
 sg13g2_fill_1 FILLER_57_2307 ();
 sg13g2_fill_1 FILLER_57_2360 ();
 sg13g2_decap_8 FILLER_57_2367 ();
 sg13g2_decap_4 FILLER_57_2374 ();
 sg13g2_fill_1 FILLER_57_2413 ();
 sg13g2_decap_8 FILLER_57_2440 ();
 sg13g2_fill_2 FILLER_57_2447 ();
 sg13g2_fill_1 FILLER_57_2449 ();
 sg13g2_decap_4 FILLER_57_2454 ();
 sg13g2_fill_2 FILLER_57_2458 ();
 sg13g2_fill_1 FILLER_57_2480 ();
 sg13g2_fill_2 FILLER_57_2497 ();
 sg13g2_decap_8 FILLER_57_2555 ();
 sg13g2_decap_8 FILLER_57_2562 ();
 sg13g2_decap_8 FILLER_57_2569 ();
 sg13g2_decap_8 FILLER_57_2576 ();
 sg13g2_decap_8 FILLER_57_2583 ();
 sg13g2_decap_8 FILLER_57_2590 ();
 sg13g2_decap_8 FILLER_57_2597 ();
 sg13g2_decap_8 FILLER_57_2604 ();
 sg13g2_decap_8 FILLER_57_2611 ();
 sg13g2_decap_8 FILLER_57_2618 ();
 sg13g2_decap_8 FILLER_57_2625 ();
 sg13g2_decap_8 FILLER_57_2632 ();
 sg13g2_decap_8 FILLER_57_2639 ();
 sg13g2_decap_8 FILLER_57_2646 ();
 sg13g2_decap_8 FILLER_57_2653 ();
 sg13g2_decap_8 FILLER_57_2660 ();
 sg13g2_fill_2 FILLER_57_2667 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_11 ();
 sg13g2_fill_1 FILLER_58_58 ();
 sg13g2_fill_2 FILLER_58_68 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_146 ();
 sg13g2_decap_8 FILLER_58_151 ();
 sg13g2_decap_8 FILLER_58_158 ();
 sg13g2_fill_1 FILLER_58_165 ();
 sg13g2_decap_8 FILLER_58_171 ();
 sg13g2_fill_2 FILLER_58_178 ();
 sg13g2_decap_8 FILLER_58_184 ();
 sg13g2_decap_4 FILLER_58_199 ();
 sg13g2_fill_2 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_248 ();
 sg13g2_decap_8 FILLER_58_255 ();
 sg13g2_decap_8 FILLER_58_262 ();
 sg13g2_decap_8 FILLER_58_269 ();
 sg13g2_decap_8 FILLER_58_276 ();
 sg13g2_decap_8 FILLER_58_283 ();
 sg13g2_decap_8 FILLER_58_290 ();
 sg13g2_decap_8 FILLER_58_297 ();
 sg13g2_fill_2 FILLER_58_304 ();
 sg13g2_decap_8 FILLER_58_310 ();
 sg13g2_decap_8 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_decap_8 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_58_361 ();
 sg13g2_decap_8 FILLER_58_368 ();
 sg13g2_decap_4 FILLER_58_390 ();
 sg13g2_fill_2 FILLER_58_394 ();
 sg13g2_fill_1 FILLER_58_410 ();
 sg13g2_fill_1 FILLER_58_415 ();
 sg13g2_fill_1 FILLER_58_421 ();
 sg13g2_decap_8 FILLER_58_430 ();
 sg13g2_decap_8 FILLER_58_437 ();
 sg13g2_decap_8 FILLER_58_444 ();
 sg13g2_fill_2 FILLER_58_455 ();
 sg13g2_fill_1 FILLER_58_457 ();
 sg13g2_fill_2 FILLER_58_468 ();
 sg13g2_fill_1 FILLER_58_470 ();
 sg13g2_fill_1 FILLER_58_476 ();
 sg13g2_fill_2 FILLER_58_482 ();
 sg13g2_decap_4 FILLER_58_494 ();
 sg13g2_fill_2 FILLER_58_509 ();
 sg13g2_fill_2 FILLER_58_516 ();
 sg13g2_decap_4 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_531 ();
 sg13g2_fill_2 FILLER_58_538 ();
 sg13g2_fill_1 FILLER_58_540 ();
 sg13g2_decap_8 FILLER_58_550 ();
 sg13g2_decap_4 FILLER_58_557 ();
 sg13g2_fill_2 FILLER_58_561 ();
 sg13g2_decap_8 FILLER_58_575 ();
 sg13g2_decap_8 FILLER_58_582 ();
 sg13g2_decap_8 FILLER_58_589 ();
 sg13g2_fill_2 FILLER_58_596 ();
 sg13g2_fill_1 FILLER_58_636 ();
 sg13g2_decap_8 FILLER_58_641 ();
 sg13g2_decap_8 FILLER_58_648 ();
 sg13g2_fill_1 FILLER_58_655 ();
 sg13g2_decap_8 FILLER_58_660 ();
 sg13g2_fill_2 FILLER_58_667 ();
 sg13g2_fill_2 FILLER_58_673 ();
 sg13g2_fill_1 FILLER_58_675 ();
 sg13g2_fill_1 FILLER_58_702 ();
 sg13g2_fill_1 FILLER_58_708 ();
 sg13g2_decap_8 FILLER_58_735 ();
 sg13g2_fill_2 FILLER_58_742 ();
 sg13g2_fill_1 FILLER_58_744 ();
 sg13g2_fill_2 FILLER_58_751 ();
 sg13g2_fill_2 FILLER_58_761 ();
 sg13g2_fill_1 FILLER_58_763 ();
 sg13g2_fill_1 FILLER_58_769 ();
 sg13g2_decap_4 FILLER_58_815 ();
 sg13g2_fill_1 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_4 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_844 ();
 sg13g2_fill_1 FILLER_58_851 ();
 sg13g2_decap_8 FILLER_58_864 ();
 sg13g2_decap_8 FILLER_58_871 ();
 sg13g2_decap_8 FILLER_58_878 ();
 sg13g2_decap_8 FILLER_58_885 ();
 sg13g2_decap_8 FILLER_58_892 ();
 sg13g2_decap_4 FILLER_58_899 ();
 sg13g2_fill_1 FILLER_58_903 ();
 sg13g2_decap_4 FILLER_58_914 ();
 sg13g2_fill_1 FILLER_58_918 ();
 sg13g2_fill_2 FILLER_58_955 ();
 sg13g2_fill_2 FILLER_58_968 ();
 sg13g2_decap_8 FILLER_58_976 ();
 sg13g2_fill_2 FILLER_58_983 ();
 sg13g2_fill_2 FILLER_58_990 ();
 sg13g2_fill_1 FILLER_58_992 ();
 sg13g2_fill_1 FILLER_58_997 ();
 sg13g2_decap_4 FILLER_58_1003 ();
 sg13g2_fill_1 FILLER_58_1007 ();
 sg13g2_decap_4 FILLER_58_1013 ();
 sg13g2_fill_1 FILLER_58_1017 ();
 sg13g2_fill_1 FILLER_58_1067 ();
 sg13g2_decap_8 FILLER_58_1072 ();
 sg13g2_decap_8 FILLER_58_1079 ();
 sg13g2_decap_4 FILLER_58_1091 ();
 sg13g2_fill_2 FILLER_58_1095 ();
 sg13g2_fill_2 FILLER_58_1103 ();
 sg13g2_fill_1 FILLER_58_1105 ();
 sg13g2_fill_1 FILLER_58_1124 ();
 sg13g2_decap_8 FILLER_58_1129 ();
 sg13g2_fill_1 FILLER_58_1136 ();
 sg13g2_fill_2 FILLER_58_1204 ();
 sg13g2_decap_8 FILLER_58_1215 ();
 sg13g2_decap_8 FILLER_58_1222 ();
 sg13g2_decap_4 FILLER_58_1229 ();
 sg13g2_fill_1 FILLER_58_1233 ();
 sg13g2_fill_2 FILLER_58_1241 ();
 sg13g2_fill_1 FILLER_58_1243 ();
 sg13g2_fill_2 FILLER_58_1254 ();
 sg13g2_decap_8 FILLER_58_1265 ();
 sg13g2_decap_4 FILLER_58_1272 ();
 sg13g2_fill_1 FILLER_58_1285 ();
 sg13g2_fill_2 FILLER_58_1309 ();
 sg13g2_fill_1 FILLER_58_1316 ();
 sg13g2_fill_2 FILLER_58_1322 ();
 sg13g2_fill_1 FILLER_58_1328 ();
 sg13g2_fill_1 FILLER_58_1343 ();
 sg13g2_fill_2 FILLER_58_1349 ();
 sg13g2_decap_4 FILLER_58_1378 ();
 sg13g2_fill_1 FILLER_58_1382 ();
 sg13g2_fill_1 FILLER_58_1390 ();
 sg13g2_fill_2 FILLER_58_1444 ();
 sg13g2_fill_1 FILLER_58_1446 ();
 sg13g2_fill_1 FILLER_58_1509 ();
 sg13g2_decap_4 FILLER_58_1514 ();
 sg13g2_fill_2 FILLER_58_1518 ();
 sg13g2_fill_2 FILLER_58_1546 ();
 sg13g2_fill_1 FILLER_58_1548 ();
 sg13g2_fill_1 FILLER_58_1553 ();
 sg13g2_decap_4 FILLER_58_1584 ();
 sg13g2_fill_1 FILLER_58_1610 ();
 sg13g2_decap_8 FILLER_58_1616 ();
 sg13g2_decap_8 FILLER_58_1623 ();
 sg13g2_fill_2 FILLER_58_1630 ();
 sg13g2_decap_4 FILLER_58_1654 ();
 sg13g2_fill_2 FILLER_58_1658 ();
 sg13g2_fill_2 FILLER_58_1674 ();
 sg13g2_decap_8 FILLER_58_1684 ();
 sg13g2_fill_1 FILLER_58_1691 ();
 sg13g2_fill_2 FILLER_58_1701 ();
 sg13g2_decap_8 FILLER_58_1709 ();
 sg13g2_decap_4 FILLER_58_1716 ();
 sg13g2_fill_2 FILLER_58_1720 ();
 sg13g2_fill_1 FILLER_58_1731 ();
 sg13g2_decap_4 FILLER_58_1740 ();
 sg13g2_fill_1 FILLER_58_1744 ();
 sg13g2_fill_1 FILLER_58_1749 ();
 sg13g2_fill_2 FILLER_58_1816 ();
 sg13g2_fill_1 FILLER_58_1857 ();
 sg13g2_fill_2 FILLER_58_1870 ();
 sg13g2_decap_8 FILLER_58_1882 ();
 sg13g2_decap_8 FILLER_58_1889 ();
 sg13g2_decap_8 FILLER_58_1896 ();
 sg13g2_fill_1 FILLER_58_1903 ();
 sg13g2_fill_2 FILLER_58_1970 ();
 sg13g2_fill_1 FILLER_58_1990 ();
 sg13g2_fill_2 FILLER_58_1996 ();
 sg13g2_fill_1 FILLER_58_2003 ();
 sg13g2_fill_2 FILLER_58_2030 ();
 sg13g2_decap_4 FILLER_58_2038 ();
 sg13g2_fill_1 FILLER_58_2071 ();
 sg13g2_decap_4 FILLER_58_2080 ();
 sg13g2_decap_8 FILLER_58_2115 ();
 sg13g2_decap_8 FILLER_58_2122 ();
 sg13g2_fill_1 FILLER_58_2129 ();
 sg13g2_fill_2 FILLER_58_2138 ();
 sg13g2_fill_1 FILLER_58_2150 ();
 sg13g2_fill_2 FILLER_58_2155 ();
 sg13g2_fill_1 FILLER_58_2157 ();
 sg13g2_fill_1 FILLER_58_2170 ();
 sg13g2_fill_1 FILLER_58_2258 ();
 sg13g2_fill_2 FILLER_58_2265 ();
 sg13g2_fill_1 FILLER_58_2267 ();
 sg13g2_fill_1 FILLER_58_2299 ();
 sg13g2_fill_2 FILLER_58_2305 ();
 sg13g2_decap_4 FILLER_58_2320 ();
 sg13g2_fill_2 FILLER_58_2330 ();
 sg13g2_fill_1 FILLER_58_2332 ();
 sg13g2_decap_8 FILLER_58_2339 ();
 sg13g2_fill_2 FILLER_58_2356 ();
 sg13g2_fill_1 FILLER_58_2358 ();
 sg13g2_fill_2 FILLER_58_2368 ();
 sg13g2_fill_1 FILLER_58_2370 ();
 sg13g2_decap_4 FILLER_58_2375 ();
 sg13g2_fill_2 FILLER_58_2418 ();
 sg13g2_fill_1 FILLER_58_2420 ();
 sg13g2_decap_8 FILLER_58_2429 ();
 sg13g2_decap_8 FILLER_58_2436 ();
 sg13g2_decap_8 FILLER_58_2443 ();
 sg13g2_decap_8 FILLER_58_2450 ();
 sg13g2_fill_2 FILLER_58_2457 ();
 sg13g2_fill_1 FILLER_58_2535 ();
 sg13g2_decap_4 FILLER_58_2540 ();
 sg13g2_fill_1 FILLER_58_2544 ();
 sg13g2_decap_8 FILLER_58_2549 ();
 sg13g2_decap_8 FILLER_58_2556 ();
 sg13g2_decap_8 FILLER_58_2563 ();
 sg13g2_decap_8 FILLER_58_2570 ();
 sg13g2_decap_8 FILLER_58_2577 ();
 sg13g2_decap_8 FILLER_58_2584 ();
 sg13g2_decap_8 FILLER_58_2591 ();
 sg13g2_decap_8 FILLER_58_2598 ();
 sg13g2_decap_8 FILLER_58_2605 ();
 sg13g2_decap_8 FILLER_58_2612 ();
 sg13g2_decap_8 FILLER_58_2619 ();
 sg13g2_decap_8 FILLER_58_2626 ();
 sg13g2_decap_8 FILLER_58_2633 ();
 sg13g2_decap_8 FILLER_58_2640 ();
 sg13g2_decap_8 FILLER_58_2647 ();
 sg13g2_decap_8 FILLER_58_2654 ();
 sg13g2_decap_8 FILLER_58_2661 ();
 sg13g2_fill_2 FILLER_58_2668 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_2 FILLER_59_11 ();
 sg13g2_fill_1 FILLER_59_25 ();
 sg13g2_fill_1 FILLER_59_54 ();
 sg13g2_fill_2 FILLER_59_70 ();
 sg13g2_fill_2 FILLER_59_117 ();
 sg13g2_decap_4 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_decap_8 FILLER_59_188 ();
 sg13g2_decap_8 FILLER_59_195 ();
 sg13g2_decap_8 FILLER_59_206 ();
 sg13g2_fill_2 FILLER_59_248 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_4 FILLER_59_294 ();
 sg13g2_fill_2 FILLER_59_298 ();
 sg13g2_decap_8 FILLER_59_305 ();
 sg13g2_decap_8 FILLER_59_312 ();
 sg13g2_decap_8 FILLER_59_319 ();
 sg13g2_decap_8 FILLER_59_326 ();
 sg13g2_decap_8 FILLER_59_333 ();
 sg13g2_decap_8 FILLER_59_340 ();
 sg13g2_decap_8 FILLER_59_347 ();
 sg13g2_decap_8 FILLER_59_354 ();
 sg13g2_decap_8 FILLER_59_361 ();
 sg13g2_fill_2 FILLER_59_388 ();
 sg13g2_decap_4 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_59_409 ();
 sg13g2_fill_1 FILLER_59_421 ();
 sg13g2_fill_2 FILLER_59_448 ();
 sg13g2_fill_2 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_481 ();
 sg13g2_fill_1 FILLER_59_498 ();
 sg13g2_fill_2 FILLER_59_503 ();
 sg13g2_decap_4 FILLER_59_511 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_decap_8 FILLER_59_529 ();
 sg13g2_decap_4 FILLER_59_536 ();
 sg13g2_fill_2 FILLER_59_540 ();
 sg13g2_fill_1 FILLER_59_547 ();
 sg13g2_decap_8 FILLER_59_552 ();
 sg13g2_fill_2 FILLER_59_559 ();
 sg13g2_fill_1 FILLER_59_561 ();
 sg13g2_fill_2 FILLER_59_592 ();
 sg13g2_fill_2 FILLER_59_599 ();
 sg13g2_fill_1 FILLER_59_601 ();
 sg13g2_fill_2 FILLER_59_619 ();
 sg13g2_fill_2 FILLER_59_635 ();
 sg13g2_decap_8 FILLER_59_641 ();
 sg13g2_decap_4 FILLER_59_648 ();
 sg13g2_fill_1 FILLER_59_652 ();
 sg13g2_fill_2 FILLER_59_682 ();
 sg13g2_fill_1 FILLER_59_692 ();
 sg13g2_decap_8 FILLER_59_698 ();
 sg13g2_fill_2 FILLER_59_705 ();
 sg13g2_fill_1 FILLER_59_743 ();
 sg13g2_decap_8 FILLER_59_779 ();
 sg13g2_fill_2 FILLER_59_786 ();
 sg13g2_fill_1 FILLER_59_788 ();
 sg13g2_fill_2 FILLER_59_897 ();
 sg13g2_fill_2 FILLER_59_925 ();
 sg13g2_fill_1 FILLER_59_927 ();
 sg13g2_fill_2 FILLER_59_939 ();
 sg13g2_fill_1 FILLER_59_949 ();
 sg13g2_decap_4 FILLER_59_986 ();
 sg13g2_fill_2 FILLER_59_990 ();
 sg13g2_fill_2 FILLER_59_1010 ();
 sg13g2_fill_1 FILLER_59_1012 ();
 sg13g2_fill_2 FILLER_59_1019 ();
 sg13g2_fill_1 FILLER_59_1021 ();
 sg13g2_fill_2 FILLER_59_1027 ();
 sg13g2_fill_1 FILLER_59_1029 ();
 sg13g2_decap_4 FILLER_59_1038 ();
 sg13g2_fill_2 FILLER_59_1042 ();
 sg13g2_fill_1 FILLER_59_1066 ();
 sg13g2_decap_4 FILLER_59_1081 ();
 sg13g2_fill_1 FILLER_59_1085 ();
 sg13g2_fill_2 FILLER_59_1091 ();
 sg13g2_fill_1 FILLER_59_1103 ();
 sg13g2_fill_2 FILLER_59_1121 ();
 sg13g2_fill_1 FILLER_59_1123 ();
 sg13g2_decap_4 FILLER_59_1133 ();
 sg13g2_fill_1 FILLER_59_1137 ();
 sg13g2_decap_8 FILLER_59_1217 ();
 sg13g2_decap_8 FILLER_59_1224 ();
 sg13g2_decap_8 FILLER_59_1265 ();
 sg13g2_decap_8 FILLER_59_1277 ();
 sg13g2_decap_4 FILLER_59_1284 ();
 sg13g2_fill_2 FILLER_59_1288 ();
 sg13g2_fill_1 FILLER_59_1308 ();
 sg13g2_fill_2 FILLER_59_1335 ();
 sg13g2_decap_4 FILLER_59_1361 ();
 sg13g2_fill_1 FILLER_59_1365 ();
 sg13g2_decap_4 FILLER_59_1369 ();
 sg13g2_fill_1 FILLER_59_1373 ();
 sg13g2_decap_4 FILLER_59_1379 ();
 sg13g2_fill_1 FILLER_59_1387 ();
 sg13g2_fill_2 FILLER_59_1428 ();
 sg13g2_fill_2 FILLER_59_1460 ();
 sg13g2_fill_2 FILLER_59_1501 ();
 sg13g2_fill_1 FILLER_59_1503 ();
 sg13g2_fill_1 FILLER_59_1522 ();
 sg13g2_fill_2 FILLER_59_1578 ();
 sg13g2_decap_8 FILLER_59_1610 ();
 sg13g2_decap_8 FILLER_59_1617 ();
 sg13g2_decap_8 FILLER_59_1624 ();
 sg13g2_decap_8 FILLER_59_1631 ();
 sg13g2_decap_4 FILLER_59_1638 ();
 sg13g2_fill_2 FILLER_59_1642 ();
 sg13g2_decap_4 FILLER_59_1670 ();
 sg13g2_decap_8 FILLER_59_1700 ();
 sg13g2_decap_8 FILLER_59_1707 ();
 sg13g2_fill_1 FILLER_59_1714 ();
 sg13g2_fill_2 FILLER_59_1723 ();
 sg13g2_decap_4 FILLER_59_1762 ();
 sg13g2_fill_2 FILLER_59_1766 ();
 sg13g2_fill_2 FILLER_59_1787 ();
 sg13g2_decap_8 FILLER_59_1821 ();
 sg13g2_fill_2 FILLER_59_1828 ();
 sg13g2_decap_4 FILLER_59_1835 ();
 sg13g2_fill_1 FILLER_59_1839 ();
 sg13g2_fill_1 FILLER_59_1848 ();
 sg13g2_decap_8 FILLER_59_1880 ();
 sg13g2_decap_8 FILLER_59_1887 ();
 sg13g2_decap_8 FILLER_59_1894 ();
 sg13g2_decap_4 FILLER_59_1901 ();
 sg13g2_fill_1 FILLER_59_1905 ();
 sg13g2_decap_8 FILLER_59_1933 ();
 sg13g2_decap_8 FILLER_59_1940 ();
 sg13g2_decap_4 FILLER_59_2073 ();
 sg13g2_fill_1 FILLER_59_2077 ();
 sg13g2_fill_2 FILLER_59_2082 ();
 sg13g2_fill_1 FILLER_59_2098 ();
 sg13g2_decap_8 FILLER_59_2125 ();
 sg13g2_fill_2 FILLER_59_2132 ();
 sg13g2_decap_4 FILLER_59_2160 ();
 sg13g2_fill_2 FILLER_59_2177 ();
 sg13g2_decap_8 FILLER_59_2197 ();
 sg13g2_decap_8 FILLER_59_2204 ();
 sg13g2_decap_8 FILLER_59_2211 ();
 sg13g2_decap_4 FILLER_59_2218 ();
 sg13g2_fill_2 FILLER_59_2222 ();
 sg13g2_fill_2 FILLER_59_2277 ();
 sg13g2_fill_2 FILLER_59_2296 ();
 sg13g2_decap_4 FILLER_59_2303 ();
 sg13g2_fill_2 FILLER_59_2315 ();
 sg13g2_decap_4 FILLER_59_2333 ();
 sg13g2_fill_2 FILLER_59_2341 ();
 sg13g2_decap_4 FILLER_59_2348 ();
 sg13g2_fill_1 FILLER_59_2352 ();
 sg13g2_fill_1 FILLER_59_2358 ();
 sg13g2_decap_8 FILLER_59_2395 ();
 sg13g2_decap_8 FILLER_59_2402 ();
 sg13g2_decap_8 FILLER_59_2409 ();
 sg13g2_decap_8 FILLER_59_2416 ();
 sg13g2_decap_8 FILLER_59_2423 ();
 sg13g2_decap_8 FILLER_59_2430 ();
 sg13g2_decap_8 FILLER_59_2437 ();
 sg13g2_decap_4 FILLER_59_2444 ();
 sg13g2_fill_1 FILLER_59_2492 ();
 sg13g2_decap_8 FILLER_59_2523 ();
 sg13g2_decap_4 FILLER_59_2530 ();
 sg13g2_decap_8 FILLER_59_2564 ();
 sg13g2_decap_8 FILLER_59_2571 ();
 sg13g2_decap_8 FILLER_59_2578 ();
 sg13g2_decap_8 FILLER_59_2585 ();
 sg13g2_decap_8 FILLER_59_2592 ();
 sg13g2_decap_8 FILLER_59_2599 ();
 sg13g2_decap_8 FILLER_59_2606 ();
 sg13g2_decap_8 FILLER_59_2613 ();
 sg13g2_decap_8 FILLER_59_2620 ();
 sg13g2_decap_8 FILLER_59_2627 ();
 sg13g2_decap_8 FILLER_59_2634 ();
 sg13g2_decap_8 FILLER_59_2641 ();
 sg13g2_decap_8 FILLER_59_2648 ();
 sg13g2_decap_8 FILLER_59_2655 ();
 sg13g2_decap_8 FILLER_59_2662 ();
 sg13g2_fill_1 FILLER_59_2669 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_1 FILLER_60_55 ();
 sg13g2_decap_4 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_100 ();
 sg13g2_fill_1 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_122 ();
 sg13g2_fill_2 FILLER_60_129 ();
 sg13g2_fill_1 FILLER_60_156 ();
 sg13g2_fill_1 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_193 ();
 sg13g2_fill_2 FILLER_60_200 ();
 sg13g2_fill_1 FILLER_60_202 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_259 ();
 sg13g2_fill_2 FILLER_60_265 ();
 sg13g2_fill_1 FILLER_60_267 ();
 sg13g2_fill_1 FILLER_60_275 ();
 sg13g2_fill_2 FILLER_60_286 ();
 sg13g2_decap_4 FILLER_60_297 ();
 sg13g2_decap_8 FILLER_60_319 ();
 sg13g2_fill_2 FILLER_60_334 ();
 sg13g2_fill_1 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_363 ();
 sg13g2_fill_2 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_decap_4 FILLER_60_378 ();
 sg13g2_fill_1 FILLER_60_382 ();
 sg13g2_decap_4 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_60_413 ();
 sg13g2_decap_8 FILLER_60_420 ();
 sg13g2_decap_8 FILLER_60_427 ();
 sg13g2_fill_2 FILLER_60_434 ();
 sg13g2_decap_4 FILLER_60_480 ();
 sg13g2_fill_2 FILLER_60_484 ();
 sg13g2_decap_4 FILLER_60_490 ();
 sg13g2_fill_2 FILLER_60_494 ();
 sg13g2_fill_2 FILLER_60_507 ();
 sg13g2_decap_8 FILLER_60_522 ();
 sg13g2_decap_8 FILLER_60_529 ();
 sg13g2_fill_1 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_552 ();
 sg13g2_fill_1 FILLER_60_594 ();
 sg13g2_fill_1 FILLER_60_599 ();
 sg13g2_decap_4 FILLER_60_635 ();
 sg13g2_fill_1 FILLER_60_639 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_fill_2 FILLER_60_683 ();
 sg13g2_fill_1 FILLER_60_685 ();
 sg13g2_decap_8 FILLER_60_695 ();
 sg13g2_fill_2 FILLER_60_702 ();
 sg13g2_fill_1 FILLER_60_704 ();
 sg13g2_fill_2 FILLER_60_709 ();
 sg13g2_fill_1 FILLER_60_711 ();
 sg13g2_decap_8 FILLER_60_724 ();
 sg13g2_fill_2 FILLER_60_731 ();
 sg13g2_fill_2 FILLER_60_743 ();
 sg13g2_fill_1 FILLER_60_745 ();
 sg13g2_decap_8 FILLER_60_760 ();
 sg13g2_fill_1 FILLER_60_767 ();
 sg13g2_fill_1 FILLER_60_778 ();
 sg13g2_fill_2 FILLER_60_813 ();
 sg13g2_fill_1 FILLER_60_819 ();
 sg13g2_fill_2 FILLER_60_832 ();
 sg13g2_decap_8 FILLER_60_865 ();
 sg13g2_decap_4 FILLER_60_872 ();
 sg13g2_decap_8 FILLER_60_902 ();
 sg13g2_fill_2 FILLER_60_909 ();
 sg13g2_fill_1 FILLER_60_911 ();
 sg13g2_decap_4 FILLER_60_954 ();
 sg13g2_fill_1 FILLER_60_970 ();
 sg13g2_decap_4 FILLER_60_987 ();
 sg13g2_decap_8 FILLER_60_1023 ();
 sg13g2_decap_8 FILLER_60_1030 ();
 sg13g2_decap_8 FILLER_60_1037 ();
 sg13g2_decap_4 FILLER_60_1044 ();
 sg13g2_fill_1 FILLER_60_1053 ();
 sg13g2_fill_1 FILLER_60_1064 ();
 sg13g2_fill_2 FILLER_60_1070 ();
 sg13g2_fill_1 FILLER_60_1086 ();
 sg13g2_fill_2 FILLER_60_1121 ();
 sg13g2_fill_1 FILLER_60_1154 ();
 sg13g2_fill_2 FILLER_60_1159 ();
 sg13g2_fill_2 FILLER_60_1176 ();
 sg13g2_fill_2 FILLER_60_1184 ();
 sg13g2_decap_8 FILLER_60_1217 ();
 sg13g2_decap_8 FILLER_60_1224 ();
 sg13g2_decap_8 FILLER_60_1231 ();
 sg13g2_fill_1 FILLER_60_1238 ();
 sg13g2_decap_8 FILLER_60_1243 ();
 sg13g2_fill_2 FILLER_60_1253 ();
 sg13g2_fill_1 FILLER_60_1255 ();
 sg13g2_decap_8 FILLER_60_1262 ();
 sg13g2_decap_8 FILLER_60_1269 ();
 sg13g2_decap_8 FILLER_60_1276 ();
 sg13g2_decap_8 FILLER_60_1283 ();
 sg13g2_decap_8 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1297 ();
 sg13g2_decap_4 FILLER_60_1304 ();
 sg13g2_decap_4 FILLER_60_1312 ();
 sg13g2_fill_1 FILLER_60_1316 ();
 sg13g2_fill_1 FILLER_60_1322 ();
 sg13g2_fill_2 FILLER_60_1328 ();
 sg13g2_fill_1 FILLER_60_1356 ();
 sg13g2_fill_2 FILLER_60_1376 ();
 sg13g2_fill_1 FILLER_60_1382 ();
 sg13g2_fill_1 FILLER_60_1397 ();
 sg13g2_fill_1 FILLER_60_1408 ();
 sg13g2_fill_2 FILLER_60_1415 ();
 sg13g2_decap_8 FILLER_60_1427 ();
 sg13g2_decap_8 FILLER_60_1434 ();
 sg13g2_decap_8 FILLER_60_1441 ();
 sg13g2_decap_8 FILLER_60_1448 ();
 sg13g2_decap_8 FILLER_60_1455 ();
 sg13g2_fill_1 FILLER_60_1462 ();
 sg13g2_fill_1 FILLER_60_1476 ();
 sg13g2_decap_8 FILLER_60_1507 ();
 sg13g2_decap_8 FILLER_60_1514 ();
 sg13g2_fill_2 FILLER_60_1537 ();
 sg13g2_fill_2 FILLER_60_1572 ();
 sg13g2_fill_1 FILLER_60_1574 ();
 sg13g2_decap_4 FILLER_60_1579 ();
 sg13g2_decap_4 FILLER_60_1586 ();
 sg13g2_decap_4 FILLER_60_1632 ();
 sg13g2_fill_2 FILLER_60_1636 ();
 sg13g2_fill_2 FILLER_60_1651 ();
 sg13g2_fill_1 FILLER_60_1661 ();
 sg13g2_decap_8 FILLER_60_1666 ();
 sg13g2_decap_8 FILLER_60_1678 ();
 sg13g2_decap_4 FILLER_60_1685 ();
 sg13g2_fill_2 FILLER_60_1689 ();
 sg13g2_decap_8 FILLER_60_1695 ();
 sg13g2_decap_8 FILLER_60_1702 ();
 sg13g2_fill_2 FILLER_60_1748 ();
 sg13g2_decap_8 FILLER_60_1755 ();
 sg13g2_decap_8 FILLER_60_1762 ();
 sg13g2_fill_2 FILLER_60_1769 ();
 sg13g2_fill_1 FILLER_60_1771 ();
 sg13g2_decap_8 FILLER_60_1791 ();
 sg13g2_decap_8 FILLER_60_1798 ();
 sg13g2_decap_8 FILLER_60_1805 ();
 sg13g2_decap_8 FILLER_60_1815 ();
 sg13g2_decap_8 FILLER_60_1822 ();
 sg13g2_decap_8 FILLER_60_1829 ();
 sg13g2_decap_8 FILLER_60_1836 ();
 sg13g2_fill_1 FILLER_60_1843 ();
 sg13g2_decap_8 FILLER_60_1884 ();
 sg13g2_decap_8 FILLER_60_1891 ();
 sg13g2_fill_2 FILLER_60_1898 ();
 sg13g2_fill_1 FILLER_60_1900 ();
 sg13g2_fill_1 FILLER_60_1928 ();
 sg13g2_decap_8 FILLER_60_1934 ();
 sg13g2_decap_4 FILLER_60_1941 ();
 sg13g2_fill_1 FILLER_60_1945 ();
 sg13g2_decap_8 FILLER_60_1954 ();
 sg13g2_decap_4 FILLER_60_1961 ();
 sg13g2_fill_2 FILLER_60_1965 ();
 sg13g2_decap_4 FILLER_60_2029 ();
 sg13g2_fill_1 FILLER_60_2033 ();
 sg13g2_fill_1 FILLER_60_2060 ();
 sg13g2_fill_2 FILLER_60_2069 ();
 sg13g2_decap_8 FILLER_60_2134 ();
 sg13g2_decap_8 FILLER_60_2141 ();
 sg13g2_decap_4 FILLER_60_2148 ();
 sg13g2_fill_1 FILLER_60_2152 ();
 sg13g2_decap_4 FILLER_60_2158 ();
 sg13g2_decap_4 FILLER_60_2208 ();
 sg13g2_decap_8 FILLER_60_2216 ();
 sg13g2_decap_8 FILLER_60_2223 ();
 sg13g2_fill_2 FILLER_60_2230 ();
 sg13g2_decap_8 FILLER_60_2236 ();
 sg13g2_decap_8 FILLER_60_2243 ();
 sg13g2_fill_2 FILLER_60_2250 ();
 sg13g2_decap_8 FILLER_60_2337 ();
 sg13g2_decap_8 FILLER_60_2344 ();
 sg13g2_decap_8 FILLER_60_2351 ();
 sg13g2_fill_1 FILLER_60_2358 ();
 sg13g2_fill_1 FILLER_60_2371 ();
 sg13g2_decap_8 FILLER_60_2403 ();
 sg13g2_decap_8 FILLER_60_2410 ();
 sg13g2_decap_8 FILLER_60_2417 ();
 sg13g2_decap_8 FILLER_60_2424 ();
 sg13g2_decap_4 FILLER_60_2431 ();
 sg13g2_fill_2 FILLER_60_2467 ();
 sg13g2_decap_4 FILLER_60_2516 ();
 sg13g2_fill_1 FILLER_60_2520 ();
 sg13g2_decap_8 FILLER_60_2525 ();
 sg13g2_decap_8 FILLER_60_2532 ();
 sg13g2_decap_8 FILLER_60_2539 ();
 sg13g2_decap_8 FILLER_60_2546 ();
 sg13g2_decap_8 FILLER_60_2553 ();
 sg13g2_decap_8 FILLER_60_2560 ();
 sg13g2_decap_8 FILLER_60_2567 ();
 sg13g2_decap_8 FILLER_60_2574 ();
 sg13g2_decap_8 FILLER_60_2581 ();
 sg13g2_decap_8 FILLER_60_2588 ();
 sg13g2_decap_8 FILLER_60_2595 ();
 sg13g2_decap_8 FILLER_60_2602 ();
 sg13g2_decap_8 FILLER_60_2609 ();
 sg13g2_decap_8 FILLER_60_2616 ();
 sg13g2_decap_8 FILLER_60_2623 ();
 sg13g2_decap_8 FILLER_60_2630 ();
 sg13g2_decap_8 FILLER_60_2637 ();
 sg13g2_decap_8 FILLER_60_2644 ();
 sg13g2_decap_8 FILLER_60_2651 ();
 sg13g2_decap_8 FILLER_60_2658 ();
 sg13g2_decap_4 FILLER_60_2665 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_15 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_1 FILLER_61_37 ();
 sg13g2_fill_2 FILLER_61_48 ();
 sg13g2_fill_2 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_76 ();
 sg13g2_fill_2 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_83 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_113 ();
 sg13g2_fill_1 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_1 FILLER_61_137 ();
 sg13g2_fill_1 FILLER_61_143 ();
 sg13g2_fill_2 FILLER_61_148 ();
 sg13g2_fill_1 FILLER_61_150 ();
 sg13g2_fill_2 FILLER_61_161 ();
 sg13g2_fill_2 FILLER_61_183 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_decap_4 FILLER_61_198 ();
 sg13g2_fill_2 FILLER_61_207 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_fill_1 FILLER_61_220 ();
 sg13g2_decap_4 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_289 ();
 sg13g2_decap_8 FILLER_61_296 ();
 sg13g2_decap_4 FILLER_61_303 ();
 sg13g2_decap_4 FILLER_61_311 ();
 sg13g2_fill_1 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_decap_8 FILLER_61_328 ();
 sg13g2_fill_1 FILLER_61_353 ();
 sg13g2_fill_2 FILLER_61_363 ();
 sg13g2_fill_1 FILLER_61_365 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_decap_8 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_61_435 ();
 sg13g2_decap_4 FILLER_61_442 ();
 sg13g2_fill_2 FILLER_61_446 ();
 sg13g2_decap_8 FILLER_61_452 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_decap_8 FILLER_61_466 ();
 sg13g2_decap_8 FILLER_61_473 ();
 sg13g2_decap_8 FILLER_61_480 ();
 sg13g2_fill_2 FILLER_61_487 ();
 sg13g2_fill_1 FILLER_61_489 ();
 sg13g2_fill_1 FILLER_61_506 ();
 sg13g2_fill_2 FILLER_61_512 ();
 sg13g2_fill_1 FILLER_61_519 ();
 sg13g2_fill_1 FILLER_61_528 ();
 sg13g2_fill_1 FILLER_61_547 ();
 sg13g2_fill_2 FILLER_61_619 ();
 sg13g2_fill_2 FILLER_61_624 ();
 sg13g2_fill_1 FILLER_61_626 ();
 sg13g2_fill_1 FILLER_61_632 ();
 sg13g2_decap_8 FILLER_61_692 ();
 sg13g2_decap_4 FILLER_61_699 ();
 sg13g2_fill_2 FILLER_61_752 ();
 sg13g2_fill_2 FILLER_61_786 ();
 sg13g2_fill_1 FILLER_61_788 ();
 sg13g2_decap_4 FILLER_61_798 ();
 sg13g2_fill_2 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_808 ();
 sg13g2_fill_1 FILLER_61_815 ();
 sg13g2_decap_4 FILLER_61_826 ();
 sg13g2_fill_1 FILLER_61_856 ();
 sg13g2_decap_8 FILLER_61_861 ();
 sg13g2_fill_2 FILLER_61_868 ();
 sg13g2_decap_8 FILLER_61_893 ();
 sg13g2_decap_8 FILLER_61_900 ();
 sg13g2_decap_8 FILLER_61_907 ();
 sg13g2_decap_8 FILLER_61_914 ();
 sg13g2_decap_4 FILLER_61_921 ();
 sg13g2_fill_1 FILLER_61_925 ();
 sg13g2_decap_8 FILLER_61_958 ();
 sg13g2_fill_2 FILLER_61_965 ();
 sg13g2_fill_1 FILLER_61_967 ();
 sg13g2_decap_8 FILLER_61_972 ();
 sg13g2_fill_1 FILLER_61_979 ();
 sg13g2_decap_4 FILLER_61_986 ();
 sg13g2_fill_1 FILLER_61_999 ();
 sg13g2_decap_8 FILLER_61_1009 ();
 sg13g2_fill_1 FILLER_61_1016 ();
 sg13g2_fill_1 FILLER_61_1028 ();
 sg13g2_fill_2 FILLER_61_1034 ();
 sg13g2_fill_1 FILLER_61_1036 ();
 sg13g2_fill_1 FILLER_61_1047 ();
 sg13g2_fill_2 FILLER_61_1058 ();
 sg13g2_fill_1 FILLER_61_1066 ();
 sg13g2_fill_1 FILLER_61_1094 ();
 sg13g2_fill_2 FILLER_61_1101 ();
 sg13g2_fill_2 FILLER_61_1109 ();
 sg13g2_fill_2 FILLER_61_1115 ();
 sg13g2_fill_1 FILLER_61_1117 ();
 sg13g2_decap_4 FILLER_61_1124 ();
 sg13g2_fill_1 FILLER_61_1128 ();
 sg13g2_decap_8 FILLER_61_1135 ();
 sg13g2_decap_4 FILLER_61_1142 ();
 sg13g2_fill_2 FILLER_61_1146 ();
 sg13g2_fill_2 FILLER_61_1152 ();
 sg13g2_fill_2 FILLER_61_1173 ();
 sg13g2_decap_8 FILLER_61_1179 ();
 sg13g2_fill_2 FILLER_61_1186 ();
 sg13g2_fill_1 FILLER_61_1188 ();
 sg13g2_fill_1 FILLER_61_1194 ();
 sg13g2_fill_1 FILLER_61_1201 ();
 sg13g2_fill_1 FILLER_61_1207 ();
 sg13g2_fill_1 FILLER_61_1249 ();
 sg13g2_decap_8 FILLER_61_1291 ();
 sg13g2_fill_2 FILLER_61_1298 ();
 sg13g2_fill_1 FILLER_61_1300 ();
 sg13g2_fill_1 FILLER_61_1354 ();
 sg13g2_fill_1 FILLER_61_1360 ();
 sg13g2_fill_1 FILLER_61_1374 ();
 sg13g2_fill_1 FILLER_61_1422 ();
 sg13g2_fill_2 FILLER_61_1458 ();
 sg13g2_decap_4 FILLER_61_1477 ();
 sg13g2_fill_1 FILLER_61_1481 ();
 sg13g2_decap_4 FILLER_61_1486 ();
 sg13g2_decap_8 FILLER_61_1500 ();
 sg13g2_decap_8 FILLER_61_1507 ();
 sg13g2_decap_8 FILLER_61_1514 ();
 sg13g2_fill_2 FILLER_61_1521 ();
 sg13g2_fill_1 FILLER_61_1523 ();
 sg13g2_fill_1 FILLER_61_1528 ();
 sg13g2_fill_1 FILLER_61_1535 ();
 sg13g2_fill_2 FILLER_61_1562 ();
 sg13g2_fill_2 FILLER_61_1568 ();
 sg13g2_fill_1 FILLER_61_1634 ();
 sg13g2_fill_1 FILLER_61_1666 ();
 sg13g2_fill_1 FILLER_61_1672 ();
 sg13g2_decap_8 FILLER_61_1688 ();
 sg13g2_fill_1 FILLER_61_1695 ();
 sg13g2_decap_8 FILLER_61_1722 ();
 sg13g2_decap_8 FILLER_61_1729 ();
 sg13g2_decap_8 FILLER_61_1736 ();
 sg13g2_decap_8 FILLER_61_1743 ();
 sg13g2_decap_8 FILLER_61_1750 ();
 sg13g2_fill_2 FILLER_61_1757 ();
 sg13g2_fill_1 FILLER_61_1759 ();
 sg13g2_decap_8 FILLER_61_1765 ();
 sg13g2_decap_8 FILLER_61_1772 ();
 sg13g2_decap_8 FILLER_61_1779 ();
 sg13g2_decap_4 FILLER_61_1791 ();
 sg13g2_fill_2 FILLER_61_1795 ();
 sg13g2_decap_8 FILLER_61_1807 ();
 sg13g2_decap_8 FILLER_61_1814 ();
 sg13g2_fill_2 FILLER_61_1821 ();
 sg13g2_fill_1 FILLER_61_1823 ();
 sg13g2_fill_1 FILLER_61_1838 ();
 sg13g2_decap_4 FILLER_61_1884 ();
 sg13g2_fill_1 FILLER_61_1888 ();
 sg13g2_fill_2 FILLER_61_1894 ();
 sg13g2_decap_4 FILLER_61_1928 ();
 sg13g2_fill_1 FILLER_61_1932 ();
 sg13g2_fill_1 FILLER_61_1938 ();
 sg13g2_decap_8 FILLER_61_1943 ();
 sg13g2_decap_8 FILLER_61_1950 ();
 sg13g2_fill_1 FILLER_61_1957 ();
 sg13g2_decap_8 FILLER_61_1962 ();
 sg13g2_decap_4 FILLER_61_1969 ();
 sg13g2_fill_1 FILLER_61_1973 ();
 sg13g2_fill_1 FILLER_61_1989 ();
 sg13g2_decap_4 FILLER_61_1999 ();
 sg13g2_fill_1 FILLER_61_2003 ();
 sg13g2_decap_8 FILLER_61_2030 ();
 sg13g2_decap_4 FILLER_61_2037 ();
 sg13g2_fill_1 FILLER_61_2076 ();
 sg13g2_fill_1 FILLER_61_2101 ();
 sg13g2_decap_8 FILLER_61_2125 ();
 sg13g2_fill_2 FILLER_61_2132 ();
 sg13g2_fill_2 FILLER_61_2139 ();
 sg13g2_decap_4 FILLER_61_2145 ();
 sg13g2_fill_2 FILLER_61_2149 ();
 sg13g2_decap_4 FILLER_61_2182 ();
 sg13g2_decap_8 FILLER_61_2217 ();
 sg13g2_decap_8 FILLER_61_2224 ();
 sg13g2_decap_8 FILLER_61_2231 ();
 sg13g2_decap_8 FILLER_61_2238 ();
 sg13g2_fill_1 FILLER_61_2245 ();
 sg13g2_fill_2 FILLER_61_2250 ();
 sg13g2_fill_1 FILLER_61_2252 ();
 sg13g2_fill_2 FILLER_61_2262 ();
 sg13g2_fill_2 FILLER_61_2290 ();
 sg13g2_decap_4 FILLER_61_2328 ();
 sg13g2_fill_1 FILLER_61_2332 ();
 sg13g2_decap_4 FILLER_61_2363 ();
 sg13g2_fill_1 FILLER_61_2367 ();
 sg13g2_decap_4 FILLER_61_2371 ();
 sg13g2_fill_1 FILLER_61_2384 ();
 sg13g2_fill_1 FILLER_61_2411 ();
 sg13g2_decap_8 FILLER_61_2416 ();
 sg13g2_decap_8 FILLER_61_2423 ();
 sg13g2_fill_1 FILLER_61_2430 ();
 sg13g2_fill_1 FILLER_61_2461 ();
 sg13g2_fill_1 FILLER_61_2468 ();
 sg13g2_decap_8 FILLER_61_2498 ();
 sg13g2_decap_4 FILLER_61_2505 ();
 sg13g2_fill_1 FILLER_61_2509 ();
 sg13g2_decap_8 FILLER_61_2540 ();
 sg13g2_decap_8 FILLER_61_2547 ();
 sg13g2_decap_8 FILLER_61_2554 ();
 sg13g2_decap_8 FILLER_61_2561 ();
 sg13g2_decap_8 FILLER_61_2568 ();
 sg13g2_decap_8 FILLER_61_2575 ();
 sg13g2_decap_8 FILLER_61_2582 ();
 sg13g2_decap_8 FILLER_61_2589 ();
 sg13g2_decap_8 FILLER_61_2596 ();
 sg13g2_decap_8 FILLER_61_2603 ();
 sg13g2_decap_8 FILLER_61_2610 ();
 sg13g2_decap_8 FILLER_61_2617 ();
 sg13g2_decap_8 FILLER_61_2624 ();
 sg13g2_decap_8 FILLER_61_2631 ();
 sg13g2_decap_8 FILLER_61_2638 ();
 sg13g2_decap_8 FILLER_61_2645 ();
 sg13g2_decap_8 FILLER_61_2652 ();
 sg13g2_decap_8 FILLER_61_2659 ();
 sg13g2_decap_4 FILLER_61_2666 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_4 ();
 sg13g2_fill_2 FILLER_62_10 ();
 sg13g2_fill_1 FILLER_62_25 ();
 sg13g2_fill_1 FILLER_62_49 ();
 sg13g2_fill_2 FILLER_62_55 ();
 sg13g2_fill_1 FILLER_62_85 ();
 sg13g2_fill_1 FILLER_62_99 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_fill_2 FILLER_62_145 ();
 sg13g2_fill_2 FILLER_62_151 ();
 sg13g2_fill_2 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_202 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_decap_8 FILLER_62_215 ();
 sg13g2_decap_4 FILLER_62_222 ();
 sg13g2_fill_2 FILLER_62_226 ();
 sg13g2_decap_4 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_248 ();
 sg13g2_decap_4 FILLER_62_270 ();
 sg13g2_fill_2 FILLER_62_274 ();
 sg13g2_decap_8 FILLER_62_306 ();
 sg13g2_decap_8 FILLER_62_313 ();
 sg13g2_decap_8 FILLER_62_320 ();
 sg13g2_decap_4 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_331 ();
 sg13g2_decap_4 FILLER_62_358 ();
 sg13g2_fill_1 FILLER_62_362 ();
 sg13g2_fill_2 FILLER_62_377 ();
 sg13g2_fill_2 FILLER_62_393 ();
 sg13g2_fill_1 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_431 ();
 sg13g2_decap_8 FILLER_62_473 ();
 sg13g2_decap_4 FILLER_62_480 ();
 sg13g2_fill_1 FILLER_62_484 ();
 sg13g2_fill_2 FILLER_62_493 ();
 sg13g2_fill_1 FILLER_62_495 ();
 sg13g2_fill_1 FILLER_62_519 ();
 sg13g2_decap_8 FILLER_62_525 ();
 sg13g2_decap_8 FILLER_62_532 ();
 sg13g2_fill_2 FILLER_62_539 ();
 sg13g2_fill_1 FILLER_62_555 ();
 sg13g2_decap_4 FILLER_62_579 ();
 sg13g2_fill_1 FILLER_62_592 ();
 sg13g2_decap_8 FILLER_62_620 ();
 sg13g2_decap_8 FILLER_62_627 ();
 sg13g2_decap_8 FILLER_62_634 ();
 sg13g2_fill_1 FILLER_62_641 ();
 sg13g2_fill_1 FILLER_62_659 ();
 sg13g2_decap_8 FILLER_62_689 ();
 sg13g2_decap_8 FILLER_62_696 ();
 sg13g2_decap_4 FILLER_62_703 ();
 sg13g2_fill_2 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_726 ();
 sg13g2_decap_4 FILLER_62_733 ();
 sg13g2_fill_1 FILLER_62_737 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_fill_2 FILLER_62_749 ();
 sg13g2_fill_1 FILLER_62_751 ();
 sg13g2_fill_2 FILLER_62_757 ();
 sg13g2_fill_1 FILLER_62_759 ();
 sg13g2_decap_4 FILLER_62_764 ();
 sg13g2_fill_2 FILLER_62_773 ();
 sg13g2_decap_4 FILLER_62_780 ();
 sg13g2_fill_2 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_decap_4 FILLER_62_802 ();
 sg13g2_fill_1 FILLER_62_811 ();
 sg13g2_fill_2 FILLER_62_851 ();
 sg13g2_decap_8 FILLER_62_857 ();
 sg13g2_fill_2 FILLER_62_864 ();
 sg13g2_fill_1 FILLER_62_866 ();
 sg13g2_decap_8 FILLER_62_871 ();
 sg13g2_decap_8 FILLER_62_878 ();
 sg13g2_fill_2 FILLER_62_885 ();
 sg13g2_decap_8 FILLER_62_891 ();
 sg13g2_decap_4 FILLER_62_898 ();
 sg13g2_fill_2 FILLER_62_902 ();
 sg13g2_decap_4 FILLER_62_987 ();
 sg13g2_fill_2 FILLER_62_1017 ();
 sg13g2_fill_1 FILLER_62_1019 ();
 sg13g2_fill_1 FILLER_62_1088 ();
 sg13g2_fill_1 FILLER_62_1099 ();
 sg13g2_decap_4 FILLER_62_1104 ();
 sg13g2_fill_2 FILLER_62_1131 ();
 sg13g2_fill_1 FILLER_62_1133 ();
 sg13g2_fill_2 FILLER_62_1140 ();
 sg13g2_fill_2 FILLER_62_1147 ();
 sg13g2_fill_1 FILLER_62_1154 ();
 sg13g2_fill_2 FILLER_62_1159 ();
 sg13g2_decap_8 FILLER_62_1179 ();
 sg13g2_decap_4 FILLER_62_1186 ();
 sg13g2_fill_1 FILLER_62_1190 ();
 sg13g2_decap_4 FILLER_62_1195 ();
 sg13g2_decap_8 FILLER_62_1205 ();
 sg13g2_decap_8 FILLER_62_1212 ();
 sg13g2_decap_8 FILLER_62_1219 ();
 sg13g2_decap_8 FILLER_62_1226 ();
 sg13g2_decap_8 FILLER_62_1233 ();
 sg13g2_decap_4 FILLER_62_1240 ();
 sg13g2_fill_2 FILLER_62_1244 ();
 sg13g2_fill_1 FILLER_62_1251 ();
 sg13g2_fill_1 FILLER_62_1302 ();
 sg13g2_decap_8 FILLER_62_1307 ();
 sg13g2_fill_1 FILLER_62_1314 ();
 sg13g2_fill_1 FILLER_62_1336 ();
 sg13g2_decap_8 FILLER_62_1401 ();
 sg13g2_decap_8 FILLER_62_1434 ();
 sg13g2_fill_2 FILLER_62_1441 ();
 sg13g2_fill_1 FILLER_62_1443 ();
 sg13g2_decap_8 FILLER_62_1448 ();
 sg13g2_fill_2 FILLER_62_1455 ();
 sg13g2_decap_8 FILLER_62_1465 ();
 sg13g2_fill_2 FILLER_62_1472 ();
 sg13g2_decap_8 FILLER_62_1508 ();
 sg13g2_decap_8 FILLER_62_1515 ();
 sg13g2_fill_2 FILLER_62_1522 ();
 sg13g2_fill_1 FILLER_62_1524 ();
 sg13g2_fill_2 FILLER_62_1534 ();
 sg13g2_fill_2 FILLER_62_1548 ();
 sg13g2_fill_2 FILLER_62_1569 ();
 sg13g2_fill_1 FILLER_62_1585 ();
 sg13g2_decap_4 FILLER_62_1592 ();
 sg13g2_fill_1 FILLER_62_1611 ();
 sg13g2_decap_8 FILLER_62_1645 ();
 sg13g2_fill_2 FILLER_62_1652 ();
 sg13g2_fill_1 FILLER_62_1654 ();
 sg13g2_fill_2 FILLER_62_1667 ();
 sg13g2_fill_1 FILLER_62_1669 ();
 sg13g2_fill_1 FILLER_62_1681 ();
 sg13g2_fill_2 FILLER_62_1714 ();
 sg13g2_fill_1 FILLER_62_1716 ();
 sg13g2_fill_2 FILLER_62_1743 ();
 sg13g2_fill_1 FILLER_62_1745 ();
 sg13g2_fill_2 FILLER_62_1808 ();
 sg13g2_decap_8 FILLER_62_1857 ();
 sg13g2_fill_1 FILLER_62_1864 ();
 sg13g2_decap_8 FILLER_62_1874 ();
 sg13g2_fill_2 FILLER_62_1881 ();
 sg13g2_decap_8 FILLER_62_1888 ();
 sg13g2_decap_8 FILLER_62_1895 ();
 sg13g2_decap_8 FILLER_62_1902 ();
 sg13g2_fill_1 FILLER_62_1909 ();
 sg13g2_decap_4 FILLER_62_1914 ();
 sg13g2_fill_1 FILLER_62_1918 ();
 sg13g2_decap_4 FILLER_62_1945 ();
 sg13g2_fill_2 FILLER_62_1949 ();
 sg13g2_decap_4 FILLER_62_1960 ();
 sg13g2_fill_2 FILLER_62_1993 ();
 sg13g2_fill_1 FILLER_62_1995 ();
 sg13g2_decap_8 FILLER_62_2001 ();
 sg13g2_fill_1 FILLER_62_2013 ();
 sg13g2_decap_8 FILLER_62_2018 ();
 sg13g2_decap_8 FILLER_62_2025 ();
 sg13g2_decap_4 FILLER_62_2032 ();
 sg13g2_fill_2 FILLER_62_2036 ();
 sg13g2_fill_1 FILLER_62_2051 ();
 sg13g2_fill_1 FILLER_62_2106 ();
 sg13g2_fill_2 FILLER_62_2115 ();
 sg13g2_fill_2 FILLER_62_2123 ();
 sg13g2_fill_2 FILLER_62_2151 ();
 sg13g2_decap_8 FILLER_62_2162 ();
 sg13g2_decap_8 FILLER_62_2169 ();
 sg13g2_fill_1 FILLER_62_2176 ();
 sg13g2_fill_2 FILLER_62_2218 ();
 sg13g2_decap_4 FILLER_62_2230 ();
 sg13g2_fill_2 FILLER_62_2276 ();
 sg13g2_fill_1 FILLER_62_2278 ();
 sg13g2_decap_4 FILLER_62_2308 ();
 sg13g2_decap_8 FILLER_62_2316 ();
 sg13g2_decap_8 FILLER_62_2372 ();
 sg13g2_decap_8 FILLER_62_2388 ();
 sg13g2_decap_8 FILLER_62_2395 ();
 sg13g2_decap_4 FILLER_62_2402 ();
 sg13g2_fill_2 FILLER_62_2406 ();
 sg13g2_fill_1 FILLER_62_2412 ();
 sg13g2_fill_2 FILLER_62_2439 ();
 sg13g2_fill_2 FILLER_62_2445 ();
 sg13g2_fill_2 FILLER_62_2451 ();
 sg13g2_decap_8 FILLER_62_2457 ();
 sg13g2_decap_4 FILLER_62_2464 ();
 sg13g2_fill_1 FILLER_62_2468 ();
 sg13g2_decap_8 FILLER_62_2472 ();
 sg13g2_decap_4 FILLER_62_2483 ();
 sg13g2_decap_8 FILLER_62_2491 ();
 sg13g2_decap_8 FILLER_62_2498 ();
 sg13g2_fill_2 FILLER_62_2505 ();
 sg13g2_decap_8 FILLER_62_2549 ();
 sg13g2_decap_8 FILLER_62_2556 ();
 sg13g2_decap_8 FILLER_62_2563 ();
 sg13g2_decap_8 FILLER_62_2570 ();
 sg13g2_decap_8 FILLER_62_2577 ();
 sg13g2_decap_8 FILLER_62_2584 ();
 sg13g2_decap_8 FILLER_62_2591 ();
 sg13g2_decap_8 FILLER_62_2598 ();
 sg13g2_decap_8 FILLER_62_2605 ();
 sg13g2_decap_8 FILLER_62_2612 ();
 sg13g2_decap_8 FILLER_62_2619 ();
 sg13g2_decap_8 FILLER_62_2626 ();
 sg13g2_decap_8 FILLER_62_2633 ();
 sg13g2_decap_8 FILLER_62_2640 ();
 sg13g2_decap_8 FILLER_62_2647 ();
 sg13g2_decap_8 FILLER_62_2654 ();
 sg13g2_decap_8 FILLER_62_2661 ();
 sg13g2_fill_2 FILLER_62_2668 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_11 ();
 sg13g2_fill_1 FILLER_63_31 ();
 sg13g2_fill_2 FILLER_63_46 ();
 sg13g2_fill_1 FILLER_63_48 ();
 sg13g2_fill_2 FILLER_63_114 ();
 sg13g2_fill_2 FILLER_63_135 ();
 sg13g2_fill_2 FILLER_63_142 ();
 sg13g2_fill_2 FILLER_63_149 ();
 sg13g2_fill_1 FILLER_63_157 ();
 sg13g2_fill_1 FILLER_63_179 ();
 sg13g2_fill_1 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_203 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_221 ();
 sg13g2_decap_8 FILLER_63_228 ();
 sg13g2_decap_8 FILLER_63_235 ();
 sg13g2_decap_8 FILLER_63_242 ();
 sg13g2_fill_2 FILLER_63_249 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_fill_2 FILLER_63_257 ();
 sg13g2_fill_2 FILLER_63_264 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_fill_2 FILLER_63_275 ();
 sg13g2_fill_1 FILLER_63_277 ();
 sg13g2_fill_2 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_285 ();
 sg13g2_decap_8 FILLER_63_303 ();
 sg13g2_decap_8 FILLER_63_310 ();
 sg13g2_decap_4 FILLER_63_317 ();
 sg13g2_fill_2 FILLER_63_321 ();
 sg13g2_fill_1 FILLER_63_352 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_1 FILLER_63_368 ();
 sg13g2_fill_1 FILLER_63_381 ();
 sg13g2_fill_2 FILLER_63_391 ();
 sg13g2_fill_2 FILLER_63_426 ();
 sg13g2_decap_4 FILLER_63_437 ();
 sg13g2_fill_1 FILLER_63_441 ();
 sg13g2_fill_1 FILLER_63_451 ();
 sg13g2_decap_8 FILLER_63_457 ();
 sg13g2_decap_8 FILLER_63_464 ();
 sg13g2_decap_8 FILLER_63_471 ();
 sg13g2_decap_8 FILLER_63_478 ();
 sg13g2_fill_2 FILLER_63_485 ();
 sg13g2_fill_1 FILLER_63_494 ();
 sg13g2_fill_1 FILLER_63_500 ();
 sg13g2_fill_2 FILLER_63_504 ();
 sg13g2_fill_2 FILLER_63_516 ();
 sg13g2_decap_8 FILLER_63_523 ();
 sg13g2_fill_2 FILLER_63_530 ();
 sg13g2_decap_4 FILLER_63_540 ();
 sg13g2_fill_2 FILLER_63_551 ();
 sg13g2_fill_1 FILLER_63_576 ();
 sg13g2_fill_2 FILLER_63_581 ();
 sg13g2_fill_2 FILLER_63_588 ();
 sg13g2_fill_2 FILLER_63_595 ();
 sg13g2_fill_1 FILLER_63_611 ();
 sg13g2_fill_1 FILLER_63_617 ();
 sg13g2_fill_1 FILLER_63_623 ();
 sg13g2_fill_1 FILLER_63_629 ();
 sg13g2_decap_8 FILLER_63_634 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_fill_2 FILLER_63_666 ();
 sg13g2_decap_8 FILLER_63_687 ();
 sg13g2_decap_8 FILLER_63_694 ();
 sg13g2_fill_1 FILLER_63_701 ();
 sg13g2_fill_1 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_4 FILLER_63_746 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_4 FILLER_63_770 ();
 sg13g2_fill_2 FILLER_63_774 ();
 sg13g2_decap_4 FILLER_63_806 ();
 sg13g2_fill_2 FILLER_63_810 ();
 sg13g2_decap_8 FILLER_63_842 ();
 sg13g2_fill_1 FILLER_63_849 ();
 sg13g2_decap_4 FILLER_63_915 ();
 sg13g2_fill_2 FILLER_63_923 ();
 sg13g2_fill_1 FILLER_63_925 ();
 sg13g2_fill_2 FILLER_63_964 ();
 sg13g2_decap_8 FILLER_63_972 ();
 sg13g2_decap_8 FILLER_63_979 ();
 sg13g2_fill_2 FILLER_63_986 ();
 sg13g2_fill_1 FILLER_63_988 ();
 sg13g2_fill_1 FILLER_63_998 ();
 sg13g2_decap_8 FILLER_63_1003 ();
 sg13g2_decap_8 FILLER_63_1010 ();
 sg13g2_decap_4 FILLER_63_1017 ();
 sg13g2_fill_1 FILLER_63_1021 ();
 sg13g2_decap_8 FILLER_63_1028 ();
 sg13g2_decap_8 FILLER_63_1035 ();
 sg13g2_fill_2 FILLER_63_1042 ();
 sg13g2_fill_1 FILLER_63_1044 ();
 sg13g2_fill_1 FILLER_63_1086 ();
 sg13g2_decap_8 FILLER_63_1133 ();
 sg13g2_decap_4 FILLER_63_1140 ();
 sg13g2_fill_1 FILLER_63_1180 ();
 sg13g2_decap_4 FILLER_63_1217 ();
 sg13g2_fill_2 FILLER_63_1221 ();
 sg13g2_decap_4 FILLER_63_1227 ();
 sg13g2_fill_1 FILLER_63_1231 ();
 sg13g2_fill_2 FILLER_63_1238 ();
 sg13g2_decap_4 FILLER_63_1251 ();
 sg13g2_decap_4 FILLER_63_1277 ();
 sg13g2_fill_2 FILLER_63_1281 ();
 sg13g2_decap_8 FILLER_63_1320 ();
 sg13g2_fill_2 FILLER_63_1327 ();
 sg13g2_fill_2 FILLER_63_1362 ();
 sg13g2_decap_4 FILLER_63_1369 ();
 sg13g2_fill_2 FILLER_63_1379 ();
 sg13g2_fill_1 FILLER_63_1384 ();
 sg13g2_decap_8 FILLER_63_1391 ();
 sg13g2_decap_8 FILLER_63_1398 ();
 sg13g2_decap_8 FILLER_63_1405 ();
 sg13g2_decap_8 FILLER_63_1412 ();
 sg13g2_decap_8 FILLER_63_1419 ();
 sg13g2_decap_8 FILLER_63_1426 ();
 sg13g2_fill_1 FILLER_63_1433 ();
 sg13g2_decap_4 FILLER_63_1460 ();
 sg13g2_fill_1 FILLER_63_1490 ();
 sg13g2_fill_1 FILLER_63_1497 ();
 sg13g2_fill_1 FILLER_63_1504 ();
 sg13g2_decap_4 FILLER_63_1509 ();
 sg13g2_fill_1 FILLER_63_1513 ();
 sg13g2_fill_2 FILLER_63_1553 ();
 sg13g2_decap_8 FILLER_63_1569 ();
 sg13g2_decap_4 FILLER_63_1576 ();
 sg13g2_fill_2 FILLER_63_1580 ();
 sg13g2_decap_4 FILLER_63_1588 ();
 sg13g2_fill_1 FILLER_63_1610 ();
 sg13g2_decap_4 FILLER_63_1640 ();
 sg13g2_fill_2 FILLER_63_1644 ();
 sg13g2_decap_4 FILLER_63_1669 ();
 sg13g2_fill_2 FILLER_63_1712 ();
 sg13g2_fill_1 FILLER_63_1714 ();
 sg13g2_decap_8 FILLER_63_1761 ();
 sg13g2_fill_1 FILLER_63_1768 ();
 sg13g2_fill_1 FILLER_63_1801 ();
 sg13g2_fill_1 FILLER_63_1831 ();
 sg13g2_fill_2 FILLER_63_1840 ();
 sg13g2_fill_2 FILLER_63_1870 ();
 sg13g2_fill_1 FILLER_63_1872 ();
 sg13g2_fill_2 FILLER_63_1899 ();
 sg13g2_fill_1 FILLER_63_1901 ();
 sg13g2_decap_4 FILLER_63_1906 ();
 sg13g2_fill_1 FILLER_63_1910 ();
 sg13g2_decap_4 FILLER_63_1917 ();
 sg13g2_fill_1 FILLER_63_1921 ();
 sg13g2_fill_2 FILLER_63_1927 ();
 sg13g2_fill_1 FILLER_63_1929 ();
 sg13g2_decap_8 FILLER_63_1956 ();
 sg13g2_decap_4 FILLER_63_1963 ();
 sg13g2_fill_2 FILLER_63_1967 ();
 sg13g2_decap_8 FILLER_63_2008 ();
 sg13g2_decap_8 FILLER_63_2015 ();
 sg13g2_decap_8 FILLER_63_2022 ();
 sg13g2_decap_8 FILLER_63_2029 ();
 sg13g2_fill_1 FILLER_63_2036 ();
 sg13g2_decap_8 FILLER_63_2075 ();
 sg13g2_fill_1 FILLER_63_2082 ();
 sg13g2_decap_8 FILLER_63_2086 ();
 sg13g2_decap_4 FILLER_63_2093 ();
 sg13g2_fill_2 FILLER_63_2097 ();
 sg13g2_fill_2 FILLER_63_2139 ();
 sg13g2_fill_2 FILLER_63_2147 ();
 sg13g2_fill_1 FILLER_63_2149 ();
 sg13g2_decap_4 FILLER_63_2182 ();
 sg13g2_fill_2 FILLER_63_2239 ();
 sg13g2_fill_1 FILLER_63_2265 ();
 sg13g2_decap_8 FILLER_63_2297 ();
 sg13g2_fill_1 FILLER_63_2304 ();
 sg13g2_fill_1 FILLER_63_2309 ();
 sg13g2_fill_1 FILLER_63_2319 ();
 sg13g2_fill_1 FILLER_63_2355 ();
 sg13g2_decap_8 FILLER_63_2362 ();
 sg13g2_decap_8 FILLER_63_2369 ();
 sg13g2_fill_1 FILLER_63_2376 ();
 sg13g2_fill_2 FILLER_63_2406 ();
 sg13g2_decap_8 FILLER_63_2448 ();
 sg13g2_decap_8 FILLER_63_2455 ();
 sg13g2_decap_8 FILLER_63_2462 ();
 sg13g2_fill_1 FILLER_63_2469 ();
 sg13g2_decap_4 FILLER_63_2476 ();
 sg13g2_fill_2 FILLER_63_2480 ();
 sg13g2_fill_2 FILLER_63_2512 ();
 sg13g2_fill_1 FILLER_63_2514 ();
 sg13g2_decap_8 FILLER_63_2549 ();
 sg13g2_decap_8 FILLER_63_2556 ();
 sg13g2_decap_8 FILLER_63_2563 ();
 sg13g2_decap_8 FILLER_63_2570 ();
 sg13g2_decap_8 FILLER_63_2577 ();
 sg13g2_decap_8 FILLER_63_2584 ();
 sg13g2_decap_8 FILLER_63_2591 ();
 sg13g2_decap_8 FILLER_63_2598 ();
 sg13g2_decap_8 FILLER_63_2605 ();
 sg13g2_decap_8 FILLER_63_2612 ();
 sg13g2_decap_8 FILLER_63_2619 ();
 sg13g2_decap_8 FILLER_63_2626 ();
 sg13g2_decap_8 FILLER_63_2633 ();
 sg13g2_decap_8 FILLER_63_2640 ();
 sg13g2_decap_8 FILLER_63_2647 ();
 sg13g2_decap_8 FILLER_63_2654 ();
 sg13g2_decap_8 FILLER_63_2661 ();
 sg13g2_fill_2 FILLER_63_2668 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_22 ();
 sg13g2_fill_1 FILLER_64_43 ();
 sg13g2_fill_2 FILLER_64_54 ();
 sg13g2_fill_1 FILLER_64_56 ();
 sg13g2_fill_1 FILLER_64_62 ();
 sg13g2_fill_2 FILLER_64_67 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_82 ();
 sg13g2_fill_2 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_104 ();
 sg13g2_fill_1 FILLER_64_109 ();
 sg13g2_decap_4 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_131 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_fill_1 FILLER_64_175 ();
 sg13g2_fill_2 FILLER_64_180 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_decap_4 FILLER_64_201 ();
 sg13g2_fill_1 FILLER_64_205 ();
 sg13g2_fill_1 FILLER_64_214 ();
 sg13g2_fill_2 FILLER_64_220 ();
 sg13g2_fill_2 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_240 ();
 sg13g2_decap_4 FILLER_64_258 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_269 ();
 sg13g2_fill_2 FILLER_64_286 ();
 sg13g2_decap_8 FILLER_64_296 ();
 sg13g2_decap_8 FILLER_64_303 ();
 sg13g2_decap_8 FILLER_64_310 ();
 sg13g2_decap_8 FILLER_64_317 ();
 sg13g2_decap_8 FILLER_64_324 ();
 sg13g2_decap_8 FILLER_64_331 ();
 sg13g2_decap_4 FILLER_64_338 ();
 sg13g2_fill_2 FILLER_64_367 ();
 sg13g2_fill_1 FILLER_64_369 ();
 sg13g2_fill_1 FILLER_64_375 ();
 sg13g2_fill_1 FILLER_64_381 ();
 sg13g2_fill_1 FILLER_64_392 ();
 sg13g2_fill_2 FILLER_64_413 ();
 sg13g2_decap_8 FILLER_64_432 ();
 sg13g2_decap_8 FILLER_64_439 ();
 sg13g2_decap_8 FILLER_64_446 ();
 sg13g2_decap_8 FILLER_64_453 ();
 sg13g2_fill_2 FILLER_64_460 ();
 sg13g2_fill_1 FILLER_64_462 ();
 sg13g2_decap_8 FILLER_64_468 ();
 sg13g2_fill_2 FILLER_64_480 ();
 sg13g2_decap_8 FILLER_64_500 ();
 sg13g2_decap_8 FILLER_64_507 ();
 sg13g2_decap_8 FILLER_64_514 ();
 sg13g2_decap_8 FILLER_64_521 ();
 sg13g2_fill_1 FILLER_64_528 ();
 sg13g2_decap_4 FILLER_64_533 ();
 sg13g2_decap_8 FILLER_64_541 ();
 sg13g2_decap_8 FILLER_64_548 ();
 sg13g2_decap_8 FILLER_64_555 ();
 sg13g2_decap_8 FILLER_64_583 ();
 sg13g2_decap_8 FILLER_64_590 ();
 sg13g2_decap_8 FILLER_64_597 ();
 sg13g2_decap_4 FILLER_64_604 ();
 sg13g2_fill_1 FILLER_64_608 ();
 sg13g2_decap_4 FILLER_64_613 ();
 sg13g2_decap_8 FILLER_64_626 ();
 sg13g2_fill_1 FILLER_64_633 ();
 sg13g2_decap_4 FILLER_64_731 ();
 sg13g2_fill_2 FILLER_64_735 ();
 sg13g2_fill_2 FILLER_64_811 ();
 sg13g2_decap_8 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_64_868 ();
 sg13g2_decap_8 FILLER_64_875 ();
 sg13g2_decap_4 FILLER_64_882 ();
 sg13g2_fill_2 FILLER_64_926 ();
 sg13g2_decap_4 FILLER_64_932 ();
 sg13g2_fill_2 FILLER_64_936 ();
 sg13g2_decap_8 FILLER_64_944 ();
 sg13g2_fill_2 FILLER_64_951 ();
 sg13g2_fill_1 FILLER_64_953 ();
 sg13g2_fill_2 FILLER_64_964 ();
 sg13g2_fill_2 FILLER_64_970 ();
 sg13g2_fill_1 FILLER_64_981 ();
 sg13g2_fill_2 FILLER_64_995 ();
 sg13g2_fill_1 FILLER_64_997 ();
 sg13g2_decap_8 FILLER_64_1029 ();
 sg13g2_decap_4 FILLER_64_1036 ();
 sg13g2_fill_1 FILLER_64_1040 ();
 sg13g2_fill_1 FILLER_64_1068 ();
 sg13g2_fill_2 FILLER_64_1072 ();
 sg13g2_fill_1 FILLER_64_1083 ();
 sg13g2_fill_2 FILLER_64_1087 ();
 sg13g2_fill_2 FILLER_64_1100 ();
 sg13g2_decap_8 FILLER_64_1106 ();
 sg13g2_fill_1 FILLER_64_1113 ();
 sg13g2_fill_1 FILLER_64_1118 ();
 sg13g2_decap_8 FILLER_64_1123 ();
 sg13g2_fill_2 FILLER_64_1130 ();
 sg13g2_decap_4 FILLER_64_1136 ();
 sg13g2_decap_8 FILLER_64_1144 ();
 sg13g2_decap_8 FILLER_64_1151 ();
 sg13g2_fill_1 FILLER_64_1158 ();
 sg13g2_fill_2 FILLER_64_1196 ();
 sg13g2_fill_1 FILLER_64_1198 ();
 sg13g2_fill_1 FILLER_64_1227 ();
 sg13g2_fill_2 FILLER_64_1257 ();
 sg13g2_fill_1 FILLER_64_1259 ();
 sg13g2_decap_8 FILLER_64_1265 ();
 sg13g2_decap_8 FILLER_64_1306 ();
 sg13g2_decap_8 FILLER_64_1313 ();
 sg13g2_decap_4 FILLER_64_1320 ();
 sg13g2_fill_2 FILLER_64_1324 ();
 sg13g2_fill_2 FILLER_64_1355 ();
 sg13g2_decap_4 FILLER_64_1361 ();
 sg13g2_fill_2 FILLER_64_1365 ();
 sg13g2_fill_1 FILLER_64_1377 ();
 sg13g2_fill_1 FILLER_64_1387 ();
 sg13g2_fill_2 FILLER_64_1394 ();
 sg13g2_decap_4 FILLER_64_1402 ();
 sg13g2_fill_2 FILLER_64_1411 ();
 sg13g2_fill_1 FILLER_64_1413 ();
 sg13g2_decap_8 FILLER_64_1422 ();
 sg13g2_decap_8 FILLER_64_1429 ();
 sg13g2_decap_4 FILLER_64_1442 ();
 sg13g2_decap_4 FILLER_64_1466 ();
 sg13g2_fill_1 FILLER_64_1470 ();
 sg13g2_fill_2 FILLER_64_1478 ();
 sg13g2_fill_1 FILLER_64_1480 ();
 sg13g2_fill_1 FILLER_64_1524 ();
 sg13g2_fill_1 FILLER_64_1541 ();
 sg13g2_fill_2 FILLER_64_1568 ();
 sg13g2_decap_4 FILLER_64_1575 ();
 sg13g2_fill_1 FILLER_64_1591 ();
 sg13g2_decap_4 FILLER_64_1598 ();
 sg13g2_fill_1 FILLER_64_1602 ();
 sg13g2_fill_2 FILLER_64_1625 ();
 sg13g2_decap_4 FILLER_64_1694 ();
 sg13g2_fill_1 FILLER_64_1698 ();
 sg13g2_fill_2 FILLER_64_1707 ();
 sg13g2_decap_8 FILLER_64_1723 ();
 sg13g2_fill_2 FILLER_64_1730 ();
 sg13g2_fill_1 FILLER_64_1732 ();
 sg13g2_decap_4 FILLER_64_1743 ();
 sg13g2_decap_4 FILLER_64_1823 ();
 sg13g2_fill_1 FILLER_64_1827 ();
 sg13g2_decap_4 FILLER_64_1838 ();
 sg13g2_fill_1 FILLER_64_1852 ();
 sg13g2_fill_2 FILLER_64_1859 ();
 sg13g2_decap_4 FILLER_64_1887 ();
 sg13g2_fill_1 FILLER_64_1896 ();
 sg13g2_fill_2 FILLER_64_1923 ();
 sg13g2_fill_1 FILLER_64_1929 ();
 sg13g2_fill_2 FILLER_64_1935 ();
 sg13g2_decap_8 FILLER_64_1986 ();
 sg13g2_fill_2 FILLER_64_1993 ();
 sg13g2_decap_8 FILLER_64_1998 ();
 sg13g2_fill_2 FILLER_64_2005 ();
 sg13g2_fill_1 FILLER_64_2007 ();
 sg13g2_fill_2 FILLER_64_2012 ();
 sg13g2_fill_2 FILLER_64_2019 ();
 sg13g2_decap_4 FILLER_64_2025 ();
 sg13g2_fill_2 FILLER_64_2029 ();
 sg13g2_fill_2 FILLER_64_2048 ();
 sg13g2_fill_1 FILLER_64_2050 ();
 sg13g2_fill_2 FILLER_64_2057 ();
 sg13g2_fill_1 FILLER_64_2059 ();
 sg13g2_fill_1 FILLER_64_2072 ();
 sg13g2_fill_1 FILLER_64_2103 ();
 sg13g2_decap_4 FILLER_64_2153 ();
 sg13g2_fill_1 FILLER_64_2157 ();
 sg13g2_decap_8 FILLER_64_2162 ();
 sg13g2_fill_2 FILLER_64_2169 ();
 sg13g2_fill_1 FILLER_64_2171 ();
 sg13g2_fill_2 FILLER_64_2180 ();
 sg13g2_fill_1 FILLER_64_2211 ();
 sg13g2_fill_2 FILLER_64_2218 ();
 sg13g2_fill_1 FILLER_64_2252 ();
 sg13g2_fill_1 FILLER_64_2285 ();
 sg13g2_fill_1 FILLER_64_2291 ();
 sg13g2_fill_1 FILLER_64_2318 ();
 sg13g2_fill_2 FILLER_64_2332 ();
 sg13g2_fill_1 FILLER_64_2334 ();
 sg13g2_fill_2 FILLER_64_2341 ();
 sg13g2_fill_2 FILLER_64_2366 ();
 sg13g2_fill_2 FILLER_64_2372 ();
 sg13g2_fill_2 FILLER_64_2409 ();
 sg13g2_fill_1 FILLER_64_2430 ();
 sg13g2_fill_2 FILLER_64_2461 ();
 sg13g2_decap_8 FILLER_64_2468 ();
 sg13g2_decap_4 FILLER_64_2475 ();
 sg13g2_fill_1 FILLER_64_2479 ();
 sg13g2_decap_4 FILLER_64_2490 ();
 sg13g2_fill_1 FILLER_64_2494 ();
 sg13g2_decap_4 FILLER_64_2525 ();
 sg13g2_fill_1 FILLER_64_2529 ();
 sg13g2_decap_8 FILLER_64_2538 ();
 sg13g2_decap_8 FILLER_64_2545 ();
 sg13g2_decap_8 FILLER_64_2552 ();
 sg13g2_decap_8 FILLER_64_2559 ();
 sg13g2_decap_8 FILLER_64_2566 ();
 sg13g2_decap_8 FILLER_64_2573 ();
 sg13g2_decap_8 FILLER_64_2580 ();
 sg13g2_decap_8 FILLER_64_2587 ();
 sg13g2_decap_8 FILLER_64_2594 ();
 sg13g2_decap_8 FILLER_64_2601 ();
 sg13g2_decap_8 FILLER_64_2608 ();
 sg13g2_decap_8 FILLER_64_2615 ();
 sg13g2_decap_8 FILLER_64_2622 ();
 sg13g2_decap_8 FILLER_64_2629 ();
 sg13g2_decap_8 FILLER_64_2636 ();
 sg13g2_decap_8 FILLER_64_2643 ();
 sg13g2_decap_8 FILLER_64_2650 ();
 sg13g2_decap_8 FILLER_64_2657 ();
 sg13g2_decap_4 FILLER_64_2664 ();
 sg13g2_fill_2 FILLER_64_2668 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_51 ();
 sg13g2_fill_1 FILLER_65_58 ();
 sg13g2_fill_2 FILLER_65_68 ();
 sg13g2_fill_1 FILLER_65_75 ();
 sg13g2_fill_1 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_86 ();
 sg13g2_fill_1 FILLER_65_91 ();
 sg13g2_fill_2 FILLER_65_101 ();
 sg13g2_fill_2 FILLER_65_108 ();
 sg13g2_fill_1 FILLER_65_147 ();
 sg13g2_decap_4 FILLER_65_215 ();
 sg13g2_fill_2 FILLER_65_219 ();
 sg13g2_decap_8 FILLER_65_229 ();
 sg13g2_decap_4 FILLER_65_236 ();
 sg13g2_fill_1 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_272 ();
 sg13g2_decap_4 FILLER_65_286 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_decap_8 FILLER_65_327 ();
 sg13g2_decap_8 FILLER_65_334 ();
 sg13g2_fill_2 FILLER_65_341 ();
 sg13g2_fill_1 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_349 ();
 sg13g2_decap_4 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_360 ();
 sg13g2_fill_1 FILLER_65_373 ();
 sg13g2_fill_2 FILLER_65_384 ();
 sg13g2_fill_1 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_421 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_decap_8 FILLER_65_434 ();
 sg13g2_decap_8 FILLER_65_441 ();
 sg13g2_decap_4 FILLER_65_465 ();
 sg13g2_decap_8 FILLER_65_473 ();
 sg13g2_decap_8 FILLER_65_480 ();
 sg13g2_decap_8 FILLER_65_487 ();
 sg13g2_decap_4 FILLER_65_524 ();
 sg13g2_fill_1 FILLER_65_528 ();
 sg13g2_decap_8 FILLER_65_533 ();
 sg13g2_decap_4 FILLER_65_549 ();
 sg13g2_fill_2 FILLER_65_553 ();
 sg13g2_decap_8 FILLER_65_589 ();
 sg13g2_decap_8 FILLER_65_596 ();
 sg13g2_decap_8 FILLER_65_603 ();
 sg13g2_decap_8 FILLER_65_610 ();
 sg13g2_decap_4 FILLER_65_617 ();
 sg13g2_fill_1 FILLER_65_625 ();
 sg13g2_fill_2 FILLER_65_640 ();
 sg13g2_fill_1 FILLER_65_650 ();
 sg13g2_fill_1 FILLER_65_659 ();
 sg13g2_fill_1 FILLER_65_666 ();
 sg13g2_fill_1 FILLER_65_685 ();
 sg13g2_decap_8 FILLER_65_691 ();
 sg13g2_decap_4 FILLER_65_702 ();
 sg13g2_fill_2 FILLER_65_706 ();
 sg13g2_decap_8 FILLER_65_712 ();
 sg13g2_decap_8 FILLER_65_719 ();
 sg13g2_decap_4 FILLER_65_726 ();
 sg13g2_fill_2 FILLER_65_730 ();
 sg13g2_fill_1 FILLER_65_737 ();
 sg13g2_fill_2 FILLER_65_746 ();
 sg13g2_fill_1 FILLER_65_748 ();
 sg13g2_decap_8 FILLER_65_753 ();
 sg13g2_fill_1 FILLER_65_760 ();
 sg13g2_fill_2 FILLER_65_776 ();
 sg13g2_fill_1 FILLER_65_778 ();
 sg13g2_decap_4 FILLER_65_783 ();
 sg13g2_fill_1 FILLER_65_787 ();
 sg13g2_decap_8 FILLER_65_793 ();
 sg13g2_decap_8 FILLER_65_800 ();
 sg13g2_fill_2 FILLER_65_820 ();
 sg13g2_decap_8 FILLER_65_832 ();
 sg13g2_fill_2 FILLER_65_839 ();
 sg13g2_fill_2 FILLER_65_872 ();
 sg13g2_decap_4 FILLER_65_882 ();
 sg13g2_fill_2 FILLER_65_886 ();
 sg13g2_decap_8 FILLER_65_931 ();
 sg13g2_decap_8 FILLER_65_938 ();
 sg13g2_decap_8 FILLER_65_945 ();
 sg13g2_decap_8 FILLER_65_952 ();
 sg13g2_decap_4 FILLER_65_959 ();
 sg13g2_fill_2 FILLER_65_963 ();
 sg13g2_decap_8 FILLER_65_970 ();
 sg13g2_fill_2 FILLER_65_977 ();
 sg13g2_decap_8 FILLER_65_983 ();
 sg13g2_decap_8 FILLER_65_994 ();
 sg13g2_fill_2 FILLER_65_1001 ();
 sg13g2_fill_1 FILLER_65_1003 ();
 sg13g2_fill_1 FILLER_65_1010 ();
 sg13g2_fill_2 FILLER_65_1017 ();
 sg13g2_fill_1 FILLER_65_1019 ();
 sg13g2_decap_4 FILLER_65_1024 ();
 sg13g2_fill_1 FILLER_65_1028 ();
 sg13g2_fill_2 FILLER_65_1034 ();
 sg13g2_fill_2 FILLER_65_1087 ();
 sg13g2_fill_2 FILLER_65_1143 ();
 sg13g2_fill_1 FILLER_65_1145 ();
 sg13g2_decap_8 FILLER_65_1151 ();
 sg13g2_decap_8 FILLER_65_1158 ();
 sg13g2_fill_1 FILLER_65_1165 ();
 sg13g2_fill_2 FILLER_65_1196 ();
 sg13g2_fill_1 FILLER_65_1198 ();
 sg13g2_fill_1 FILLER_65_1234 ();
 sg13g2_fill_1 FILLER_65_1246 ();
 sg13g2_fill_2 FILLER_65_1253 ();
 sg13g2_fill_1 FILLER_65_1255 ();
 sg13g2_decap_4 FILLER_65_1264 ();
 sg13g2_fill_1 FILLER_65_1296 ();
 sg13g2_decap_4 FILLER_65_1313 ();
 sg13g2_fill_2 FILLER_65_1373 ();
 sg13g2_fill_1 FILLER_65_1391 ();
 sg13g2_fill_1 FILLER_65_1406 ();
 sg13g2_fill_2 FILLER_65_1443 ();
 sg13g2_fill_1 FILLER_65_1445 ();
 sg13g2_decap_8 FILLER_65_1450 ();
 sg13g2_decap_4 FILLER_65_1457 ();
 sg13g2_fill_2 FILLER_65_1461 ();
 sg13g2_fill_1 FILLER_65_1466 ();
 sg13g2_fill_1 FILLER_65_1481 ();
 sg13g2_fill_2 FILLER_65_1594 ();
 sg13g2_fill_1 FILLER_65_1596 ();
 sg13g2_fill_2 FILLER_65_1606 ();
 sg13g2_fill_1 FILLER_65_1617 ();
 sg13g2_fill_1 FILLER_65_1652 ();
 sg13g2_decap_4 FILLER_65_1658 ();
 sg13g2_decap_8 FILLER_65_1688 ();
 sg13g2_decap_8 FILLER_65_1695 ();
 sg13g2_decap_8 FILLER_65_1702 ();
 sg13g2_decap_8 FILLER_65_1715 ();
 sg13g2_fill_2 FILLER_65_1722 ();
 sg13g2_fill_1 FILLER_65_1724 ();
 sg13g2_decap_4 FILLER_65_1730 ();
 sg13g2_fill_1 FILLER_65_1734 ();
 sg13g2_fill_2 FILLER_65_1761 ();
 sg13g2_fill_1 FILLER_65_1763 ();
 sg13g2_fill_1 FILLER_65_1782 ();
 sg13g2_fill_2 FILLER_65_1797 ();
 sg13g2_decap_8 FILLER_65_1803 ();
 sg13g2_decap_8 FILLER_65_1810 ();
 sg13g2_decap_8 FILLER_65_1817 ();
 sg13g2_decap_4 FILLER_65_1824 ();
 sg13g2_fill_2 FILLER_65_1828 ();
 sg13g2_fill_1 FILLER_65_1848 ();
 sg13g2_decap_8 FILLER_65_1894 ();
 sg13g2_decap_8 FILLER_65_1901 ();
 sg13g2_decap_8 FILLER_65_1908 ();
 sg13g2_decap_8 FILLER_65_1915 ();
 sg13g2_decap_8 FILLER_65_1922 ();
 sg13g2_decap_8 FILLER_65_1929 ();
 sg13g2_fill_2 FILLER_65_1936 ();
 sg13g2_fill_2 FILLER_65_1944 ();
 sg13g2_fill_1 FILLER_65_1946 ();
 sg13g2_decap_4 FILLER_65_1953 ();
 sg13g2_decap_8 FILLER_65_1963 ();
 sg13g2_decap_8 FILLER_65_1970 ();
 sg13g2_fill_2 FILLER_65_1977 ();
 sg13g2_fill_1 FILLER_65_1979 ();
 sg13g2_fill_1 FILLER_65_2001 ();
 sg13g2_fill_2 FILLER_65_2007 ();
 sg13g2_fill_2 FILLER_65_2035 ();
 sg13g2_fill_1 FILLER_65_2037 ();
 sg13g2_fill_2 FILLER_65_2128 ();
 sg13g2_fill_1 FILLER_65_2130 ();
 sg13g2_fill_2 FILLER_65_2140 ();
 sg13g2_decap_4 FILLER_65_2156 ();
 sg13g2_fill_1 FILLER_65_2186 ();
 sg13g2_fill_1 FILLER_65_2200 ();
 sg13g2_fill_2 FILLER_65_2228 ();
 sg13g2_fill_2 FILLER_65_2248 ();
 sg13g2_fill_2 FILLER_65_2256 ();
 sg13g2_decap_8 FILLER_65_2270 ();
 sg13g2_fill_2 FILLER_65_2277 ();
 sg13g2_fill_1 FILLER_65_2279 ();
 sg13g2_decap_4 FILLER_65_2293 ();
 sg13g2_fill_1 FILLER_65_2302 ();
 sg13g2_decap_8 FILLER_65_2307 ();
 sg13g2_fill_1 FILLER_65_2314 ();
 sg13g2_decap_8 FILLER_65_2341 ();
 sg13g2_decap_8 FILLER_65_2348 ();
 sg13g2_decap_8 FILLER_65_2355 ();
 sg13g2_fill_1 FILLER_65_2367 ();
 sg13g2_decap_4 FILLER_65_2382 ();
 sg13g2_fill_1 FILLER_65_2386 ();
 sg13g2_decap_4 FILLER_65_2413 ();
 sg13g2_fill_2 FILLER_65_2421 ();
 sg13g2_fill_2 FILLER_65_2449 ();
 sg13g2_fill_1 FILLER_65_2451 ();
 sg13g2_fill_2 FILLER_65_2456 ();
 sg13g2_fill_1 FILLER_65_2458 ();
 sg13g2_decap_8 FILLER_65_2485 ();
 sg13g2_fill_2 FILLER_65_2492 ();
 sg13g2_decap_8 FILLER_65_2521 ();
 sg13g2_decap_8 FILLER_65_2528 ();
 sg13g2_decap_8 FILLER_65_2535 ();
 sg13g2_decap_8 FILLER_65_2542 ();
 sg13g2_decap_8 FILLER_65_2549 ();
 sg13g2_decap_8 FILLER_65_2556 ();
 sg13g2_decap_8 FILLER_65_2563 ();
 sg13g2_decap_8 FILLER_65_2570 ();
 sg13g2_decap_8 FILLER_65_2577 ();
 sg13g2_decap_8 FILLER_65_2584 ();
 sg13g2_decap_8 FILLER_65_2591 ();
 sg13g2_decap_8 FILLER_65_2598 ();
 sg13g2_decap_8 FILLER_65_2605 ();
 sg13g2_decap_8 FILLER_65_2612 ();
 sg13g2_decap_8 FILLER_65_2619 ();
 sg13g2_decap_8 FILLER_65_2626 ();
 sg13g2_decap_8 FILLER_65_2633 ();
 sg13g2_decap_8 FILLER_65_2640 ();
 sg13g2_decap_8 FILLER_65_2647 ();
 sg13g2_decap_8 FILLER_65_2654 ();
 sg13g2_decap_8 FILLER_65_2661 ();
 sg13g2_fill_2 FILLER_65_2668 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_fill_1 FILLER_66_45 ();
 sg13g2_fill_2 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_76 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_107 ();
 sg13g2_fill_1 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_167 ();
 sg13g2_decap_4 FILLER_66_182 ();
 sg13g2_fill_2 FILLER_66_186 ();
 sg13g2_fill_1 FILLER_66_206 ();
 sg13g2_fill_1 FILLER_66_213 ();
 sg13g2_fill_2 FILLER_66_217 ();
 sg13g2_fill_1 FILLER_66_219 ();
 sg13g2_decap_8 FILLER_66_225 ();
 sg13g2_decap_8 FILLER_66_232 ();
 sg13g2_decap_4 FILLER_66_239 ();
 sg13g2_fill_1 FILLER_66_243 ();
 sg13g2_decap_4 FILLER_66_264 ();
 sg13g2_fill_2 FILLER_66_268 ();
 sg13g2_decap_8 FILLER_66_274 ();
 sg13g2_decap_8 FILLER_66_281 ();
 sg13g2_decap_8 FILLER_66_293 ();
 sg13g2_decap_4 FILLER_66_313 ();
 sg13g2_fill_2 FILLER_66_317 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_fill_1 FILLER_66_383 ();
 sg13g2_fill_1 FILLER_66_390 ();
 sg13g2_fill_1 FILLER_66_396 ();
 sg13g2_decap_4 FILLER_66_416 ();
 sg13g2_decap_8 FILLER_66_426 ();
 sg13g2_decap_4 FILLER_66_433 ();
 sg13g2_fill_1 FILLER_66_437 ();
 sg13g2_decap_8 FILLER_66_464 ();
 sg13g2_fill_2 FILLER_66_475 ();
 sg13g2_fill_2 FILLER_66_481 ();
 sg13g2_fill_1 FILLER_66_483 ();
 sg13g2_fill_2 FILLER_66_489 ();
 sg13g2_fill_1 FILLER_66_491 ();
 sg13g2_decap_4 FILLER_66_496 ();
 sg13g2_fill_1 FILLER_66_500 ();
 sg13g2_decap_8 FILLER_66_504 ();
 sg13g2_fill_2 FILLER_66_511 ();
 sg13g2_fill_2 FILLER_66_539 ();
 sg13g2_decap_8 FILLER_66_553 ();
 sg13g2_fill_1 FILLER_66_560 ();
 sg13g2_decap_8 FILLER_66_566 ();
 sg13g2_fill_2 FILLER_66_573 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_decap_8 FILLER_66_598 ();
 sg13g2_decap_8 FILLER_66_605 ();
 sg13g2_decap_8 FILLER_66_612 ();
 sg13g2_fill_2 FILLER_66_644 ();
 sg13g2_fill_2 FILLER_66_722 ();
 sg13g2_decap_8 FILLER_66_745 ();
 sg13g2_fill_1 FILLER_66_752 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_4 FILLER_66_786 ();
 sg13g2_fill_1 FILLER_66_790 ();
 sg13g2_decap_8 FILLER_66_804 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_8 FILLER_66_857 ();
 sg13g2_decap_8 FILLER_66_864 ();
 sg13g2_decap_8 FILLER_66_871 ();
 sg13g2_decap_8 FILLER_66_878 ();
 sg13g2_fill_2 FILLER_66_885 ();
 sg13g2_decap_8 FILLER_66_897 ();
 sg13g2_fill_1 FILLER_66_904 ();
 sg13g2_fill_2 FILLER_66_914 ();
 sg13g2_fill_1 FILLER_66_916 ();
 sg13g2_fill_1 FILLER_66_943 ();
 sg13g2_decap_8 FILLER_66_986 ();
 sg13g2_decap_8 FILLER_66_993 ();
 sg13g2_decap_4 FILLER_66_1000 ();
 sg13g2_fill_1 FILLER_66_1008 ();
 sg13g2_fill_2 FILLER_66_1015 ();
 sg13g2_fill_1 FILLER_66_1020 ();
 sg13g2_fill_2 FILLER_66_1026 ();
 sg13g2_fill_1 FILLER_66_1092 ();
 sg13g2_fill_2 FILLER_66_1111 ();
 sg13g2_decap_8 FILLER_66_1118 ();
 sg13g2_fill_2 FILLER_66_1202 ();
 sg13g2_fill_1 FILLER_66_1204 ();
 sg13g2_decap_4 FILLER_66_1243 ();
 sg13g2_fill_1 FILLER_66_1247 ();
 sg13g2_fill_1 FILLER_66_1252 ();
 sg13g2_decap_8 FILLER_66_1265 ();
 sg13g2_decap_8 FILLER_66_1272 ();
 sg13g2_decap_8 FILLER_66_1279 ();
 sg13g2_fill_1 FILLER_66_1286 ();
 sg13g2_fill_2 FILLER_66_1291 ();
 sg13g2_decap_8 FILLER_66_1311 ();
 sg13g2_decap_8 FILLER_66_1318 ();
 sg13g2_fill_2 FILLER_66_1325 ();
 sg13g2_fill_1 FILLER_66_1327 ();
 sg13g2_fill_1 FILLER_66_1369 ();
 sg13g2_fill_1 FILLER_66_1375 ();
 sg13g2_decap_4 FILLER_66_1420 ();
 sg13g2_fill_2 FILLER_66_1424 ();
 sg13g2_fill_2 FILLER_66_1435 ();
 sg13g2_decap_4 FILLER_66_1469 ();
 sg13g2_fill_1 FILLER_66_1473 ();
 sg13g2_decap_8 FILLER_66_1500 ();
 sg13g2_fill_1 FILLER_66_1507 ();
 sg13g2_fill_1 FILLER_66_1537 ();
 sg13g2_fill_2 FILLER_66_1547 ();
 sg13g2_fill_2 FILLER_66_1555 ();
 sg13g2_decap_4 FILLER_66_1565 ();
 sg13g2_fill_1 FILLER_66_1643 ();
 sg13g2_decap_8 FILLER_66_1649 ();
 sg13g2_fill_2 FILLER_66_1656 ();
 sg13g2_fill_1 FILLER_66_1658 ();
 sg13g2_decap_8 FILLER_66_1664 ();
 sg13g2_decap_8 FILLER_66_1671 ();
 sg13g2_fill_1 FILLER_66_1678 ();
 sg13g2_fill_2 FILLER_66_1691 ();
 sg13g2_decap_4 FILLER_66_1700 ();
 sg13g2_fill_2 FILLER_66_1704 ();
 sg13g2_decap_8 FILLER_66_1714 ();
 sg13g2_decap_8 FILLER_66_1721 ();
 sg13g2_decap_8 FILLER_66_1728 ();
 sg13g2_decap_8 FILLER_66_1735 ();
 sg13g2_fill_2 FILLER_66_1742 ();
 sg13g2_fill_2 FILLER_66_1754 ();
 sg13g2_fill_1 FILLER_66_1756 ();
 sg13g2_decap_4 FILLER_66_1800 ();
 sg13g2_decap_8 FILLER_66_1814 ();
 sg13g2_decap_4 FILLER_66_1821 ();
 sg13g2_fill_2 FILLER_66_1825 ();
 sg13g2_fill_1 FILLER_66_1839 ();
 sg13g2_decap_8 FILLER_66_1866 ();
 sg13g2_decap_8 FILLER_66_1873 ();
 sg13g2_decap_8 FILLER_66_1880 ();
 sg13g2_decap_8 FILLER_66_1887 ();
 sg13g2_fill_1 FILLER_66_1894 ();
 sg13g2_decap_4 FILLER_66_1931 ();
 sg13g2_fill_2 FILLER_66_1935 ();
 sg13g2_decap_4 FILLER_66_1943 ();
 sg13g2_decap_8 FILLER_66_1951 ();
 sg13g2_decap_8 FILLER_66_1958 ();
 sg13g2_decap_4 FILLER_66_1965 ();
 sg13g2_fill_1 FILLER_66_1969 ();
 sg13g2_decap_8 FILLER_66_2027 ();
 sg13g2_decap_8 FILLER_66_2034 ();
 sg13g2_fill_2 FILLER_66_2041 ();
 sg13g2_fill_1 FILLER_66_2043 ();
 sg13g2_decap_8 FILLER_66_2059 ();
 sg13g2_decap_8 FILLER_66_2066 ();
 sg13g2_decap_4 FILLER_66_2073 ();
 sg13g2_fill_2 FILLER_66_2077 ();
 sg13g2_fill_2 FILLER_66_2084 ();
 sg13g2_fill_2 FILLER_66_2099 ();
 sg13g2_fill_2 FILLER_66_2106 ();
 sg13g2_fill_2 FILLER_66_2116 ();
 sg13g2_fill_1 FILLER_66_2118 ();
 sg13g2_decap_8 FILLER_66_2133 ();
 sg13g2_decap_8 FILLER_66_2140 ();
 sg13g2_decap_8 FILLER_66_2147 ();
 sg13g2_decap_8 FILLER_66_2154 ();
 sg13g2_fill_1 FILLER_66_2161 ();
 sg13g2_fill_2 FILLER_66_2170 ();
 sg13g2_fill_1 FILLER_66_2184 ();
 sg13g2_fill_2 FILLER_66_2215 ();
 sg13g2_fill_1 FILLER_66_2226 ();
 sg13g2_fill_2 FILLER_66_2267 ();
 sg13g2_decap_8 FILLER_66_2278 ();
 sg13g2_decap_8 FILLER_66_2285 ();
 sg13g2_decap_8 FILLER_66_2292 ();
 sg13g2_fill_2 FILLER_66_2299 ();
 sg13g2_fill_1 FILLER_66_2313 ();
 sg13g2_decap_4 FILLER_66_2327 ();
 sg13g2_decap_8 FILLER_66_2338 ();
 sg13g2_decap_8 FILLER_66_2345 ();
 sg13g2_fill_2 FILLER_66_2352 ();
 sg13g2_decap_8 FILLER_66_2406 ();
 sg13g2_decap_8 FILLER_66_2413 ();
 sg13g2_decap_8 FILLER_66_2420 ();
 sg13g2_fill_2 FILLER_66_2427 ();
 sg13g2_decap_8 FILLER_66_2433 ();
 sg13g2_decap_4 FILLER_66_2440 ();
 sg13g2_fill_2 FILLER_66_2444 ();
 sg13g2_fill_1 FILLER_66_2460 ();
 sg13g2_decap_4 FILLER_66_2487 ();
 sg13g2_fill_2 FILLER_66_2491 ();
 sg13g2_decap_8 FILLER_66_2533 ();
 sg13g2_decap_8 FILLER_66_2540 ();
 sg13g2_decap_8 FILLER_66_2547 ();
 sg13g2_decap_8 FILLER_66_2554 ();
 sg13g2_decap_8 FILLER_66_2561 ();
 sg13g2_decap_8 FILLER_66_2568 ();
 sg13g2_decap_8 FILLER_66_2575 ();
 sg13g2_decap_8 FILLER_66_2582 ();
 sg13g2_decap_8 FILLER_66_2589 ();
 sg13g2_decap_8 FILLER_66_2596 ();
 sg13g2_decap_8 FILLER_66_2603 ();
 sg13g2_decap_8 FILLER_66_2610 ();
 sg13g2_decap_8 FILLER_66_2617 ();
 sg13g2_decap_8 FILLER_66_2624 ();
 sg13g2_decap_8 FILLER_66_2631 ();
 sg13g2_decap_8 FILLER_66_2638 ();
 sg13g2_decap_8 FILLER_66_2645 ();
 sg13g2_decap_8 FILLER_66_2652 ();
 sg13g2_decap_8 FILLER_66_2659 ();
 sg13g2_decap_4 FILLER_66_2666 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_fill_1 FILLER_67_25 ();
 sg13g2_fill_1 FILLER_67_31 ();
 sg13g2_fill_1 FILLER_67_36 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_48 ();
 sg13g2_fill_1 FILLER_67_50 ();
 sg13g2_fill_2 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_68 ();
 sg13g2_fill_1 FILLER_67_74 ();
 sg13g2_fill_1 FILLER_67_99 ();
 sg13g2_fill_2 FILLER_67_105 ();
 sg13g2_fill_2 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_135 ();
 sg13g2_fill_1 FILLER_67_142 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_fill_2 FILLER_67_176 ();
 sg13g2_decap_4 FILLER_67_192 ();
 sg13g2_fill_1 FILLER_67_196 ();
 sg13g2_fill_1 FILLER_67_217 ();
 sg13g2_decap_4 FILLER_67_222 ();
 sg13g2_decap_8 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_241 ();
 sg13g2_fill_2 FILLER_67_248 ();
 sg13g2_fill_2 FILLER_67_261 ();
 sg13g2_fill_1 FILLER_67_263 ();
 sg13g2_decap_8 FILLER_67_270 ();
 sg13g2_decap_4 FILLER_67_277 ();
 sg13g2_decap_8 FILLER_67_286 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_decap_8 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_338 ();
 sg13g2_decap_4 FILLER_67_345 ();
 sg13g2_fill_1 FILLER_67_349 ();
 sg13g2_fill_1 FILLER_67_371 ();
 sg13g2_fill_1 FILLER_67_378 ();
 sg13g2_fill_1 FILLER_67_384 ();
 sg13g2_fill_1 FILLER_67_390 ();
 sg13g2_fill_1 FILLER_67_396 ();
 sg13g2_fill_1 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_407 ();
 sg13g2_fill_1 FILLER_67_415 ();
 sg13g2_decap_8 FILLER_67_421 ();
 sg13g2_decap_8 FILLER_67_428 ();
 sg13g2_fill_2 FILLER_67_435 ();
 sg13g2_fill_1 FILLER_67_437 ();
 sg13g2_fill_1 FILLER_67_480 ();
 sg13g2_fill_1 FILLER_67_486 ();
 sg13g2_fill_1 FILLER_67_492 ();
 sg13g2_fill_1 FILLER_67_498 ();
 sg13g2_decap_8 FILLER_67_509 ();
 sg13g2_decap_4 FILLER_67_516 ();
 sg13g2_fill_2 FILLER_67_520 ();
 sg13g2_decap_8 FILLER_67_532 ();
 sg13g2_decap_4 FILLER_67_539 ();
 sg13g2_fill_1 FILLER_67_548 ();
 sg13g2_fill_2 FILLER_67_554 ();
 sg13g2_fill_1 FILLER_67_556 ();
 sg13g2_fill_2 FILLER_67_567 ();
 sg13g2_fill_1 FILLER_67_569 ();
 sg13g2_decap_4 FILLER_67_581 ();
 sg13g2_fill_2 FILLER_67_585 ();
 sg13g2_decap_8 FILLER_67_590 ();
 sg13g2_fill_1 FILLER_67_597 ();
 sg13g2_decap_8 FILLER_67_605 ();
 sg13g2_fill_2 FILLER_67_612 ();
 sg13g2_fill_1 FILLER_67_614 ();
 sg13g2_fill_2 FILLER_67_620 ();
 sg13g2_fill_1 FILLER_67_622 ();
 sg13g2_fill_2 FILLER_67_636 ();
 sg13g2_fill_2 FILLER_67_665 ();
 sg13g2_fill_1 FILLER_67_673 ();
 sg13g2_decap_8 FILLER_67_683 ();
 sg13g2_fill_2 FILLER_67_708 ();
 sg13g2_fill_2 FILLER_67_723 ();
 sg13g2_fill_1 FILLER_67_725 ();
 sg13g2_decap_8 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_743 ();
 sg13g2_fill_1 FILLER_67_750 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_fill_1 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_fill_1 FILLER_67_816 ();
 sg13g2_fill_1 FILLER_67_835 ();
 sg13g2_decap_8 FILLER_67_872 ();
 sg13g2_decap_8 FILLER_67_879 ();
 sg13g2_decap_4 FILLER_67_886 ();
 sg13g2_fill_1 FILLER_67_890 ();
 sg13g2_fill_1 FILLER_67_907 ();
 sg13g2_decap_8 FILLER_67_934 ();
 sg13g2_decap_4 FILLER_67_949 ();
 sg13g2_fill_2 FILLER_67_962 ();
 sg13g2_fill_1 FILLER_67_970 ();
 sg13g2_fill_2 FILLER_67_989 ();
 sg13g2_decap_4 FILLER_67_995 ();
 sg13g2_fill_1 FILLER_67_999 ();
 sg13g2_fill_2 FILLER_67_1008 ();
 sg13g2_fill_1 FILLER_67_1010 ();
 sg13g2_fill_1 FILLER_67_1055 ();
 sg13g2_fill_2 FILLER_67_1062 ();
 sg13g2_fill_2 FILLER_67_1102 ();
 sg13g2_decap_8 FILLER_67_1110 ();
 sg13g2_decap_8 FILLER_67_1117 ();
 sg13g2_fill_1 FILLER_67_1124 ();
 sg13g2_fill_2 FILLER_67_1137 ();
 sg13g2_fill_1 FILLER_67_1139 ();
 sg13g2_decap_4 FILLER_67_1150 ();
 sg13g2_decap_8 FILLER_67_1158 ();
 sg13g2_decap_4 FILLER_67_1165 ();
 sg13g2_fill_1 FILLER_67_1169 ();
 sg13g2_fill_2 FILLER_67_1179 ();
 sg13g2_fill_1 FILLER_67_1181 ();
 sg13g2_fill_1 FILLER_67_1188 ();
 sg13g2_fill_2 FILLER_67_1197 ();
 sg13g2_fill_1 FILLER_67_1229 ();
 sg13g2_decap_8 FILLER_67_1234 ();
 sg13g2_fill_2 FILLER_67_1241 ();
 sg13g2_fill_1 FILLER_67_1243 ();
 sg13g2_decap_8 FILLER_67_1276 ();
 sg13g2_fill_2 FILLER_67_1283 ();
 sg13g2_fill_2 FILLER_67_1290 ();
 sg13g2_fill_1 FILLER_67_1292 ();
 sg13g2_decap_8 FILLER_67_1305 ();
 sg13g2_fill_2 FILLER_67_1312 ();
 sg13g2_fill_1 FILLER_67_1314 ();
 sg13g2_decap_8 FILLER_67_1322 ();
 sg13g2_fill_2 FILLER_67_1329 ();
 sg13g2_fill_1 FILLER_67_1331 ();
 sg13g2_decap_8 FILLER_67_1335 ();
 sg13g2_decap_8 FILLER_67_1346 ();
 sg13g2_decap_8 FILLER_67_1353 ();
 sg13g2_fill_2 FILLER_67_1365 ();
 sg13g2_fill_1 FILLER_67_1367 ();
 sg13g2_fill_2 FILLER_67_1387 ();
 sg13g2_fill_1 FILLER_67_1389 ();
 sg13g2_fill_2 FILLER_67_1407 ();
 sg13g2_decap_8 FILLER_67_1435 ();
 sg13g2_decap_4 FILLER_67_1442 ();
 sg13g2_decap_8 FILLER_67_1454 ();
 sg13g2_decap_8 FILLER_67_1461 ();
 sg13g2_fill_1 FILLER_67_1468 ();
 sg13g2_fill_2 FILLER_67_1473 ();
 sg13g2_fill_1 FILLER_67_1475 ();
 sg13g2_fill_1 FILLER_67_1483 ();
 sg13g2_decap_8 FILLER_67_1501 ();
 sg13g2_fill_2 FILLER_67_1508 ();
 sg13g2_fill_1 FILLER_67_1510 ();
 sg13g2_fill_1 FILLER_67_1515 ();
 sg13g2_decap_8 FILLER_67_1531 ();
 sg13g2_decap_8 FILLER_67_1538 ();
 sg13g2_decap_8 FILLER_67_1545 ();
 sg13g2_decap_8 FILLER_67_1563 ();
 sg13g2_fill_1 FILLER_67_1599 ();
 sg13g2_fill_1 FILLER_67_1624 ();
 sg13g2_fill_1 FILLER_67_1638 ();
 sg13g2_decap_4 FILLER_67_1664 ();
 sg13g2_fill_1 FILLER_67_1674 ();
 sg13g2_fill_1 FILLER_67_1684 ();
 sg13g2_fill_1 FILLER_67_1690 ();
 sg13g2_fill_2 FILLER_67_1699 ();
 sg13g2_decap_8 FILLER_67_1707 ();
 sg13g2_decap_4 FILLER_67_1714 ();
 sg13g2_decap_8 FILLER_67_1722 ();
 sg13g2_fill_2 FILLER_67_1729 ();
 sg13g2_fill_2 FILLER_67_1777 ();
 sg13g2_fill_2 FILLER_67_1808 ();
 sg13g2_fill_1 FILLER_67_1810 ();
 sg13g2_decap_4 FILLER_67_1840 ();
 sg13g2_decap_4 FILLER_67_1868 ();
 sg13g2_fill_1 FILLER_67_1876 ();
 sg13g2_decap_4 FILLER_67_1883 ();
 sg13g2_fill_1 FILLER_67_1887 ();
 sg13g2_fill_1 FILLER_67_1897 ();
 sg13g2_decap_4 FILLER_67_1903 ();
 sg13g2_fill_1 FILLER_67_1907 ();
 sg13g2_fill_2 FILLER_67_1934 ();
 sg13g2_fill_1 FILLER_67_1941 ();
 sg13g2_fill_2 FILLER_67_1968 ();
 sg13g2_decap_8 FILLER_67_1996 ();
 sg13g2_decap_8 FILLER_67_2003 ();
 sg13g2_decap_8 FILLER_67_2010 ();
 sg13g2_decap_8 FILLER_67_2017 ();
 sg13g2_decap_8 FILLER_67_2024 ();
 sg13g2_decap_8 FILLER_67_2031 ();
 sg13g2_decap_4 FILLER_67_2038 ();
 sg13g2_fill_2 FILLER_67_2042 ();
 sg13g2_decap_8 FILLER_67_2050 ();
 sg13g2_decap_4 FILLER_67_2057 ();
 sg13g2_fill_2 FILLER_67_2061 ();
 sg13g2_fill_2 FILLER_67_2096 ();
 sg13g2_decap_8 FILLER_67_2159 ();
 sg13g2_decap_4 FILLER_67_2166 ();
 sg13g2_fill_2 FILLER_67_2170 ();
 sg13g2_fill_2 FILLER_67_2225 ();
 sg13g2_fill_1 FILLER_67_2256 ();
 sg13g2_fill_1 FILLER_67_2301 ();
 sg13g2_fill_1 FILLER_67_2360 ();
 sg13g2_fill_1 FILLER_67_2364 ();
 sg13g2_decap_8 FILLER_67_2384 ();
 sg13g2_decap_8 FILLER_67_2391 ();
 sg13g2_decap_8 FILLER_67_2398 ();
 sg13g2_decap_8 FILLER_67_2405 ();
 sg13g2_decap_8 FILLER_67_2412 ();
 sg13g2_decap_4 FILLER_67_2419 ();
 sg13g2_fill_1 FILLER_67_2423 ();
 sg13g2_decap_8 FILLER_67_2438 ();
 sg13g2_decap_8 FILLER_67_2445 ();
 sg13g2_decap_4 FILLER_67_2452 ();
 sg13g2_fill_1 FILLER_67_2456 ();
 sg13g2_decap_8 FILLER_67_2461 ();
 sg13g2_fill_1 FILLER_67_2468 ();
 sg13g2_decap_4 FILLER_67_2473 ();
 sg13g2_fill_1 FILLER_67_2477 ();
 sg13g2_decap_4 FILLER_67_2482 ();
 sg13g2_fill_2 FILLER_67_2486 ();
 sg13g2_fill_1 FILLER_67_2505 ();
 sg13g2_decap_8 FILLER_67_2532 ();
 sg13g2_decap_8 FILLER_67_2539 ();
 sg13g2_decap_8 FILLER_67_2546 ();
 sg13g2_decap_8 FILLER_67_2553 ();
 sg13g2_decap_8 FILLER_67_2560 ();
 sg13g2_decap_8 FILLER_67_2567 ();
 sg13g2_decap_8 FILLER_67_2574 ();
 sg13g2_decap_8 FILLER_67_2581 ();
 sg13g2_decap_8 FILLER_67_2588 ();
 sg13g2_decap_8 FILLER_67_2595 ();
 sg13g2_decap_8 FILLER_67_2602 ();
 sg13g2_decap_8 FILLER_67_2609 ();
 sg13g2_decap_8 FILLER_67_2616 ();
 sg13g2_decap_8 FILLER_67_2623 ();
 sg13g2_decap_8 FILLER_67_2630 ();
 sg13g2_decap_8 FILLER_67_2637 ();
 sg13g2_decap_8 FILLER_67_2644 ();
 sg13g2_decap_8 FILLER_67_2651 ();
 sg13g2_decap_8 FILLER_67_2658 ();
 sg13g2_decap_4 FILLER_67_2665 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_19 ();
 sg13g2_fill_1 FILLER_68_26 ();
 sg13g2_decap_4 FILLER_68_41 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_fill_1 FILLER_68_88 ();
 sg13g2_decap_4 FILLER_68_94 ();
 sg13g2_fill_1 FILLER_68_104 ();
 sg13g2_fill_2 FILLER_68_115 ();
 sg13g2_fill_1 FILLER_68_117 ();
 sg13g2_decap_4 FILLER_68_122 ();
 sg13g2_fill_1 FILLER_68_126 ();
 sg13g2_decap_4 FILLER_68_132 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_fill_2 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_145 ();
 sg13g2_fill_2 FILLER_68_167 ();
 sg13g2_decap_4 FILLER_68_174 ();
 sg13g2_decap_8 FILLER_68_194 ();
 sg13g2_fill_1 FILLER_68_201 ();
 sg13g2_decap_8 FILLER_68_206 ();
 sg13g2_decap_8 FILLER_68_213 ();
 sg13g2_decap_8 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_229 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_4 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_decap_8 FILLER_68_268 ();
 sg13g2_decap_8 FILLER_68_275 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_decap_8 FILLER_68_289 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_decap_8 FILLER_68_310 ();
 sg13g2_decap_8 FILLER_68_317 ();
 sg13g2_decap_8 FILLER_68_324 ();
 sg13g2_decap_8 FILLER_68_331 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_409 ();
 sg13g2_fill_1 FILLER_68_431 ();
 sg13g2_fill_1 FILLER_68_441 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_8 FILLER_68_453 ();
 sg13g2_decap_8 FILLER_68_460 ();
 sg13g2_decap_4 FILLER_68_467 ();
 sg13g2_fill_2 FILLER_68_471 ();
 sg13g2_fill_2 FILLER_68_510 ();
 sg13g2_fill_2 FILLER_68_517 ();
 sg13g2_fill_1 FILLER_68_519 ();
 sg13g2_decap_8 FILLER_68_525 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_4 FILLER_68_539 ();
 sg13g2_decap_8 FILLER_68_547 ();
 sg13g2_decap_8 FILLER_68_554 ();
 sg13g2_decap_4 FILLER_68_561 ();
 sg13g2_fill_1 FILLER_68_600 ();
 sg13g2_fill_2 FILLER_68_612 ();
 sg13g2_fill_2 FILLER_68_623 ();
 sg13g2_fill_1 FILLER_68_625 ();
 sg13g2_fill_2 FILLER_68_637 ();
 sg13g2_fill_1 FILLER_68_639 ();
 sg13g2_decap_4 FILLER_68_644 ();
 sg13g2_decap_8 FILLER_68_660 ();
 sg13g2_decap_8 FILLER_68_667 ();
 sg13g2_fill_1 FILLER_68_674 ();
 sg13g2_decap_4 FILLER_68_680 ();
 sg13g2_fill_2 FILLER_68_684 ();
 sg13g2_fill_1 FILLER_68_734 ();
 sg13g2_decap_8 FILLER_68_750 ();
 sg13g2_fill_1 FILLER_68_757 ();
 sg13g2_decap_8 FILLER_68_771 ();
 sg13g2_fill_1 FILLER_68_778 ();
 sg13g2_fill_1 FILLER_68_783 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_fill_1 FILLER_68_846 ();
 sg13g2_decap_4 FILLER_68_853 ();
 sg13g2_fill_1 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_888 ();
 sg13g2_decap_8 FILLER_68_897 ();
 sg13g2_decap_8 FILLER_68_904 ();
 sg13g2_fill_1 FILLER_68_911 ();
 sg13g2_decap_8 FILLER_68_925 ();
 sg13g2_fill_2 FILLER_68_944 ();
 sg13g2_decap_4 FILLER_68_952 ();
 sg13g2_fill_1 FILLER_68_1000 ();
 sg13g2_fill_1 FILLER_68_1005 ();
 sg13g2_fill_1 FILLER_68_1016 ();
 sg13g2_fill_2 FILLER_68_1037 ();
 sg13g2_fill_1 FILLER_68_1065 ();
 sg13g2_fill_1 FILLER_68_1110 ();
 sg13g2_decap_8 FILLER_68_1161 ();
 sg13g2_fill_2 FILLER_68_1168 ();
 sg13g2_fill_1 FILLER_68_1224 ();
 sg13g2_fill_2 FILLER_68_1251 ();
 sg13g2_decap_8 FILLER_68_1315 ();
 sg13g2_decap_8 FILLER_68_1322 ();
 sg13g2_decap_4 FILLER_68_1329 ();
 sg13g2_decap_8 FILLER_68_1336 ();
 sg13g2_decap_8 FILLER_68_1343 ();
 sg13g2_decap_4 FILLER_68_1350 ();
 sg13g2_fill_2 FILLER_68_1354 ();
 sg13g2_decap_4 FILLER_68_1405 ();
 sg13g2_fill_1 FILLER_68_1426 ();
 sg13g2_fill_1 FILLER_68_1431 ();
 sg13g2_fill_1 FILLER_68_1437 ();
 sg13g2_fill_2 FILLER_68_1464 ();
 sg13g2_fill_1 FILLER_68_1466 ();
 sg13g2_fill_2 FILLER_68_1471 ();
 sg13g2_fill_2 FILLER_68_1481 ();
 sg13g2_fill_1 FILLER_68_1483 ();
 sg13g2_fill_2 FILLER_68_1499 ();
 sg13g2_fill_1 FILLER_68_1501 ();
 sg13g2_fill_2 FILLER_68_1528 ();
 sg13g2_fill_1 FILLER_68_1530 ();
 sg13g2_decap_8 FILLER_68_1557 ();
 sg13g2_decap_4 FILLER_68_1570 ();
 sg13g2_fill_1 FILLER_68_1574 ();
 sg13g2_fill_2 FILLER_68_1594 ();
 sg13g2_fill_1 FILLER_68_1611 ();
 sg13g2_fill_2 FILLER_68_1620 ();
 sg13g2_fill_1 FILLER_68_1635 ();
 sg13g2_fill_1 FILLER_68_1704 ();
 sg13g2_fill_1 FILLER_68_1708 ();
 sg13g2_fill_1 FILLER_68_1715 ();
 sg13g2_fill_2 FILLER_68_1754 ();
 sg13g2_fill_1 FILLER_68_1756 ();
 sg13g2_fill_2 FILLER_68_1777 ();
 sg13g2_fill_2 FILLER_68_1796 ();
 sg13g2_fill_2 FILLER_68_1806 ();
 sg13g2_fill_1 FILLER_68_1808 ();
 sg13g2_fill_2 FILLER_68_1824 ();
 sg13g2_decap_4 FILLER_68_1858 ();
 sg13g2_decap_8 FILLER_68_1898 ();
 sg13g2_decap_8 FILLER_68_1941 ();
 sg13g2_decap_8 FILLER_68_1948 ();
 sg13g2_fill_2 FILLER_68_1955 ();
 sg13g2_decap_8 FILLER_68_1979 ();
 sg13g2_decap_8 FILLER_68_1986 ();
 sg13g2_decap_4 FILLER_68_1993 ();
 sg13g2_fill_1 FILLER_68_2005 ();
 sg13g2_fill_1 FILLER_68_2015 ();
 sg13g2_fill_1 FILLER_68_2020 ();
 sg13g2_decap_8 FILLER_68_2056 ();
 sg13g2_decap_4 FILLER_68_2063 ();
 sg13g2_fill_2 FILLER_68_2072 ();
 sg13g2_fill_2 FILLER_68_2087 ();
 sg13g2_fill_1 FILLER_68_2089 ();
 sg13g2_fill_2 FILLER_68_2097 ();
 sg13g2_fill_1 FILLER_68_2125 ();
 sg13g2_fill_1 FILLER_68_2150 ();
 sg13g2_fill_1 FILLER_68_2217 ();
 sg13g2_fill_1 FILLER_68_2247 ();
 sg13g2_fill_1 FILLER_68_2256 ();
 sg13g2_fill_2 FILLER_68_2263 ();
 sg13g2_decap_4 FILLER_68_2296 ();
 sg13g2_fill_1 FILLER_68_2300 ();
 sg13g2_decap_8 FILLER_68_2311 ();
 sg13g2_fill_2 FILLER_68_2355 ();
 sg13g2_fill_1 FILLER_68_2357 ();
 sg13g2_decap_8 FILLER_68_2405 ();
 sg13g2_fill_2 FILLER_68_2412 ();
 sg13g2_fill_2 FILLER_68_2453 ();
 sg13g2_fill_1 FILLER_68_2455 ();
 sg13g2_fill_2 FILLER_68_2504 ();
 sg13g2_decap_8 FILLER_68_2532 ();
 sg13g2_decap_8 FILLER_68_2539 ();
 sg13g2_decap_8 FILLER_68_2546 ();
 sg13g2_decap_8 FILLER_68_2553 ();
 sg13g2_decap_8 FILLER_68_2560 ();
 sg13g2_decap_8 FILLER_68_2567 ();
 sg13g2_decap_8 FILLER_68_2574 ();
 sg13g2_decap_8 FILLER_68_2581 ();
 sg13g2_decap_8 FILLER_68_2588 ();
 sg13g2_decap_8 FILLER_68_2595 ();
 sg13g2_decap_8 FILLER_68_2602 ();
 sg13g2_decap_8 FILLER_68_2609 ();
 sg13g2_decap_8 FILLER_68_2616 ();
 sg13g2_decap_8 FILLER_68_2623 ();
 sg13g2_decap_8 FILLER_68_2630 ();
 sg13g2_decap_8 FILLER_68_2637 ();
 sg13g2_decap_8 FILLER_68_2644 ();
 sg13g2_decap_8 FILLER_68_2651 ();
 sg13g2_decap_8 FILLER_68_2658 ();
 sg13g2_decap_4 FILLER_68_2665 ();
 sg13g2_fill_1 FILLER_68_2669 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_11 ();
 sg13g2_fill_2 FILLER_69_39 ();
 sg13g2_fill_1 FILLER_69_41 ();
 sg13g2_fill_2 FILLER_69_56 ();
 sg13g2_decap_4 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_91 ();
 sg13g2_fill_1 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_114 ();
 sg13g2_fill_1 FILLER_69_122 ();
 sg13g2_fill_2 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_137 ();
 sg13g2_decap_8 FILLER_69_141 ();
 sg13g2_fill_2 FILLER_69_148 ();
 sg13g2_fill_1 FILLER_69_150 ();
 sg13g2_fill_1 FILLER_69_155 ();
 sg13g2_fill_2 FILLER_69_161 ();
 sg13g2_fill_1 FILLER_69_173 ();
 sg13g2_fill_2 FILLER_69_184 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_fill_2 FILLER_69_207 ();
 sg13g2_decap_8 FILLER_69_214 ();
 sg13g2_decap_4 FILLER_69_221 ();
 sg13g2_decap_8 FILLER_69_230 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_276 ();
 sg13g2_decap_8 FILLER_69_284 ();
 sg13g2_fill_2 FILLER_69_291 ();
 sg13g2_fill_1 FILLER_69_366 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_fill_2 FILLER_69_387 ();
 sg13g2_fill_1 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_69_433 ();
 sg13g2_fill_1 FILLER_69_440 ();
 sg13g2_decap_8 FILLER_69_446 ();
 sg13g2_decap_8 FILLER_69_453 ();
 sg13g2_decap_8 FILLER_69_460 ();
 sg13g2_decap_8 FILLER_69_467 ();
 sg13g2_decap_8 FILLER_69_474 ();
 sg13g2_decap_4 FILLER_69_481 ();
 sg13g2_fill_1 FILLER_69_485 ();
 sg13g2_fill_2 FILLER_69_519 ();
 sg13g2_decap_8 FILLER_69_526 ();
 sg13g2_decap_8 FILLER_69_533 ();
 sg13g2_decap_4 FILLER_69_540 ();
 sg13g2_fill_2 FILLER_69_544 ();
 sg13g2_fill_2 FILLER_69_551 ();
 sg13g2_fill_2 FILLER_69_557 ();
 sg13g2_fill_2 FILLER_69_564 ();
 sg13g2_fill_1 FILLER_69_566 ();
 sg13g2_fill_1 FILLER_69_572 ();
 sg13g2_fill_2 FILLER_69_578 ();
 sg13g2_fill_1 FILLER_69_580 ();
 sg13g2_decap_8 FILLER_69_585 ();
 sg13g2_decap_8 FILLER_69_592 ();
 sg13g2_fill_1 FILLER_69_604 ();
 sg13g2_fill_1 FILLER_69_631 ();
 sg13g2_fill_2 FILLER_69_646 ();
 sg13g2_fill_1 FILLER_69_648 ();
 sg13g2_decap_4 FILLER_69_657 ();
 sg13g2_fill_2 FILLER_69_661 ();
 sg13g2_decap_4 FILLER_69_668 ();
 sg13g2_fill_1 FILLER_69_672 ();
 sg13g2_decap_8 FILLER_69_677 ();
 sg13g2_decap_8 FILLER_69_684 ();
 sg13g2_fill_1 FILLER_69_698 ();
 sg13g2_fill_1 FILLER_69_725 ();
 sg13g2_decap_4 FILLER_69_761 ();
 sg13g2_fill_2 FILLER_69_765 ();
 sg13g2_fill_2 FILLER_69_797 ();
 sg13g2_fill_1 FILLER_69_799 ();
 sg13g2_fill_1 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_4 FILLER_69_857 ();
 sg13g2_fill_2 FILLER_69_861 ();
 sg13g2_fill_2 FILLER_69_867 ();
 sg13g2_fill_1 FILLER_69_869 ();
 sg13g2_decap_4 FILLER_69_914 ();
 sg13g2_fill_2 FILLER_69_918 ();
 sg13g2_decap_8 FILLER_69_945 ();
 sg13g2_fill_2 FILLER_69_952 ();
 sg13g2_fill_1 FILLER_69_954 ();
 sg13g2_decap_4 FILLER_69_961 ();
 sg13g2_fill_2 FILLER_69_965 ();
 sg13g2_decap_8 FILLER_69_988 ();
 sg13g2_fill_1 FILLER_69_995 ();
 sg13g2_fill_1 FILLER_69_1008 ();
 sg13g2_fill_2 FILLER_69_1015 ();
 sg13g2_fill_1 FILLER_69_1071 ();
 sg13g2_fill_1 FILLER_69_1081 ();
 sg13g2_fill_2 FILLER_69_1092 ();
 sg13g2_decap_8 FILLER_69_1115 ();
 sg13g2_decap_8 FILLER_69_1122 ();
 sg13g2_decap_4 FILLER_69_1129 ();
 sg13g2_fill_1 FILLER_69_1137 ();
 sg13g2_fill_2 FILLER_69_1168 ();
 sg13g2_decap_8 FILLER_69_1176 ();
 sg13g2_decap_4 FILLER_69_1183 ();
 sg13g2_fill_2 FILLER_69_1187 ();
 sg13g2_fill_1 FILLER_69_1211 ();
 sg13g2_fill_1 FILLER_69_1227 ();
 sg13g2_decap_8 FILLER_69_1233 ();
 sg13g2_decap_4 FILLER_69_1240 ();
 sg13g2_fill_2 FILLER_69_1263 ();
 sg13g2_decap_4 FILLER_69_1269 ();
 sg13g2_fill_1 FILLER_69_1297 ();
 sg13g2_fill_2 FILLER_69_1304 ();
 sg13g2_fill_1 FILLER_69_1332 ();
 sg13g2_decap_8 FILLER_69_1410 ();
 sg13g2_fill_2 FILLER_69_1417 ();
 sg13g2_fill_2 FILLER_69_1427 ();
 sg13g2_fill_1 FILLER_69_1429 ();
 sg13g2_fill_2 FILLER_69_1463 ();
 sg13g2_decap_8 FILLER_69_1470 ();
 sg13g2_decap_8 FILLER_69_1477 ();
 sg13g2_fill_2 FILLER_69_1484 ();
 sg13g2_fill_1 FILLER_69_1486 ();
 sg13g2_decap_8 FILLER_69_1490 ();
 sg13g2_fill_2 FILLER_69_1510 ();
 sg13g2_decap_4 FILLER_69_1552 ();
 sg13g2_fill_1 FILLER_69_1584 ();
 sg13g2_fill_1 FILLER_69_1597 ();
 sg13g2_fill_2 FILLER_69_1627 ();
 sg13g2_decap_4 FILLER_69_1638 ();
 sg13g2_fill_2 FILLER_69_1642 ();
 sg13g2_fill_2 FILLER_69_1650 ();
 sg13g2_fill_1 FILLER_69_1652 ();
 sg13g2_decap_4 FILLER_69_1671 ();
 sg13g2_fill_1 FILLER_69_1675 ();
 sg13g2_fill_1 FILLER_69_1724 ();
 sg13g2_decap_8 FILLER_69_1747 ();
 sg13g2_decap_8 FILLER_69_1754 ();
 sg13g2_decap_4 FILLER_69_1761 ();
 sg13g2_fill_2 FILLER_69_1765 ();
 sg13g2_fill_2 FILLER_69_1771 ();
 sg13g2_fill_2 FILLER_69_1808 ();
 sg13g2_fill_1 FILLER_69_1810 ();
 sg13g2_fill_1 FILLER_69_1817 ();
 sg13g2_fill_2 FILLER_69_1831 ();
 sg13g2_fill_1 FILLER_69_1836 ();
 sg13g2_fill_2 FILLER_69_1890 ();
 sg13g2_fill_1 FILLER_69_1901 ();
 sg13g2_fill_1 FILLER_69_1908 ();
 sg13g2_decap_8 FILLER_69_1920 ();
 sg13g2_decap_4 FILLER_69_1927 ();
 sg13g2_fill_1 FILLER_69_1931 ();
 sg13g2_fill_2 FILLER_69_1941 ();
 sg13g2_fill_1 FILLER_69_1948 ();
 sg13g2_fill_1 FILLER_69_1953 ();
 sg13g2_decap_8 FILLER_69_1960 ();
 sg13g2_decap_8 FILLER_69_1967 ();
 sg13g2_decap_8 FILLER_69_1974 ();
 sg13g2_decap_8 FILLER_69_2026 ();
 sg13g2_fill_2 FILLER_69_2033 ();
 sg13g2_fill_1 FILLER_69_2035 ();
 sg13g2_decap_8 FILLER_69_2041 ();
 sg13g2_decap_8 FILLER_69_2048 ();
 sg13g2_decap_8 FILLER_69_2055 ();
 sg13g2_decap_8 FILLER_69_2093 ();
 sg13g2_decap_8 FILLER_69_2100 ();
 sg13g2_decap_4 FILLER_69_2107 ();
 sg13g2_fill_1 FILLER_69_2114 ();
 sg13g2_fill_1 FILLER_69_2124 ();
 sg13g2_fill_2 FILLER_69_2133 ();
 sg13g2_fill_1 FILLER_69_2140 ();
 sg13g2_decap_8 FILLER_69_2159 ();
 sg13g2_fill_1 FILLER_69_2166 ();
 sg13g2_fill_1 FILLER_69_2172 ();
 sg13g2_decap_8 FILLER_69_2177 ();
 sg13g2_fill_1 FILLER_69_2184 ();
 sg13g2_fill_1 FILLER_69_2209 ();
 sg13g2_fill_1 FILLER_69_2221 ();
 sg13g2_decap_8 FILLER_69_2282 ();
 sg13g2_decap_4 FILLER_69_2289 ();
 sg13g2_fill_1 FILLER_69_2293 ();
 sg13g2_decap_4 FILLER_69_2331 ();
 sg13g2_fill_1 FILLER_69_2340 ();
 sg13g2_decap_4 FILLER_69_2346 ();
 sg13g2_fill_1 FILLER_69_2350 ();
 sg13g2_fill_1 FILLER_69_2364 ();
 sg13g2_fill_1 FILLER_69_2375 ();
 sg13g2_decap_8 FILLER_69_2405 ();
 sg13g2_decap_8 FILLER_69_2412 ();
 sg13g2_decap_4 FILLER_69_2419 ();
 sg13g2_fill_2 FILLER_69_2423 ();
 sg13g2_fill_1 FILLER_69_2501 ();
 sg13g2_decap_8 FILLER_69_2506 ();
 sg13g2_decap_8 FILLER_69_2517 ();
 sg13g2_decap_8 FILLER_69_2524 ();
 sg13g2_decap_8 FILLER_69_2531 ();
 sg13g2_decap_8 FILLER_69_2538 ();
 sg13g2_decap_8 FILLER_69_2545 ();
 sg13g2_decap_8 FILLER_69_2552 ();
 sg13g2_decap_8 FILLER_69_2559 ();
 sg13g2_decap_8 FILLER_69_2566 ();
 sg13g2_decap_8 FILLER_69_2573 ();
 sg13g2_decap_8 FILLER_69_2580 ();
 sg13g2_decap_8 FILLER_69_2587 ();
 sg13g2_decap_8 FILLER_69_2594 ();
 sg13g2_decap_8 FILLER_69_2601 ();
 sg13g2_decap_8 FILLER_69_2608 ();
 sg13g2_decap_8 FILLER_69_2615 ();
 sg13g2_decap_8 FILLER_69_2622 ();
 sg13g2_decap_8 FILLER_69_2629 ();
 sg13g2_decap_8 FILLER_69_2636 ();
 sg13g2_decap_8 FILLER_69_2643 ();
 sg13g2_decap_8 FILLER_69_2650 ();
 sg13g2_decap_8 FILLER_69_2657 ();
 sg13g2_decap_4 FILLER_69_2664 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_40 ();
 sg13g2_decap_4 FILLER_70_57 ();
 sg13g2_fill_2 FILLER_70_61 ();
 sg13g2_fill_2 FILLER_70_79 ();
 sg13g2_fill_1 FILLER_70_81 ();
 sg13g2_fill_2 FILLER_70_90 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_decap_4 FILLER_70_116 ();
 sg13g2_fill_1 FILLER_70_120 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_132 ();
 sg13g2_fill_1 FILLER_70_134 ();
 sg13g2_fill_2 FILLER_70_144 ();
 sg13g2_fill_1 FILLER_70_166 ();
 sg13g2_fill_1 FILLER_70_172 ();
 sg13g2_fill_1 FILLER_70_183 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_196 ();
 sg13g2_decap_4 FILLER_70_211 ();
 sg13g2_decap_8 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_230 ();
 sg13g2_fill_1 FILLER_70_236 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_270 ();
 sg13g2_decap_4 FILLER_70_293 ();
 sg13g2_fill_2 FILLER_70_302 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_fill_1 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_351 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_fill_2 FILLER_70_375 ();
 sg13g2_fill_1 FILLER_70_405 ();
 sg13g2_fill_1 FILLER_70_410 ();
 sg13g2_fill_1 FILLER_70_421 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_fill_1 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_439 ();
 sg13g2_decap_8 FILLER_70_446 ();
 sg13g2_decap_4 FILLER_70_453 ();
 sg13g2_fill_2 FILLER_70_457 ();
 sg13g2_fill_1 FILLER_70_464 ();
 sg13g2_fill_2 FILLER_70_469 ();
 sg13g2_fill_1 FILLER_70_497 ();
 sg13g2_fill_1 FILLER_70_514 ();
 sg13g2_fill_1 FILLER_70_521 ();
 sg13g2_decap_8 FILLER_70_536 ();
 sg13g2_fill_1 FILLER_70_543 ();
 sg13g2_fill_1 FILLER_70_576 ();
 sg13g2_fill_2 FILLER_70_650 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_decap_4 FILLER_70_674 ();
 sg13g2_fill_2 FILLER_70_678 ();
 sg13g2_decap_4 FILLER_70_684 ();
 sg13g2_fill_2 FILLER_70_722 ();
 sg13g2_fill_1 FILLER_70_724 ();
 sg13g2_decap_8 FILLER_70_745 ();
 sg13g2_decap_8 FILLER_70_752 ();
 sg13g2_decap_8 FILLER_70_759 ();
 sg13g2_decap_8 FILLER_70_766 ();
 sg13g2_decap_8 FILLER_70_773 ();
 sg13g2_decap_8 FILLER_70_780 ();
 sg13g2_decap_8 FILLER_70_787 ();
 sg13g2_fill_1 FILLER_70_794 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_decap_4 FILLER_70_845 ();
 sg13g2_fill_1 FILLER_70_849 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_decap_4 FILLER_70_871 ();
 sg13g2_fill_2 FILLER_70_894 ();
 sg13g2_fill_2 FILLER_70_901 ();
 sg13g2_fill_2 FILLER_70_929 ();
 sg13g2_decap_8 FILLER_70_957 ();
 sg13g2_decap_8 FILLER_70_964 ();
 sg13g2_fill_1 FILLER_70_971 ();
 sg13g2_fill_2 FILLER_70_1037 ();
 sg13g2_fill_1 FILLER_70_1096 ();
 sg13g2_decap_8 FILLER_70_1112 ();
 sg13g2_decap_8 FILLER_70_1119 ();
 sg13g2_decap_4 FILLER_70_1126 ();
 sg13g2_fill_2 FILLER_70_1130 ();
 sg13g2_fill_2 FILLER_70_1137 ();
 sg13g2_decap_8 FILLER_70_1185 ();
 sg13g2_fill_2 FILLER_70_1192 ();
 sg13g2_decap_4 FILLER_70_1228 ();
 sg13g2_decap_8 FILLER_70_1258 ();
 sg13g2_fill_2 FILLER_70_1270 ();
 sg13g2_fill_1 FILLER_70_1272 ();
 sg13g2_fill_1 FILLER_70_1281 ();
 sg13g2_decap_8 FILLER_70_1288 ();
 sg13g2_fill_1 FILLER_70_1295 ();
 sg13g2_decap_8 FILLER_70_1302 ();
 sg13g2_decap_4 FILLER_70_1309 ();
 sg13g2_fill_2 FILLER_70_1317 ();
 sg13g2_fill_1 FILLER_70_1319 ();
 sg13g2_fill_1 FILLER_70_1329 ();
 sg13g2_decap_8 FILLER_70_1348 ();
 sg13g2_fill_2 FILLER_70_1355 ();
 sg13g2_fill_2 FILLER_70_1373 ();
 sg13g2_decap_8 FILLER_70_1400 ();
 sg13g2_decap_8 FILLER_70_1412 ();
 sg13g2_decap_8 FILLER_70_1419 ();
 sg13g2_decap_8 FILLER_70_1426 ();
 sg13g2_decap_4 FILLER_70_1433 ();
 sg13g2_fill_2 FILLER_70_1466 ();
 sg13g2_fill_1 FILLER_70_1468 ();
 sg13g2_fill_1 FILLER_70_1503 ();
 sg13g2_fill_1 FILLER_70_1524 ();
 sg13g2_decap_8 FILLER_70_1602 ();
 sg13g2_decap_8 FILLER_70_1609 ();
 sg13g2_decap_8 FILLER_70_1616 ();
 sg13g2_decap_4 FILLER_70_1623 ();
 sg13g2_fill_2 FILLER_70_1627 ();
 sg13g2_fill_2 FILLER_70_1638 ();
 sg13g2_fill_2 FILLER_70_1650 ();
 sg13g2_fill_1 FILLER_70_1652 ();
 sg13g2_fill_1 FILLER_70_1665 ();
 sg13g2_fill_1 FILLER_70_1676 ();
 sg13g2_fill_1 FILLER_70_1737 ();
 sg13g2_decap_8 FILLER_70_1747 ();
 sg13g2_decap_8 FILLER_70_1754 ();
 sg13g2_decap_8 FILLER_70_1761 ();
 sg13g2_fill_1 FILLER_70_1768 ();
 sg13g2_fill_1 FILLER_70_1794 ();
 sg13g2_decap_4 FILLER_70_1869 ();
 sg13g2_fill_2 FILLER_70_1881 ();
 sg13g2_fill_1 FILLER_70_1883 ();
 sg13g2_fill_1 FILLER_70_1893 ();
 sg13g2_fill_1 FILLER_70_1942 ();
 sg13g2_fill_2 FILLER_70_1969 ();
 sg13g2_decap_4 FILLER_70_1976 ();
 sg13g2_fill_1 FILLER_70_1980 ();
 sg13g2_fill_2 FILLER_70_1985 ();
 sg13g2_fill_1 FILLER_70_1987 ();
 sg13g2_decap_8 FILLER_70_1991 ();
 sg13g2_decap_8 FILLER_70_1998 ();
 sg13g2_decap_8 FILLER_70_2005 ();
 sg13g2_fill_1 FILLER_70_2012 ();
 sg13g2_decap_8 FILLER_70_2016 ();
 sg13g2_decap_4 FILLER_70_2023 ();
 sg13g2_decap_8 FILLER_70_2063 ();
 sg13g2_decap_8 FILLER_70_2070 ();
 sg13g2_decap_4 FILLER_70_2077 ();
 sg13g2_fill_2 FILLER_70_2081 ();
 sg13g2_decap_8 FILLER_70_2096 ();
 sg13g2_decap_4 FILLER_70_2103 ();
 sg13g2_fill_1 FILLER_70_2107 ();
 sg13g2_fill_1 FILLER_70_2117 ();
 sg13g2_fill_1 FILLER_70_2198 ();
 sg13g2_fill_2 FILLER_70_2211 ();
 sg13g2_fill_2 FILLER_70_2252 ();
 sg13g2_decap_4 FILLER_70_2299 ();
 sg13g2_fill_1 FILLER_70_2303 ();
 sg13g2_fill_2 FILLER_70_2312 ();
 sg13g2_fill_2 FILLER_70_2379 ();
 sg13g2_decap_8 FILLER_70_2394 ();
 sg13g2_decap_8 FILLER_70_2401 ();
 sg13g2_decap_8 FILLER_70_2408 ();
 sg13g2_decap_8 FILLER_70_2415 ();
 sg13g2_decap_8 FILLER_70_2422 ();
 sg13g2_fill_2 FILLER_70_2429 ();
 sg13g2_decap_4 FILLER_70_2435 ();
 sg13g2_fill_1 FILLER_70_2439 ();
 sg13g2_fill_1 FILLER_70_2444 ();
 sg13g2_decap_8 FILLER_70_2501 ();
 sg13g2_decap_8 FILLER_70_2508 ();
 sg13g2_decap_8 FILLER_70_2515 ();
 sg13g2_decap_8 FILLER_70_2522 ();
 sg13g2_decap_8 FILLER_70_2529 ();
 sg13g2_decap_8 FILLER_70_2536 ();
 sg13g2_decap_8 FILLER_70_2543 ();
 sg13g2_decap_8 FILLER_70_2550 ();
 sg13g2_decap_8 FILLER_70_2557 ();
 sg13g2_decap_8 FILLER_70_2564 ();
 sg13g2_decap_8 FILLER_70_2571 ();
 sg13g2_decap_8 FILLER_70_2578 ();
 sg13g2_decap_8 FILLER_70_2585 ();
 sg13g2_decap_8 FILLER_70_2592 ();
 sg13g2_decap_8 FILLER_70_2599 ();
 sg13g2_decap_8 FILLER_70_2606 ();
 sg13g2_decap_8 FILLER_70_2613 ();
 sg13g2_decap_8 FILLER_70_2620 ();
 sg13g2_decap_8 FILLER_70_2627 ();
 sg13g2_decap_8 FILLER_70_2634 ();
 sg13g2_decap_8 FILLER_70_2641 ();
 sg13g2_decap_8 FILLER_70_2648 ();
 sg13g2_decap_8 FILLER_70_2655 ();
 sg13g2_decap_8 FILLER_70_2662 ();
 sg13g2_fill_1 FILLER_70_2669 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_4 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_22 ();
 sg13g2_decap_4 FILLER_71_36 ();
 sg13g2_fill_2 FILLER_71_40 ();
 sg13g2_decap_4 FILLER_71_46 ();
 sg13g2_fill_2 FILLER_71_50 ();
 sg13g2_decap_4 FILLER_71_58 ();
 sg13g2_fill_1 FILLER_71_62 ();
 sg13g2_fill_1 FILLER_71_74 ();
 sg13g2_fill_1 FILLER_71_88 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_131 ();
 sg13g2_fill_2 FILLER_71_136 ();
 sg13g2_fill_2 FILLER_71_156 ();
 sg13g2_fill_1 FILLER_71_163 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_175 ();
 sg13g2_fill_2 FILLER_71_186 ();
 sg13g2_fill_1 FILLER_71_188 ();
 sg13g2_fill_2 FILLER_71_194 ();
 sg13g2_fill_2 FILLER_71_201 ();
 sg13g2_fill_2 FILLER_71_213 ();
 sg13g2_fill_1 FILLER_71_219 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_fill_2 FILLER_71_231 ();
 sg13g2_fill_1 FILLER_71_242 ();
 sg13g2_fill_1 FILLER_71_247 ();
 sg13g2_fill_1 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_267 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_decap_4 FILLER_71_325 ();
 sg13g2_fill_2 FILLER_71_329 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_fill_1 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_388 ();
 sg13g2_fill_2 FILLER_71_395 ();
 sg13g2_fill_1 FILLER_71_397 ();
 sg13g2_fill_1 FILLER_71_417 ();
 sg13g2_decap_4 FILLER_71_428 ();
 sg13g2_decap_4 FILLER_71_441 ();
 sg13g2_fill_2 FILLER_71_445 ();
 sg13g2_decap_8 FILLER_71_452 ();
 sg13g2_decap_8 FILLER_71_459 ();
 sg13g2_fill_2 FILLER_71_466 ();
 sg13g2_fill_1 FILLER_71_468 ();
 sg13g2_decap_4 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_506 ();
 sg13g2_fill_2 FILLER_71_522 ();
 sg13g2_decap_8 FILLER_71_532 ();
 sg13g2_decap_8 FILLER_71_539 ();
 sg13g2_decap_4 FILLER_71_546 ();
 sg13g2_fill_1 FILLER_71_550 ();
 sg13g2_decap_4 FILLER_71_555 ();
 sg13g2_decap_4 FILLER_71_563 ();
 sg13g2_fill_1 FILLER_71_567 ();
 sg13g2_fill_1 FILLER_71_572 ();
 sg13g2_decap_8 FILLER_71_578 ();
 sg13g2_decap_8 FILLER_71_585 ();
 sg13g2_fill_1 FILLER_71_592 ();
 sg13g2_decap_8 FILLER_71_597 ();
 sg13g2_decap_8 FILLER_71_604 ();
 sg13g2_fill_2 FILLER_71_611 ();
 sg13g2_fill_1 FILLER_71_613 ();
 sg13g2_decap_8 FILLER_71_635 ();
 sg13g2_decap_8 FILLER_71_642 ();
 sg13g2_decap_8 FILLER_71_649 ();
 sg13g2_decap_4 FILLER_71_656 ();
 sg13g2_decap_8 FILLER_71_670 ();
 sg13g2_decap_4 FILLER_71_677 ();
 sg13g2_fill_1 FILLER_71_681 ();
 sg13g2_decap_4 FILLER_71_695 ();
 sg13g2_fill_2 FILLER_71_699 ();
 sg13g2_fill_2 FILLER_71_735 ();
 sg13g2_decap_8 FILLER_71_741 ();
 sg13g2_decap_8 FILLER_71_748 ();
 sg13g2_fill_2 FILLER_71_759 ();
 sg13g2_fill_2 FILLER_71_765 ();
 sg13g2_fill_1 FILLER_71_803 ();
 sg13g2_fill_2 FILLER_71_862 ();
 sg13g2_fill_1 FILLER_71_881 ();
 sg13g2_fill_2 FILLER_71_899 ();
 sg13g2_decap_4 FILLER_71_937 ();
 sg13g2_fill_2 FILLER_71_941 ();
 sg13g2_decap_8 FILLER_71_953 ();
 sg13g2_decap_4 FILLER_71_960 ();
 sg13g2_decap_4 FILLER_71_974 ();
 sg13g2_fill_1 FILLER_71_978 ();
 sg13g2_fill_2 FILLER_71_992 ();
 sg13g2_fill_1 FILLER_71_1050 ();
 sg13g2_fill_1 FILLER_71_1058 ();
 sg13g2_fill_1 FILLER_71_1068 ();
 sg13g2_fill_1 FILLER_71_1093 ();
 sg13g2_fill_1 FILLER_71_1110 ();
 sg13g2_decap_8 FILLER_71_1142 ();
 sg13g2_decap_8 FILLER_71_1149 ();
 sg13g2_decap_8 FILLER_71_1196 ();
 sg13g2_decap_4 FILLER_71_1203 ();
 sg13g2_fill_2 FILLER_71_1223 ();
 sg13g2_decap_8 FILLER_71_1251 ();
 sg13g2_decap_8 FILLER_71_1258 ();
 sg13g2_decap_8 FILLER_71_1265 ();
 sg13g2_decap_8 FILLER_71_1272 ();
 sg13g2_decap_8 FILLER_71_1279 ();
 sg13g2_decap_8 FILLER_71_1286 ();
 sg13g2_fill_1 FILLER_71_1293 ();
 sg13g2_fill_1 FILLER_71_1313 ();
 sg13g2_fill_2 FILLER_71_1337 ();
 sg13g2_fill_1 FILLER_71_1339 ();
 sg13g2_decap_8 FILLER_71_1366 ();
 sg13g2_decap_8 FILLER_71_1373 ();
 sg13g2_decap_8 FILLER_71_1380 ();
 sg13g2_decap_8 FILLER_71_1387 ();
 sg13g2_decap_8 FILLER_71_1394 ();
 sg13g2_decap_4 FILLER_71_1401 ();
 sg13g2_fill_2 FILLER_71_1405 ();
 sg13g2_fill_1 FILLER_71_1468 ();
 sg13g2_fill_2 FILLER_71_1498 ();
 sg13g2_fill_1 FILLER_71_1527 ();
 sg13g2_fill_2 FILLER_71_1560 ();
 sg13g2_fill_1 FILLER_71_1562 ();
 sg13g2_decap_8 FILLER_71_1592 ();
 sg13g2_decap_8 FILLER_71_1599 ();
 sg13g2_fill_2 FILLER_71_1606 ();
 sg13g2_decap_8 FILLER_71_1614 ();
 sg13g2_decap_8 FILLER_71_1621 ();
 sg13g2_fill_1 FILLER_71_1682 ();
 sg13g2_fill_2 FILLER_71_1693 ();
 sg13g2_fill_2 FILLER_71_1734 ();
 sg13g2_fill_1 FILLER_71_1772 ();
 sg13g2_fill_1 FILLER_71_1787 ();
 sg13g2_fill_1 FILLER_71_1793 ();
 sg13g2_fill_1 FILLER_71_1799 ();
 sg13g2_fill_2 FILLER_71_1838 ();
 sg13g2_fill_2 FILLER_71_1843 ();
 sg13g2_fill_2 FILLER_71_1881 ();
 sg13g2_fill_2 FILLER_71_1916 ();
 sg13g2_fill_1 FILLER_71_1926 ();
 sg13g2_decap_8 FILLER_71_1999 ();
 sg13g2_fill_2 FILLER_71_2006 ();
 sg13g2_fill_1 FILLER_71_2008 ();
 sg13g2_decap_8 FILLER_71_2019 ();
 sg13g2_fill_1 FILLER_71_2026 ();
 sg13g2_fill_1 FILLER_71_2036 ();
 sg13g2_decap_4 FILLER_71_2063 ();
 sg13g2_fill_2 FILLER_71_2067 ();
 sg13g2_decap_4 FILLER_71_2107 ();
 sg13g2_decap_8 FILLER_71_2119 ();
 sg13g2_decap_4 FILLER_71_2126 ();
 sg13g2_fill_1 FILLER_71_2139 ();
 sg13g2_fill_2 FILLER_71_2183 ();
 sg13g2_fill_1 FILLER_71_2185 ();
 sg13g2_fill_2 FILLER_71_2211 ();
 sg13g2_fill_1 FILLER_71_2251 ();
 sg13g2_decap_4 FILLER_71_2267 ();
 sg13g2_fill_1 FILLER_71_2271 ();
 sg13g2_decap_4 FILLER_71_2285 ();
 sg13g2_fill_1 FILLER_71_2289 ();
 sg13g2_decap_4 FILLER_71_2301 ();
 sg13g2_decap_8 FILLER_71_2310 ();
 sg13g2_decap_8 FILLER_71_2317 ();
 sg13g2_decap_8 FILLER_71_2329 ();
 sg13g2_decap_8 FILLER_71_2336 ();
 sg13g2_decap_8 FILLER_71_2343 ();
 sg13g2_decap_8 FILLER_71_2350 ();
 sg13g2_decap_8 FILLER_71_2391 ();
 sg13g2_decap_8 FILLER_71_2398 ();
 sg13g2_fill_1 FILLER_71_2405 ();
 sg13g2_decap_4 FILLER_71_2450 ();
 sg13g2_decap_8 FILLER_71_2458 ();
 sg13g2_decap_8 FILLER_71_2465 ();
 sg13g2_decap_8 FILLER_71_2472 ();
 sg13g2_decap_8 FILLER_71_2491 ();
 sg13g2_decap_8 FILLER_71_2498 ();
 sg13g2_decap_8 FILLER_71_2505 ();
 sg13g2_decap_8 FILLER_71_2512 ();
 sg13g2_decap_8 FILLER_71_2519 ();
 sg13g2_decap_8 FILLER_71_2526 ();
 sg13g2_decap_8 FILLER_71_2533 ();
 sg13g2_decap_8 FILLER_71_2540 ();
 sg13g2_decap_8 FILLER_71_2547 ();
 sg13g2_decap_8 FILLER_71_2554 ();
 sg13g2_decap_8 FILLER_71_2561 ();
 sg13g2_decap_8 FILLER_71_2568 ();
 sg13g2_decap_8 FILLER_71_2575 ();
 sg13g2_decap_8 FILLER_71_2582 ();
 sg13g2_decap_8 FILLER_71_2589 ();
 sg13g2_decap_8 FILLER_71_2596 ();
 sg13g2_decap_8 FILLER_71_2603 ();
 sg13g2_decap_8 FILLER_71_2610 ();
 sg13g2_decap_8 FILLER_71_2617 ();
 sg13g2_decap_8 FILLER_71_2624 ();
 sg13g2_decap_8 FILLER_71_2631 ();
 sg13g2_decap_8 FILLER_71_2638 ();
 sg13g2_decap_8 FILLER_71_2645 ();
 sg13g2_decap_8 FILLER_71_2652 ();
 sg13g2_decap_8 FILLER_71_2659 ();
 sg13g2_decap_4 FILLER_71_2666 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_9 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_43 ();
 sg13g2_decap_4 FILLER_72_55 ();
 sg13g2_fill_1 FILLER_72_63 ();
 sg13g2_decap_4 FILLER_72_68 ();
 sg13g2_fill_2 FILLER_72_96 ();
 sg13g2_fill_1 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_129 ();
 sg13g2_fill_2 FILLER_72_151 ();
 sg13g2_fill_1 FILLER_72_153 ();
 sg13g2_fill_2 FILLER_72_169 ();
 sg13g2_fill_2 FILLER_72_175 ();
 sg13g2_fill_2 FILLER_72_181 ();
 sg13g2_fill_1 FILLER_72_193 ();
 sg13g2_fill_2 FILLER_72_198 ();
 sg13g2_fill_1 FILLER_72_200 ();
 sg13g2_decap_4 FILLER_72_207 ();
 sg13g2_decap_8 FILLER_72_215 ();
 sg13g2_fill_1 FILLER_72_222 ();
 sg13g2_decap_8 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_260 ();
 sg13g2_fill_2 FILLER_72_269 ();
 sg13g2_fill_1 FILLER_72_275 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_fill_2 FILLER_72_290 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_fill_1 FILLER_72_300 ();
 sg13g2_fill_2 FILLER_72_305 ();
 sg13g2_fill_2 FILLER_72_342 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_fill_2 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_390 ();
 sg13g2_decap_8 FILLER_72_397 ();
 sg13g2_decap_8 FILLER_72_409 ();
 sg13g2_fill_2 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_429 ();
 sg13g2_decap_4 FILLER_72_436 ();
 sg13g2_fill_1 FILLER_72_466 ();
 sg13g2_fill_2 FILLER_72_472 ();
 sg13g2_fill_1 FILLER_72_474 ();
 sg13g2_fill_1 FILLER_72_542 ();
 sg13g2_decap_4 FILLER_72_547 ();
 sg13g2_decap_4 FILLER_72_561 ();
 sg13g2_decap_4 FILLER_72_570 ();
 sg13g2_fill_2 FILLER_72_578 ();
 sg13g2_fill_1 FILLER_72_580 ();
 sg13g2_decap_8 FILLER_72_584 ();
 sg13g2_fill_2 FILLER_72_591 ();
 sg13g2_decap_4 FILLER_72_598 ();
 sg13g2_fill_1 FILLER_72_602 ();
 sg13g2_fill_2 FILLER_72_607 ();
 sg13g2_fill_1 FILLER_72_617 ();
 sg13g2_decap_8 FILLER_72_627 ();
 sg13g2_decap_8 FILLER_72_634 ();
 sg13g2_fill_2 FILLER_72_641 ();
 sg13g2_decap_8 FILLER_72_647 ();
 sg13g2_decap_8 FILLER_72_654 ();
 sg13g2_fill_1 FILLER_72_661 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_8 FILLER_72_679 ();
 sg13g2_decap_8 FILLER_72_686 ();
 sg13g2_decap_4 FILLER_72_693 ();
 sg13g2_decap_4 FILLER_72_702 ();
 sg13g2_fill_1 FILLER_72_706 ();
 sg13g2_decap_4 FILLER_72_720 ();
 sg13g2_decap_4 FILLER_72_737 ();
 sg13g2_fill_2 FILLER_72_741 ();
 sg13g2_fill_2 FILLER_72_773 ();
 sg13g2_fill_1 FILLER_72_775 ();
 sg13g2_decap_4 FILLER_72_782 ();
 sg13g2_fill_2 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_fill_2 FILLER_72_799 ();
 sg13g2_fill_2 FILLER_72_820 ();
 sg13g2_fill_1 FILLER_72_827 ();
 sg13g2_fill_1 FILLER_72_850 ();
 sg13g2_fill_2 FILLER_72_877 ();
 sg13g2_fill_1 FILLER_72_890 ();
 sg13g2_decap_8 FILLER_72_910 ();
 sg13g2_decap_8 FILLER_72_917 ();
 sg13g2_decap_8 FILLER_72_924 ();
 sg13g2_fill_2 FILLER_72_931 ();
 sg13g2_fill_1 FILLER_72_933 ();
 sg13g2_fill_2 FILLER_72_948 ();
 sg13g2_decap_4 FILLER_72_968 ();
 sg13g2_fill_1 FILLER_72_976 ();
 sg13g2_fill_2 FILLER_72_995 ();
 sg13g2_fill_1 FILLER_72_1008 ();
 sg13g2_fill_1 FILLER_72_1022 ();
 sg13g2_fill_2 FILLER_72_1069 ();
 sg13g2_fill_1 FILLER_72_1075 ();
 sg13g2_fill_2 FILLER_72_1080 ();
 sg13g2_fill_2 FILLER_72_1095 ();
 sg13g2_decap_8 FILLER_72_1180 ();
 sg13g2_decap_8 FILLER_72_1187 ();
 sg13g2_decap_8 FILLER_72_1194 ();
 sg13g2_decap_4 FILLER_72_1201 ();
 sg13g2_fill_1 FILLER_72_1205 ();
 sg13g2_fill_2 FILLER_72_1210 ();
 sg13g2_fill_1 FILLER_72_1212 ();
 sg13g2_decap_8 FILLER_72_1224 ();
 sg13g2_decap_8 FILLER_72_1231 ();
 sg13g2_decap_4 FILLER_72_1238 ();
 sg13g2_fill_1 FILLER_72_1272 ();
 sg13g2_fill_1 FILLER_72_1277 ();
 sg13g2_fill_2 FILLER_72_1304 ();
 sg13g2_fill_1 FILLER_72_1345 ();
 sg13g2_fill_2 FILLER_72_1364 ();
 sg13g2_fill_2 FILLER_72_1370 ();
 sg13g2_fill_1 FILLER_72_1372 ();
 sg13g2_decap_8 FILLER_72_1377 ();
 sg13g2_decap_8 FILLER_72_1384 ();
 sg13g2_fill_2 FILLER_72_1391 ();
 sg13g2_decap_8 FILLER_72_1414 ();
 sg13g2_decap_8 FILLER_72_1421 ();
 sg13g2_decap_8 FILLER_72_1428 ();
 sg13g2_decap_8 FILLER_72_1435 ();
 sg13g2_decap_8 FILLER_72_1442 ();
 sg13g2_fill_2 FILLER_72_1449 ();
 sg13g2_fill_2 FILLER_72_1487 ();
 sg13g2_fill_2 FILLER_72_1503 ();
 sg13g2_decap_4 FILLER_72_1572 ();
 sg13g2_decap_4 FILLER_72_1585 ();
 sg13g2_decap_8 FILLER_72_1595 ();
 sg13g2_fill_2 FILLER_72_1644 ();
 sg13g2_decap_8 FILLER_72_1685 ();
 sg13g2_fill_2 FILLER_72_1692 ();
 sg13g2_fill_1 FILLER_72_1825 ();
 sg13g2_fill_2 FILLER_72_1835 ();
 sg13g2_fill_1 FILLER_72_1855 ();
 sg13g2_fill_1 FILLER_72_1882 ();
 sg13g2_fill_1 FILLER_72_1888 ();
 sg13g2_fill_1 FILLER_72_1918 ();
 sg13g2_decap_4 FILLER_72_1971 ();
 sg13g2_fill_2 FILLER_72_1975 ();
 sg13g2_decap_4 FILLER_72_1991 ();
 sg13g2_decap_8 FILLER_72_2053 ();
 sg13g2_fill_2 FILLER_72_2060 ();
 sg13g2_decap_4 FILLER_72_2096 ();
 sg13g2_fill_1 FILLER_72_2100 ();
 sg13g2_fill_2 FILLER_72_2110 ();
 sg13g2_fill_1 FILLER_72_2112 ();
 sg13g2_decap_4 FILLER_72_2121 ();
 sg13g2_fill_1 FILLER_72_2125 ();
 sg13g2_decap_4 FILLER_72_2178 ();
 sg13g2_fill_1 FILLER_72_2182 ();
 sg13g2_fill_1 FILLER_72_2209 ();
 sg13g2_fill_1 FILLER_72_2232 ();
 sg13g2_fill_2 FILLER_72_2245 ();
 sg13g2_fill_1 FILLER_72_2247 ();
 sg13g2_fill_2 FILLER_72_2251 ();
 sg13g2_fill_1 FILLER_72_2253 ();
 sg13g2_fill_2 FILLER_72_2312 ();
 sg13g2_fill_2 FILLER_72_2319 ();
 sg13g2_fill_2 FILLER_72_2382 ();
 sg13g2_decap_4 FILLER_72_2405 ();
 sg13g2_fill_2 FILLER_72_2439 ();
 sg13g2_decap_8 FILLER_72_2445 ();
 sg13g2_decap_8 FILLER_72_2452 ();
 sg13g2_decap_8 FILLER_72_2459 ();
 sg13g2_decap_8 FILLER_72_2466 ();
 sg13g2_decap_8 FILLER_72_2473 ();
 sg13g2_decap_8 FILLER_72_2480 ();
 sg13g2_decap_8 FILLER_72_2487 ();
 sg13g2_decap_8 FILLER_72_2494 ();
 sg13g2_decap_8 FILLER_72_2501 ();
 sg13g2_decap_8 FILLER_72_2508 ();
 sg13g2_decap_8 FILLER_72_2515 ();
 sg13g2_decap_8 FILLER_72_2522 ();
 sg13g2_decap_8 FILLER_72_2529 ();
 sg13g2_decap_8 FILLER_72_2536 ();
 sg13g2_decap_8 FILLER_72_2543 ();
 sg13g2_decap_8 FILLER_72_2550 ();
 sg13g2_decap_8 FILLER_72_2557 ();
 sg13g2_decap_8 FILLER_72_2564 ();
 sg13g2_decap_8 FILLER_72_2571 ();
 sg13g2_decap_8 FILLER_72_2578 ();
 sg13g2_decap_8 FILLER_72_2585 ();
 sg13g2_decap_8 FILLER_72_2592 ();
 sg13g2_decap_8 FILLER_72_2599 ();
 sg13g2_decap_8 FILLER_72_2606 ();
 sg13g2_decap_8 FILLER_72_2613 ();
 sg13g2_decap_8 FILLER_72_2620 ();
 sg13g2_decap_8 FILLER_72_2627 ();
 sg13g2_decap_8 FILLER_72_2634 ();
 sg13g2_decap_8 FILLER_72_2641 ();
 sg13g2_decap_8 FILLER_72_2648 ();
 sg13g2_decap_8 FILLER_72_2655 ();
 sg13g2_decap_8 FILLER_72_2662 ();
 sg13g2_fill_1 FILLER_72_2669 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_9 ();
 sg13g2_fill_2 FILLER_73_30 ();
 sg13g2_fill_2 FILLER_73_52 ();
 sg13g2_decap_8 FILLER_73_60 ();
 sg13g2_decap_4 FILLER_73_67 ();
 sg13g2_fill_1 FILLER_73_71 ();
 sg13g2_fill_2 FILLER_73_76 ();
 sg13g2_fill_1 FILLER_73_82 ();
 sg13g2_fill_2 FILLER_73_88 ();
 sg13g2_fill_1 FILLER_73_90 ();
 sg13g2_fill_1 FILLER_73_152 ();
 sg13g2_decap_4 FILLER_73_164 ();
 sg13g2_decap_4 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_fill_2 FILLER_73_200 ();
 sg13g2_decap_8 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_216 ();
 sg13g2_decap_8 FILLER_73_223 ();
 sg13g2_decap_8 FILLER_73_230 ();
 sg13g2_decap_8 FILLER_73_237 ();
 sg13g2_decap_8 FILLER_73_248 ();
 sg13g2_decap_4 FILLER_73_264 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_4 FILLER_73_328 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_decap_8 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_345 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_73_409 ();
 sg13g2_decap_4 FILLER_73_416 ();
 sg13g2_fill_2 FILLER_73_450 ();
 sg13g2_decap_8 FILLER_73_456 ();
 sg13g2_fill_2 FILLER_73_463 ();
 sg13g2_fill_1 FILLER_73_465 ();
 sg13g2_fill_1 FILLER_73_516 ();
 sg13g2_decap_8 FILLER_73_521 ();
 sg13g2_decap_4 FILLER_73_528 ();
 sg13g2_fill_1 FILLER_73_532 ();
 sg13g2_fill_2 FILLER_73_556 ();
 sg13g2_fill_2 FILLER_73_571 ();
 sg13g2_decap_4 FILLER_73_578 ();
 sg13g2_fill_2 FILLER_73_582 ();
 sg13g2_decap_8 FILLER_73_592 ();
 sg13g2_fill_1 FILLER_73_599 ();
 sg13g2_decap_8 FILLER_73_620 ();
 sg13g2_fill_2 FILLER_73_627 ();
 sg13g2_fill_1 FILLER_73_629 ();
 sg13g2_fill_1 FILLER_73_639 ();
 sg13g2_fill_1 FILLER_73_648 ();
 sg13g2_fill_2 FILLER_73_654 ();
 sg13g2_fill_2 FILLER_73_661 ();
 sg13g2_fill_1 FILLER_73_663 ();
 sg13g2_fill_1 FILLER_73_669 ();
 sg13g2_decap_8 FILLER_73_675 ();
 sg13g2_decap_4 FILLER_73_682 ();
 sg13g2_fill_1 FILLER_73_698 ();
 sg13g2_decap_8 FILLER_73_734 ();
 sg13g2_fill_2 FILLER_73_741 ();
 sg13g2_fill_1 FILLER_73_743 ();
 sg13g2_fill_2 FILLER_73_748 ();
 sg13g2_fill_1 FILLER_73_750 ();
 sg13g2_decap_8 FILLER_73_781 ();
 sg13g2_fill_2 FILLER_73_818 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_fill_1 FILLER_73_858 ();
 sg13g2_fill_2 FILLER_73_864 ();
 sg13g2_fill_1 FILLER_73_892 ();
 sg13g2_decap_8 FILLER_73_900 ();
 sg13g2_fill_1 FILLER_73_907 ();
 sg13g2_fill_1 FILLER_73_934 ();
 sg13g2_fill_1 FILLER_73_961 ();
 sg13g2_fill_1 FILLER_73_991 ();
 sg13g2_fill_2 FILLER_73_1003 ();
 sg13g2_fill_1 FILLER_73_1012 ();
 sg13g2_fill_1 FILLER_73_1054 ();
 sg13g2_fill_1 FILLER_73_1073 ();
 sg13g2_fill_1 FILLER_73_1133 ();
 sg13g2_decap_8 FILLER_73_1144 ();
 sg13g2_decap_4 FILLER_73_1151 ();
 sg13g2_fill_1 FILLER_73_1155 ();
 sg13g2_decap_8 FILLER_73_1229 ();
 sg13g2_decap_8 FILLER_73_1245 ();
 sg13g2_decap_4 FILLER_73_1252 ();
 sg13g2_fill_2 FILLER_73_1336 ();
 sg13g2_fill_1 FILLER_73_1338 ();
 sg13g2_fill_1 FILLER_73_1348 ();
 sg13g2_fill_1 FILLER_73_1364 ();
 sg13g2_fill_2 FILLER_73_1395 ();
 sg13g2_decap_8 FILLER_73_1423 ();
 sg13g2_fill_2 FILLER_73_1430 ();
 sg13g2_decap_4 FILLER_73_1451 ();
 sg13g2_decap_8 FILLER_73_1472 ();
 sg13g2_fill_1 FILLER_73_1511 ();
 sg13g2_decap_4 FILLER_73_1602 ();
 sg13g2_fill_2 FILLER_73_1679 ();
 sg13g2_decap_8 FILLER_73_1765 ();
 sg13g2_decap_4 FILLER_73_1772 ();
 sg13g2_fill_2 FILLER_73_1776 ();
 sg13g2_fill_2 FILLER_73_1790 ();
 sg13g2_fill_1 FILLER_73_1831 ();
 sg13g2_decap_8 FILLER_73_1868 ();
 sg13g2_decap_4 FILLER_73_1875 ();
 sg13g2_fill_1 FILLER_73_1879 ();
 sg13g2_fill_1 FILLER_73_1923 ();
 sg13g2_fill_2 FILLER_73_1929 ();
 sg13g2_fill_2 FILLER_73_1956 ();
 sg13g2_fill_1 FILLER_73_1958 ();
 sg13g2_decap_8 FILLER_73_1963 ();
 sg13g2_decap_8 FILLER_73_1970 ();
 sg13g2_fill_2 FILLER_73_1977 ();
 sg13g2_decap_4 FILLER_73_1996 ();
 sg13g2_fill_2 FILLER_73_2000 ();
 sg13g2_decap_8 FILLER_73_2015 ();
 sg13g2_decap_4 FILLER_73_2022 ();
 sg13g2_fill_2 FILLER_73_2026 ();
 sg13g2_decap_4 FILLER_73_2032 ();
 sg13g2_fill_2 FILLER_73_2107 ();
 sg13g2_fill_1 FILLER_73_2109 ();
 sg13g2_fill_2 FILLER_73_2136 ();
 sg13g2_fill_2 FILLER_73_2142 ();
 sg13g2_fill_2 FILLER_73_2152 ();
 sg13g2_fill_1 FILLER_73_2154 ();
 sg13g2_decap_4 FILLER_73_2165 ();
 sg13g2_fill_2 FILLER_73_2169 ();
 sg13g2_decap_8 FILLER_73_2175 ();
 sg13g2_decap_4 FILLER_73_2182 ();
 sg13g2_fill_2 FILLER_73_2186 ();
 sg13g2_fill_2 FILLER_73_2203 ();
 sg13g2_fill_1 FILLER_73_2222 ();
 sg13g2_fill_2 FILLER_73_2265 ();
 sg13g2_fill_1 FILLER_73_2267 ();
 sg13g2_decap_8 FILLER_73_2273 ();
 sg13g2_decap_4 FILLER_73_2280 ();
 sg13g2_fill_1 FILLER_73_2284 ();
 sg13g2_decap_4 FILLER_73_2296 ();
 sg13g2_fill_2 FILLER_73_2300 ();
 sg13g2_fill_2 FILLER_73_2311 ();
 sg13g2_fill_1 FILLER_73_2313 ();
 sg13g2_decap_4 FILLER_73_2345 ();
 sg13g2_fill_2 FILLER_73_2430 ();
 sg13g2_decap_8 FILLER_73_2436 ();
 sg13g2_decap_8 FILLER_73_2443 ();
 sg13g2_decap_8 FILLER_73_2450 ();
 sg13g2_decap_8 FILLER_73_2457 ();
 sg13g2_decap_8 FILLER_73_2464 ();
 sg13g2_decap_8 FILLER_73_2471 ();
 sg13g2_decap_8 FILLER_73_2478 ();
 sg13g2_decap_8 FILLER_73_2485 ();
 sg13g2_decap_8 FILLER_73_2492 ();
 sg13g2_decap_8 FILLER_73_2499 ();
 sg13g2_decap_8 FILLER_73_2506 ();
 sg13g2_decap_8 FILLER_73_2513 ();
 sg13g2_decap_8 FILLER_73_2520 ();
 sg13g2_decap_8 FILLER_73_2527 ();
 sg13g2_decap_8 FILLER_73_2534 ();
 sg13g2_decap_8 FILLER_73_2541 ();
 sg13g2_decap_8 FILLER_73_2548 ();
 sg13g2_decap_8 FILLER_73_2555 ();
 sg13g2_decap_8 FILLER_73_2562 ();
 sg13g2_decap_8 FILLER_73_2569 ();
 sg13g2_decap_8 FILLER_73_2576 ();
 sg13g2_decap_8 FILLER_73_2583 ();
 sg13g2_decap_8 FILLER_73_2590 ();
 sg13g2_decap_8 FILLER_73_2597 ();
 sg13g2_decap_8 FILLER_73_2604 ();
 sg13g2_decap_8 FILLER_73_2611 ();
 sg13g2_decap_8 FILLER_73_2618 ();
 sg13g2_decap_8 FILLER_73_2625 ();
 sg13g2_decap_8 FILLER_73_2632 ();
 sg13g2_decap_8 FILLER_73_2639 ();
 sg13g2_decap_8 FILLER_73_2646 ();
 sg13g2_decap_8 FILLER_73_2653 ();
 sg13g2_decap_8 FILLER_73_2660 ();
 sg13g2_fill_2 FILLER_73_2667 ();
 sg13g2_fill_1 FILLER_73_2669 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_4 FILLER_74_14 ();
 sg13g2_fill_2 FILLER_74_76 ();
 sg13g2_fill_2 FILLER_74_102 ();
 sg13g2_fill_1 FILLER_74_130 ();
 sg13g2_fill_2 FILLER_74_158 ();
 sg13g2_fill_1 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_decap_8 FILLER_74_183 ();
 sg13g2_decap_4 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_194 ();
 sg13g2_fill_2 FILLER_74_204 ();
 sg13g2_fill_1 FILLER_74_206 ();
 sg13g2_fill_2 FILLER_74_211 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_fill_1 FILLER_74_231 ();
 sg13g2_fill_2 FILLER_74_237 ();
 sg13g2_fill_1 FILLER_74_239 ();
 sg13g2_decap_8 FILLER_74_243 ();
 sg13g2_decap_8 FILLER_74_250 ();
 sg13g2_decap_8 FILLER_74_257 ();
 sg13g2_decap_8 FILLER_74_264 ();
 sg13g2_decap_8 FILLER_74_271 ();
 sg13g2_decap_8 FILLER_74_278 ();
 sg13g2_decap_4 FILLER_74_285 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_fill_2 FILLER_74_301 ();
 sg13g2_fill_1 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_74_335 ();
 sg13g2_decap_8 FILLER_74_342 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_384 ();
 sg13g2_decap_8 FILLER_74_391 ();
 sg13g2_decap_4 FILLER_74_490 ();
 sg13g2_fill_1 FILLER_74_494 ();
 sg13g2_decap_8 FILLER_74_517 ();
 sg13g2_decap_8 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_531 ();
 sg13g2_decap_4 FILLER_74_538 ();
 sg13g2_fill_1 FILLER_74_556 ();
 sg13g2_decap_8 FILLER_74_568 ();
 sg13g2_fill_1 FILLER_74_575 ();
 sg13g2_fill_1 FILLER_74_610 ();
 sg13g2_fill_1 FILLER_74_616 ();
 sg13g2_fill_1 FILLER_74_679 ();
 sg13g2_fill_2 FILLER_74_741 ();
 sg13g2_fill_1 FILLER_74_743 ();
 sg13g2_decap_8 FILLER_74_770 ();
 sg13g2_decap_4 FILLER_74_777 ();
 sg13g2_fill_1 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_787 ();
 sg13g2_decap_4 FILLER_74_794 ();
 sg13g2_fill_1 FILLER_74_798 ();
 sg13g2_decap_4 FILLER_74_803 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_4 FILLER_74_818 ();
 sg13g2_fill_1 FILLER_74_822 ();
 sg13g2_fill_1 FILLER_74_836 ();
 sg13g2_decap_4 FILLER_74_861 ();
 sg13g2_fill_1 FILLER_74_880 ();
 sg13g2_fill_2 FILLER_74_942 ();
 sg13g2_fill_2 FILLER_74_996 ();
 sg13g2_fill_2 FILLER_74_1036 ();
 sg13g2_fill_2 FILLER_74_1101 ();
 sg13g2_decap_4 FILLER_74_1117 ();
 sg13g2_fill_2 FILLER_74_1121 ();
 sg13g2_decap_4 FILLER_74_1128 ();
 sg13g2_fill_1 FILLER_74_1136 ();
 sg13g2_decap_4 FILLER_74_1163 ();
 sg13g2_decap_8 FILLER_74_1171 ();
 sg13g2_decap_4 FILLER_74_1178 ();
 sg13g2_fill_1 FILLER_74_1182 ();
 sg13g2_decap_4 FILLER_74_1192 ();
 sg13g2_fill_2 FILLER_74_1201 ();
 sg13g2_fill_1 FILLER_74_1203 ();
 sg13g2_decap_4 FILLER_74_1209 ();
 sg13g2_fill_1 FILLER_74_1265 ();
 sg13g2_decap_8 FILLER_74_1327 ();
 sg13g2_fill_2 FILLER_74_1334 ();
 sg13g2_decap_4 FILLER_74_1341 ();
 sg13g2_fill_2 FILLER_74_1400 ();
 sg13g2_fill_2 FILLER_74_1432 ();
 sg13g2_fill_1 FILLER_74_1434 ();
 sg13g2_decap_4 FILLER_74_1474 ();
 sg13g2_fill_2 FILLER_74_1478 ();
 sg13g2_fill_1 FILLER_74_1487 ();
 sg13g2_decap_8 FILLER_74_1557 ();
 sg13g2_decap_8 FILLER_74_1564 ();
 sg13g2_decap_8 FILLER_74_1571 ();
 sg13g2_decap_8 FILLER_74_1578 ();
 sg13g2_decap_8 FILLER_74_1590 ();
 sg13g2_decap_8 FILLER_74_1597 ();
 sg13g2_fill_1 FILLER_74_1604 ();
 sg13g2_fill_1 FILLER_74_1651 ();
 sg13g2_decap_4 FILLER_74_1694 ();
 sg13g2_fill_1 FILLER_74_1714 ();
 sg13g2_decap_8 FILLER_74_1766 ();
 sg13g2_decap_8 FILLER_74_1773 ();
 sg13g2_decap_4 FILLER_74_1803 ();
 sg13g2_fill_2 FILLER_74_1812 ();
 sg13g2_fill_2 FILLER_74_1857 ();
 sg13g2_fill_1 FILLER_74_1859 ();
 sg13g2_decap_8 FILLER_74_1876 ();
 sg13g2_fill_1 FILLER_74_1889 ();
 sg13g2_fill_2 FILLER_74_1911 ();
 sg13g2_fill_1 FILLER_74_1913 ();
 sg13g2_fill_2 FILLER_74_1919 ();
 sg13g2_fill_1 FILLER_74_1955 ();
 sg13g2_decap_8 FILLER_74_1991 ();
 sg13g2_decap_8 FILLER_74_1998 ();
 sg13g2_fill_1 FILLER_74_2005 ();
 sg13g2_decap_8 FILLER_74_2036 ();
 sg13g2_decap_4 FILLER_74_2043 ();
 sg13g2_fill_1 FILLER_74_2047 ();
 sg13g2_fill_1 FILLER_74_2053 ();
 sg13g2_fill_1 FILLER_74_2089 ();
 sg13g2_fill_1 FILLER_74_2129 ();
 sg13g2_fill_1 FILLER_74_2153 ();
 sg13g2_decap_8 FILLER_74_2157 ();
 sg13g2_decap_8 FILLER_74_2164 ();
 sg13g2_decap_8 FILLER_74_2171 ();
 sg13g2_decap_4 FILLER_74_2178 ();
 sg13g2_fill_1 FILLER_74_2182 ();
 sg13g2_decap_4 FILLER_74_2261 ();
 sg13g2_fill_1 FILLER_74_2265 ();
 sg13g2_decap_4 FILLER_74_2283 ();
 sg13g2_decap_4 FILLER_74_2296 ();
 sg13g2_fill_2 FILLER_74_2300 ();
 sg13g2_fill_1 FILLER_74_2310 ();
 sg13g2_decap_8 FILLER_74_2315 ();
 sg13g2_decap_8 FILLER_74_2322 ();
 sg13g2_fill_2 FILLER_74_2329 ();
 sg13g2_fill_1 FILLER_74_2337 ();
 sg13g2_decap_4 FILLER_74_2344 ();
 sg13g2_fill_2 FILLER_74_2365 ();
 sg13g2_decap_4 FILLER_74_2380 ();
 sg13g2_fill_2 FILLER_74_2384 ();
 sg13g2_decap_8 FILLER_74_2454 ();
 sg13g2_decap_8 FILLER_74_2461 ();
 sg13g2_decap_8 FILLER_74_2468 ();
 sg13g2_decap_8 FILLER_74_2475 ();
 sg13g2_decap_8 FILLER_74_2482 ();
 sg13g2_decap_8 FILLER_74_2489 ();
 sg13g2_decap_8 FILLER_74_2496 ();
 sg13g2_decap_8 FILLER_74_2503 ();
 sg13g2_decap_8 FILLER_74_2510 ();
 sg13g2_decap_8 FILLER_74_2517 ();
 sg13g2_decap_8 FILLER_74_2524 ();
 sg13g2_decap_8 FILLER_74_2531 ();
 sg13g2_decap_8 FILLER_74_2538 ();
 sg13g2_decap_8 FILLER_74_2545 ();
 sg13g2_decap_8 FILLER_74_2552 ();
 sg13g2_decap_8 FILLER_74_2559 ();
 sg13g2_decap_8 FILLER_74_2566 ();
 sg13g2_decap_8 FILLER_74_2573 ();
 sg13g2_decap_8 FILLER_74_2580 ();
 sg13g2_decap_8 FILLER_74_2587 ();
 sg13g2_decap_8 FILLER_74_2594 ();
 sg13g2_decap_8 FILLER_74_2601 ();
 sg13g2_decap_8 FILLER_74_2608 ();
 sg13g2_decap_8 FILLER_74_2615 ();
 sg13g2_decap_8 FILLER_74_2622 ();
 sg13g2_decap_8 FILLER_74_2629 ();
 sg13g2_decap_8 FILLER_74_2636 ();
 sg13g2_decap_8 FILLER_74_2643 ();
 sg13g2_decap_8 FILLER_74_2650 ();
 sg13g2_decap_8 FILLER_74_2657 ();
 sg13g2_decap_4 FILLER_74_2664 ();
 sg13g2_fill_2 FILLER_74_2668 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_21 ();
 sg13g2_fill_2 FILLER_75_68 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_fill_1 FILLER_75_82 ();
 sg13g2_fill_1 FILLER_75_96 ();
 sg13g2_fill_2 FILLER_75_134 ();
 sg13g2_fill_1 FILLER_75_156 ();
 sg13g2_fill_1 FILLER_75_164 ();
 sg13g2_decap_4 FILLER_75_171 ();
 sg13g2_fill_2 FILLER_75_209 ();
 sg13g2_fill_1 FILLER_75_211 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_fill_2 FILLER_75_224 ();
 sg13g2_fill_1 FILLER_75_226 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_decap_4 FILLER_75_248 ();
 sg13g2_fill_1 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_286 ();
 sg13g2_decap_8 FILLER_75_319 ();
 sg13g2_fill_1 FILLER_75_326 ();
 sg13g2_fill_1 FILLER_75_371 ();
 sg13g2_fill_2 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_389 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_decap_8 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_410 ();
 sg13g2_decap_4 FILLER_75_424 ();
 sg13g2_fill_1 FILLER_75_428 ();
 sg13g2_fill_2 FILLER_75_453 ();
 sg13g2_fill_2 FILLER_75_459 ();
 sg13g2_decap_4 FILLER_75_465 ();
 sg13g2_fill_1 FILLER_75_469 ();
 sg13g2_decap_8 FILLER_75_480 ();
 sg13g2_decap_8 FILLER_75_497 ();
 sg13g2_decap_4 FILLER_75_504 ();
 sg13g2_fill_1 FILLER_75_508 ();
 sg13g2_fill_2 FILLER_75_513 ();
 sg13g2_decap_8 FILLER_75_519 ();
 sg13g2_fill_1 FILLER_75_526 ();
 sg13g2_fill_1 FILLER_75_536 ();
 sg13g2_fill_1 FILLER_75_541 ();
 sg13g2_fill_2 FILLER_75_557 ();
 sg13g2_decap_8 FILLER_75_590 ();
 sg13g2_fill_2 FILLER_75_597 ();
 sg13g2_fill_1 FILLER_75_599 ();
 sg13g2_fill_1 FILLER_75_620 ();
 sg13g2_fill_1 FILLER_75_631 ();
 sg13g2_fill_1 FILLER_75_637 ();
 sg13g2_decap_8 FILLER_75_656 ();
 sg13g2_fill_2 FILLER_75_667 ();
 sg13g2_decap_8 FILLER_75_673 ();
 sg13g2_decap_4 FILLER_75_685 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_731 ();
 sg13g2_decap_8 FILLER_75_738 ();
 sg13g2_decap_4 FILLER_75_745 ();
 sg13g2_fill_2 FILLER_75_749 ();
 sg13g2_fill_1 FILLER_75_755 ();
 sg13g2_fill_2 FILLER_75_760 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_4 FILLER_75_780 ();
 sg13g2_fill_1 FILLER_75_784 ();
 sg13g2_decap_4 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_fill_1 FILLER_75_832 ();
 sg13g2_fill_1 FILLER_75_845 ();
 sg13g2_fill_1 FILLER_75_872 ();
 sg13g2_fill_2 FILLER_75_909 ();
 sg13g2_decap_8 FILLER_75_915 ();
 sg13g2_fill_2 FILLER_75_922 ();
 sg13g2_fill_1 FILLER_75_924 ();
 sg13g2_fill_1 FILLER_75_940 ();
 sg13g2_fill_1 FILLER_75_999 ();
 sg13g2_fill_2 FILLER_75_1059 ();
 sg13g2_fill_2 FILLER_75_1121 ();
 sg13g2_fill_2 FILLER_75_1162 ();
 sg13g2_decap_8 FILLER_75_1174 ();
 sg13g2_fill_1 FILLER_75_1181 ();
 sg13g2_decap_4 FILLER_75_1208 ();
 sg13g2_fill_1 FILLER_75_1212 ();
 sg13g2_fill_2 FILLER_75_1239 ();
 sg13g2_fill_2 FILLER_75_1245 ();
 sg13g2_decap_8 FILLER_75_1255 ();
 sg13g2_decap_8 FILLER_75_1262 ();
 sg13g2_decap_8 FILLER_75_1269 ();
 sg13g2_decap_8 FILLER_75_1276 ();
 sg13g2_decap_8 FILLER_75_1283 ();
 sg13g2_decap_8 FILLER_75_1290 ();
 sg13g2_fill_2 FILLER_75_1297 ();
 sg13g2_fill_1 FILLER_75_1299 ();
 sg13g2_decap_8 FILLER_75_1330 ();
 sg13g2_decap_8 FILLER_75_1337 ();
 sg13g2_decap_8 FILLER_75_1344 ();
 sg13g2_decap_4 FILLER_75_1351 ();
 sg13g2_fill_2 FILLER_75_1355 ();
 sg13g2_decap_4 FILLER_75_1360 ();
 sg13g2_decap_4 FILLER_75_1394 ();
 sg13g2_decap_8 FILLER_75_1402 ();
 sg13g2_fill_2 FILLER_75_1409 ();
 sg13g2_fill_1 FILLER_75_1411 ();
 sg13g2_fill_1 FILLER_75_1452 ();
 sg13g2_decap_8 FILLER_75_1457 ();
 sg13g2_decap_8 FILLER_75_1464 ();
 sg13g2_fill_2 FILLER_75_1471 ();
 sg13g2_fill_1 FILLER_75_1473 ();
 sg13g2_fill_1 FILLER_75_1513 ();
 sg13g2_decap_8 FILLER_75_1561 ();
 sg13g2_decap_8 FILLER_75_1573 ();
 sg13g2_decap_8 FILLER_75_1580 ();
 sg13g2_decap_4 FILLER_75_1587 ();
 sg13g2_decap_8 FILLER_75_1595 ();
 sg13g2_decap_8 FILLER_75_1602 ();
 sg13g2_fill_2 FILLER_75_1609 ();
 sg13g2_fill_1 FILLER_75_1611 ();
 sg13g2_decap_8 FILLER_75_1638 ();
 sg13g2_decap_8 FILLER_75_1645 ();
 sg13g2_fill_2 FILLER_75_1652 ();
 sg13g2_decap_8 FILLER_75_1676 ();
 sg13g2_decap_8 FILLER_75_1683 ();
 sg13g2_decap_4 FILLER_75_1690 ();
 sg13g2_fill_1 FILLER_75_1694 ();
 sg13g2_decap_4 FILLER_75_1702 ();
 sg13g2_fill_1 FILLER_75_1706 ();
 sg13g2_decap_8 FILLER_75_1711 ();
 sg13g2_decap_8 FILLER_75_1718 ();
 sg13g2_decap_4 FILLER_75_1725 ();
 sg13g2_fill_1 FILLER_75_1729 ();
 sg13g2_fill_2 FILLER_75_1739 ();
 sg13g2_fill_1 FILLER_75_1741 ();
 sg13g2_fill_2 FILLER_75_1751 ();
 sg13g2_fill_1 FILLER_75_1756 ();
 sg13g2_decap_4 FILLER_75_1783 ();
 sg13g2_fill_2 FILLER_75_1787 ();
 sg13g2_fill_1 FILLER_75_1845 ();
 sg13g2_decap_8 FILLER_75_1872 ();
 sg13g2_decap_8 FILLER_75_1879 ();
 sg13g2_decap_8 FILLER_75_1886 ();
 sg13g2_decap_8 FILLER_75_1893 ();
 sg13g2_decap_8 FILLER_75_1900 ();
 sg13g2_decap_4 FILLER_75_1907 ();
 sg13g2_fill_2 FILLER_75_1911 ();
 sg13g2_decap_8 FILLER_75_1943 ();
 sg13g2_fill_2 FILLER_75_1950 ();
 sg13g2_decap_8 FILLER_75_1957 ();
 sg13g2_fill_2 FILLER_75_1964 ();
 sg13g2_fill_2 FILLER_75_1975 ();
 sg13g2_decap_8 FILLER_75_2016 ();
 sg13g2_decap_8 FILLER_75_2023 ();
 sg13g2_decap_8 FILLER_75_2030 ();
 sg13g2_decap_8 FILLER_75_2037 ();
 sg13g2_decap_8 FILLER_75_2044 ();
 sg13g2_decap_8 FILLER_75_2051 ();
 sg13g2_fill_2 FILLER_75_2071 ();
 sg13g2_fill_2 FILLER_75_2125 ();
 sg13g2_fill_1 FILLER_75_2135 ();
 sg13g2_fill_2 FILLER_75_2152 ();
 sg13g2_decap_8 FILLER_75_2167 ();
 sg13g2_decap_4 FILLER_75_2174 ();
 sg13g2_fill_2 FILLER_75_2178 ();
 sg13g2_decap_8 FILLER_75_2186 ();
 sg13g2_fill_2 FILLER_75_2193 ();
 sg13g2_fill_1 FILLER_75_2225 ();
 sg13g2_decap_8 FILLER_75_2231 ();
 sg13g2_decap_8 FILLER_75_2238 ();
 sg13g2_fill_2 FILLER_75_2245 ();
 sg13g2_decap_8 FILLER_75_2260 ();
 sg13g2_fill_1 FILLER_75_2267 ();
 sg13g2_decap_8 FILLER_75_2293 ();
 sg13g2_decap_4 FILLER_75_2300 ();
 sg13g2_fill_2 FILLER_75_2308 ();
 sg13g2_fill_2 FILLER_75_2314 ();
 sg13g2_fill_1 FILLER_75_2316 ();
 sg13g2_decap_4 FILLER_75_2335 ();
 sg13g2_fill_1 FILLER_75_2339 ();
 sg13g2_decap_8 FILLER_75_2344 ();
 sg13g2_decap_8 FILLER_75_2351 ();
 sg13g2_decap_8 FILLER_75_2358 ();
 sg13g2_decap_8 FILLER_75_2365 ();
 sg13g2_decap_8 FILLER_75_2377 ();
 sg13g2_decap_8 FILLER_75_2384 ();
 sg13g2_fill_1 FILLER_75_2391 ();
 sg13g2_decap_8 FILLER_75_2404 ();
 sg13g2_decap_8 FILLER_75_2411 ();
 sg13g2_decap_8 FILLER_75_2418 ();
 sg13g2_fill_2 FILLER_75_2425 ();
 sg13g2_fill_1 FILLER_75_2427 ();
 sg13g2_decap_8 FILLER_75_2454 ();
 sg13g2_decap_8 FILLER_75_2461 ();
 sg13g2_decap_8 FILLER_75_2468 ();
 sg13g2_decap_8 FILLER_75_2475 ();
 sg13g2_decap_8 FILLER_75_2482 ();
 sg13g2_decap_8 FILLER_75_2489 ();
 sg13g2_decap_8 FILLER_75_2496 ();
 sg13g2_decap_8 FILLER_75_2503 ();
 sg13g2_decap_8 FILLER_75_2510 ();
 sg13g2_decap_8 FILLER_75_2517 ();
 sg13g2_decap_8 FILLER_75_2524 ();
 sg13g2_decap_8 FILLER_75_2531 ();
 sg13g2_decap_8 FILLER_75_2538 ();
 sg13g2_decap_8 FILLER_75_2545 ();
 sg13g2_decap_8 FILLER_75_2552 ();
 sg13g2_decap_8 FILLER_75_2559 ();
 sg13g2_decap_8 FILLER_75_2566 ();
 sg13g2_decap_8 FILLER_75_2573 ();
 sg13g2_decap_8 FILLER_75_2580 ();
 sg13g2_decap_8 FILLER_75_2587 ();
 sg13g2_decap_8 FILLER_75_2594 ();
 sg13g2_decap_8 FILLER_75_2601 ();
 sg13g2_decap_8 FILLER_75_2608 ();
 sg13g2_decap_8 FILLER_75_2615 ();
 sg13g2_decap_8 FILLER_75_2622 ();
 sg13g2_decap_8 FILLER_75_2629 ();
 sg13g2_decap_8 FILLER_75_2636 ();
 sg13g2_decap_8 FILLER_75_2643 ();
 sg13g2_decap_8 FILLER_75_2650 ();
 sg13g2_decap_8 FILLER_75_2657 ();
 sg13g2_decap_4 FILLER_75_2664 ();
 sg13g2_fill_2 FILLER_75_2668 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_47 ();
 sg13g2_fill_2 FILLER_76_51 ();
 sg13g2_decap_4 FILLER_76_90 ();
 sg13g2_fill_2 FILLER_76_103 ();
 sg13g2_fill_1 FILLER_76_119 ();
 sg13g2_fill_1 FILLER_76_125 ();
 sg13g2_fill_1 FILLER_76_132 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_160 ();
 sg13g2_fill_2 FILLER_76_179 ();
 sg13g2_fill_1 FILLER_76_181 ();
 sg13g2_fill_1 FILLER_76_187 ();
 sg13g2_fill_2 FILLER_76_193 ();
 sg13g2_fill_2 FILLER_76_220 ();
 sg13g2_fill_2 FILLER_76_268 ();
 sg13g2_fill_1 FILLER_76_270 ();
 sg13g2_decap_4 FILLER_76_288 ();
 sg13g2_fill_2 FILLER_76_292 ();
 sg13g2_fill_2 FILLER_76_299 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_328 ();
 sg13g2_decap_8 FILLER_76_335 ();
 sg13g2_decap_8 FILLER_76_342 ();
 sg13g2_decap_8 FILLER_76_349 ();
 sg13g2_decap_8 FILLER_76_356 ();
 sg13g2_decap_8 FILLER_76_363 ();
 sg13g2_decap_8 FILLER_76_370 ();
 sg13g2_fill_2 FILLER_76_377 ();
 sg13g2_fill_1 FILLER_76_379 ();
 sg13g2_fill_2 FILLER_76_393 ();
 sg13g2_fill_1 FILLER_76_395 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_fill_2 FILLER_76_413 ();
 sg13g2_fill_1 FILLER_76_415 ();
 sg13g2_fill_2 FILLER_76_429 ();
 sg13g2_fill_2 FILLER_76_465 ();
 sg13g2_fill_1 FILLER_76_467 ();
 sg13g2_fill_2 FILLER_76_477 ();
 sg13g2_decap_4 FILLER_76_522 ();
 sg13g2_decap_8 FILLER_76_531 ();
 sg13g2_fill_2 FILLER_76_538 ();
 sg13g2_decap_4 FILLER_76_560 ();
 sg13g2_decap_4 FILLER_76_567 ();
 sg13g2_fill_2 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_fill_1 FILLER_76_585 ();
 sg13g2_decap_4 FILLER_76_590 ();
 sg13g2_fill_1 FILLER_76_594 ();
 sg13g2_decap_8 FILLER_76_600 ();
 sg13g2_decap_4 FILLER_76_607 ();
 sg13g2_decap_4 FILLER_76_618 ();
 sg13g2_fill_1 FILLER_76_622 ();
 sg13g2_fill_2 FILLER_76_629 ();
 sg13g2_decap_4 FILLER_76_641 ();
 sg13g2_fill_2 FILLER_76_652 ();
 sg13g2_fill_1 FILLER_76_654 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_decap_8 FILLER_76_665 ();
 sg13g2_decap_8 FILLER_76_672 ();
 sg13g2_decap_8 FILLER_76_679 ();
 sg13g2_decap_8 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_693 ();
 sg13g2_decap_8 FILLER_76_700 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_714 ();
 sg13g2_fill_1 FILLER_76_721 ();
 sg13g2_fill_2 FILLER_76_752 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_fill_1 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_fill_2 FILLER_76_844 ();
 sg13g2_fill_2 FILLER_76_853 ();
 sg13g2_decap_8 FILLER_76_917 ();
 sg13g2_decap_4 FILLER_76_928 ();
 sg13g2_fill_1 FILLER_76_938 ();
 sg13g2_decap_8 FILLER_76_946 ();
 sg13g2_decap_8 FILLER_76_953 ();
 sg13g2_decap_8 FILLER_76_960 ();
 sg13g2_decap_8 FILLER_76_967 ();
 sg13g2_decap_4 FILLER_76_974 ();
 sg13g2_fill_1 FILLER_76_978 ();
 sg13g2_decap_8 FILLER_76_983 ();
 sg13g2_fill_1 FILLER_76_1044 ();
 sg13g2_fill_2 FILLER_76_1054 ();
 sg13g2_fill_1 FILLER_76_1063 ();
 sg13g2_fill_1 FILLER_76_1098 ();
 sg13g2_decap_8 FILLER_76_1121 ();
 sg13g2_decap_8 FILLER_76_1128 ();
 sg13g2_decap_8 FILLER_76_1135 ();
 sg13g2_decap_8 FILLER_76_1142 ();
 sg13g2_decap_8 FILLER_76_1149 ();
 sg13g2_decap_8 FILLER_76_1156 ();
 sg13g2_decap_8 FILLER_76_1163 ();
 sg13g2_decap_8 FILLER_76_1170 ();
 sg13g2_fill_1 FILLER_76_1177 ();
 sg13g2_decap_8 FILLER_76_1182 ();
 sg13g2_decap_4 FILLER_76_1189 ();
 sg13g2_decap_4 FILLER_76_1208 ();
 sg13g2_decap_8 FILLER_76_1229 ();
 sg13g2_decap_8 FILLER_76_1236 ();
 sg13g2_fill_2 FILLER_76_1283 ();
 sg13g2_fill_1 FILLER_76_1285 ();
 sg13g2_decap_8 FILLER_76_1290 ();
 sg13g2_decap_8 FILLER_76_1297 ();
 sg13g2_decap_8 FILLER_76_1304 ();
 sg13g2_decap_8 FILLER_76_1311 ();
 sg13g2_decap_8 FILLER_76_1322 ();
 sg13g2_decap_4 FILLER_76_1329 ();
 sg13g2_fill_1 FILLER_76_1333 ();
 sg13g2_fill_2 FILLER_76_1364 ();
 sg13g2_decap_8 FILLER_76_1379 ();
 sg13g2_fill_1 FILLER_76_1386 ();
 sg13g2_decap_8 FILLER_76_1392 ();
 sg13g2_fill_1 FILLER_76_1399 ();
 sg13g2_decap_4 FILLER_76_1404 ();
 sg13g2_decap_4 FILLER_76_1412 ();
 sg13g2_decap_8 FILLER_76_1420 ();
 sg13g2_decap_8 FILLER_76_1427 ();
 sg13g2_fill_2 FILLER_76_1443 ();
 sg13g2_decap_4 FILLER_76_1478 ();
 sg13g2_decap_8 FILLER_76_1486 ();
 sg13g2_fill_2 FILLER_76_1493 ();
 sg13g2_decap_8 FILLER_76_1521 ();
 sg13g2_fill_2 FILLER_76_1528 ();
 sg13g2_fill_1 FILLER_76_1530 ();
 sg13g2_decap_8 FILLER_76_1544 ();
 sg13g2_decap_4 FILLER_76_1551 ();
 sg13g2_fill_1 FILLER_76_1555 ();
 sg13g2_fill_2 FILLER_76_1595 ();
 sg13g2_fill_1 FILLER_76_1597 ();
 sg13g2_decap_8 FILLER_76_1625 ();
 sg13g2_decap_8 FILLER_76_1632 ();
 sg13g2_decap_4 FILLER_76_1639 ();
 sg13g2_decap_4 FILLER_76_1679 ();
 sg13g2_fill_2 FILLER_76_1687 ();
 sg13g2_fill_1 FILLER_76_1689 ();
 sg13g2_decap_4 FILLER_76_1695 ();
 sg13g2_decap_4 FILLER_76_1707 ();
 sg13g2_decap_4 FILLER_76_1715 ();
 sg13g2_fill_1 FILLER_76_1719 ();
 sg13g2_fill_1 FILLER_76_1725 ();
 sg13g2_fill_1 FILLER_76_1730 ();
 sg13g2_decap_8 FILLER_76_1766 ();
 sg13g2_decap_8 FILLER_76_1773 ();
 sg13g2_decap_8 FILLER_76_1780 ();
 sg13g2_fill_1 FILLER_76_1813 ();
 sg13g2_fill_1 FILLER_76_1817 ();
 sg13g2_decap_8 FILLER_76_1893 ();
 sg13g2_decap_4 FILLER_76_1900 ();
 sg13g2_fill_2 FILLER_76_1904 ();
 sg13g2_fill_2 FILLER_76_1935 ();
 sg13g2_fill_1 FILLER_76_1946 ();
 sg13g2_decap_8 FILLER_76_1951 ();
 sg13g2_decap_4 FILLER_76_1958 ();
 sg13g2_decap_8 FILLER_76_1996 ();
 sg13g2_decap_8 FILLER_76_2003 ();
 sg13g2_fill_2 FILLER_76_2010 ();
 sg13g2_fill_1 FILLER_76_2012 ();
 sg13g2_fill_1 FILLER_76_2044 ();
 sg13g2_fill_1 FILLER_76_2049 ();
 sg13g2_fill_1 FILLER_76_2055 ();
 sg13g2_fill_1 FILLER_76_2060 ();
 sg13g2_decap_8 FILLER_76_2091 ();
 sg13g2_decap_8 FILLER_76_2098 ();
 sg13g2_fill_2 FILLER_76_2105 ();
 sg13g2_fill_2 FILLER_76_2127 ();
 sg13g2_decap_8 FILLER_76_2185 ();
 sg13g2_fill_1 FILLER_76_2192 ();
 sg13g2_fill_2 FILLER_76_2206 ();
 sg13g2_fill_1 FILLER_76_2208 ();
 sg13g2_decap_8 FILLER_76_2234 ();
 sg13g2_decap_4 FILLER_76_2241 ();
 sg13g2_fill_2 FILLER_76_2245 ();
 sg13g2_decap_8 FILLER_76_2256 ();
 sg13g2_decap_8 FILLER_76_2263 ();
 sg13g2_decap_8 FILLER_76_2270 ();
 sg13g2_decap_8 FILLER_76_2277 ();
 sg13g2_decap_8 FILLER_76_2284 ();
 sg13g2_decap_8 FILLER_76_2291 ();
 sg13g2_fill_1 FILLER_76_2298 ();
 sg13g2_fill_1 FILLER_76_2302 ();
 sg13g2_decap_8 FILLER_76_2313 ();
 sg13g2_decap_8 FILLER_76_2320 ();
 sg13g2_decap_8 FILLER_76_2327 ();
 sg13g2_decap_4 FILLER_76_2360 ();
 sg13g2_fill_1 FILLER_76_2364 ();
 sg13g2_decap_8 FILLER_76_2375 ();
 sg13g2_decap_8 FILLER_76_2382 ();
 sg13g2_decap_8 FILLER_76_2389 ();
 sg13g2_decap_8 FILLER_76_2396 ();
 sg13g2_decap_4 FILLER_76_2403 ();
 sg13g2_fill_1 FILLER_76_2407 ();
 sg13g2_decap_4 FILLER_76_2428 ();
 sg13g2_fill_2 FILLER_76_2436 ();
 sg13g2_decap_8 FILLER_76_2442 ();
 sg13g2_decap_8 FILLER_76_2449 ();
 sg13g2_decap_8 FILLER_76_2456 ();
 sg13g2_decap_8 FILLER_76_2463 ();
 sg13g2_decap_8 FILLER_76_2470 ();
 sg13g2_decap_8 FILLER_76_2477 ();
 sg13g2_decap_8 FILLER_76_2484 ();
 sg13g2_decap_8 FILLER_76_2491 ();
 sg13g2_decap_8 FILLER_76_2498 ();
 sg13g2_decap_8 FILLER_76_2505 ();
 sg13g2_decap_8 FILLER_76_2512 ();
 sg13g2_decap_8 FILLER_76_2519 ();
 sg13g2_decap_8 FILLER_76_2526 ();
 sg13g2_decap_8 FILLER_76_2533 ();
 sg13g2_decap_8 FILLER_76_2540 ();
 sg13g2_decap_8 FILLER_76_2547 ();
 sg13g2_decap_8 FILLER_76_2554 ();
 sg13g2_decap_8 FILLER_76_2561 ();
 sg13g2_decap_8 FILLER_76_2568 ();
 sg13g2_decap_8 FILLER_76_2575 ();
 sg13g2_decap_8 FILLER_76_2582 ();
 sg13g2_decap_8 FILLER_76_2589 ();
 sg13g2_decap_8 FILLER_76_2596 ();
 sg13g2_decap_8 FILLER_76_2603 ();
 sg13g2_decap_8 FILLER_76_2610 ();
 sg13g2_decap_8 FILLER_76_2617 ();
 sg13g2_decap_8 FILLER_76_2624 ();
 sg13g2_decap_8 FILLER_76_2631 ();
 sg13g2_decap_8 FILLER_76_2638 ();
 sg13g2_decap_8 FILLER_76_2645 ();
 sg13g2_decap_8 FILLER_76_2652 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_4 FILLER_76_2666 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_59 ();
 sg13g2_fill_1 FILLER_77_99 ();
 sg13g2_fill_1 FILLER_77_171 ();
 sg13g2_decap_4 FILLER_77_176 ();
 sg13g2_fill_2 FILLER_77_215 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_2 FILLER_77_246 ();
 sg13g2_decap_8 FILLER_77_256 ();
 sg13g2_fill_2 FILLER_77_263 ();
 sg13g2_fill_1 FILLER_77_265 ();
 sg13g2_decap_4 FILLER_77_297 ();
 sg13g2_fill_1 FILLER_77_306 ();
 sg13g2_fill_1 FILLER_77_367 ();
 sg13g2_fill_2 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_424 ();
 sg13g2_decap_8 FILLER_77_431 ();
 sg13g2_fill_1 FILLER_77_438 ();
 sg13g2_fill_2 FILLER_77_470 ();
 sg13g2_fill_2 FILLER_77_476 ();
 sg13g2_fill_1 FILLER_77_478 ();
 sg13g2_decap_4 FILLER_77_489 ();
 sg13g2_fill_2 FILLER_77_493 ();
 sg13g2_fill_2 FILLER_77_505 ();
 sg13g2_fill_1 FILLER_77_507 ();
 sg13g2_decap_8 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_519 ();
 sg13g2_fill_1 FILLER_77_560 ();
 sg13g2_fill_1 FILLER_77_570 ();
 sg13g2_decap_8 FILLER_77_610 ();
 sg13g2_decap_8 FILLER_77_617 ();
 sg13g2_decap_8 FILLER_77_624 ();
 sg13g2_fill_1 FILLER_77_631 ();
 sg13g2_fill_2 FILLER_77_636 ();
 sg13g2_fill_1 FILLER_77_638 ();
 sg13g2_decap_4 FILLER_77_699 ();
 sg13g2_fill_2 FILLER_77_703 ();
 sg13g2_decap_4 FILLER_77_713 ();
 sg13g2_fill_2 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_753 ();
 sg13g2_fill_1 FILLER_77_786 ();
 sg13g2_fill_2 FILLER_77_791 ();
 sg13g2_decap_4 FILLER_77_801 ();
 sg13g2_fill_1 FILLER_77_805 ();
 sg13g2_fill_1 FILLER_77_814 ();
 sg13g2_fill_1 FILLER_77_841 ();
 sg13g2_fill_1 FILLER_77_868 ();
 sg13g2_fill_2 FILLER_77_873 ();
 sg13g2_fill_1 FILLER_77_875 ();
 sg13g2_fill_2 FILLER_77_879 ();
 sg13g2_fill_1 FILLER_77_881 ();
 sg13g2_decap_8 FILLER_77_893 ();
 sg13g2_fill_1 FILLER_77_900 ();
 sg13g2_decap_4 FILLER_77_965 ();
 sg13g2_decap_4 FILLER_77_973 ();
 sg13g2_fill_2 FILLER_77_977 ();
 sg13g2_decap_4 FILLER_77_1009 ();
 sg13g2_decap_8 FILLER_77_1031 ();
 sg13g2_decap_8 FILLER_77_1038 ();
 sg13g2_fill_1 FILLER_77_1097 ();
 sg13g2_decap_8 FILLER_77_1135 ();
 sg13g2_fill_2 FILLER_77_1142 ();
 sg13g2_fill_1 FILLER_77_1144 ();
 sg13g2_decap_8 FILLER_77_1171 ();
 sg13g2_decap_4 FILLER_77_1178 ();
 sg13g2_fill_1 FILLER_77_1182 ();
 sg13g2_fill_2 FILLER_77_1191 ();
 sg13g2_decap_8 FILLER_77_1200 ();
 sg13g2_fill_2 FILLER_77_1207 ();
 sg13g2_fill_1 FILLER_77_1209 ();
 sg13g2_decap_8 FILLER_77_1244 ();
 sg13g2_decap_4 FILLER_77_1251 ();
 sg13g2_fill_2 FILLER_77_1255 ();
 sg13g2_decap_8 FILLER_77_1261 ();
 sg13g2_decap_4 FILLER_77_1268 ();
 sg13g2_fill_1 FILLER_77_1280 ();
 sg13g2_fill_1 FILLER_77_1311 ();
 sg13g2_decap_8 FILLER_77_1338 ();
 sg13g2_decap_8 FILLER_77_1345 ();
 sg13g2_fill_1 FILLER_77_1352 ();
 sg13g2_fill_2 FILLER_77_1361 ();
 sg13g2_fill_1 FILLER_77_1363 ();
 sg13g2_decap_8 FILLER_77_1368 ();
 sg13g2_decap_8 FILLER_77_1375 ();
 sg13g2_fill_2 FILLER_77_1382 ();
 sg13g2_decap_4 FILLER_77_1415 ();
 sg13g2_fill_2 FILLER_77_1419 ();
 sg13g2_fill_1 FILLER_77_1460 ();
 sg13g2_decap_8 FILLER_77_1487 ();
 sg13g2_fill_1 FILLER_77_1494 ();
 sg13g2_decap_4 FILLER_77_1530 ();
 sg13g2_fill_1 FILLER_77_1534 ();
 sg13g2_fill_2 FILLER_77_1584 ();
 sg13g2_fill_1 FILLER_77_1586 ();
 sg13g2_fill_2 FILLER_77_1613 ();
 sg13g2_fill_1 FILLER_77_1615 ();
 sg13g2_decap_4 FILLER_77_1621 ();
 sg13g2_fill_1 FILLER_77_1629 ();
 sg13g2_fill_1 FILLER_77_1635 ();
 sg13g2_fill_2 FILLER_77_1640 ();
 sg13g2_decap_4 FILLER_77_1672 ();
 sg13g2_fill_2 FILLER_77_1676 ();
 sg13g2_fill_2 FILLER_77_1709 ();
 sg13g2_fill_1 FILLER_77_1716 ();
 sg13g2_fill_1 FILLER_77_1743 ();
 sg13g2_fill_1 FILLER_77_1749 ();
 sg13g2_decap_8 FILLER_77_1776 ();
 sg13g2_fill_2 FILLER_77_1783 ();
 sg13g2_decap_8 FILLER_77_1789 ();
 sg13g2_fill_2 FILLER_77_1800 ();
 sg13g2_fill_1 FILLER_77_1802 ();
 sg13g2_fill_2 FILLER_77_1808 ();
 sg13g2_fill_1 FILLER_77_1810 ();
 sg13g2_fill_2 FILLER_77_1824 ();
 sg13g2_decap_4 FILLER_77_1856 ();
 sg13g2_fill_1 FILLER_77_1860 ();
 sg13g2_decap_4 FILLER_77_1887 ();
 sg13g2_fill_2 FILLER_77_1891 ();
 sg13g2_decap_4 FILLER_77_1898 ();
 sg13g2_fill_2 FILLER_77_1902 ();
 sg13g2_fill_2 FILLER_77_1908 ();
 sg13g2_decap_4 FILLER_77_1967 ();
 sg13g2_fill_1 FILLER_77_1971 ();
 sg13g2_decap_8 FILLER_77_1977 ();
 sg13g2_decap_4 FILLER_77_1984 ();
 sg13g2_fill_2 FILLER_77_1988 ();
 sg13g2_fill_2 FILLER_77_1995 ();
 sg13g2_fill_1 FILLER_77_1997 ();
 sg13g2_fill_1 FILLER_77_2003 ();
 sg13g2_decap_8 FILLER_77_2008 ();
 sg13g2_decap_8 FILLER_77_2015 ();
 sg13g2_fill_2 FILLER_77_2022 ();
 sg13g2_fill_1 FILLER_77_2024 ();
 sg13g2_fill_1 FILLER_77_2060 ();
 sg13g2_fill_2 FILLER_77_2090 ();
 sg13g2_fill_1 FILLER_77_2092 ();
 sg13g2_fill_2 FILLER_77_2097 ();
 sg13g2_decap_4 FILLER_77_2103 ();
 sg13g2_fill_2 FILLER_77_2112 ();
 sg13g2_fill_2 FILLER_77_2149 ();
 sg13g2_fill_1 FILLER_77_2177 ();
 sg13g2_fill_2 FILLER_77_2181 ();
 sg13g2_fill_2 FILLER_77_2209 ();
 sg13g2_fill_1 FILLER_77_2211 ();
 sg13g2_decap_4 FILLER_77_2220 ();
 sg13g2_fill_1 FILLER_77_2224 ();
 sg13g2_decap_8 FILLER_77_2251 ();
 sg13g2_fill_1 FILLER_77_2258 ();
 sg13g2_decap_8 FILLER_77_2285 ();
 sg13g2_decap_8 FILLER_77_2292 ();
 sg13g2_fill_2 FILLER_77_2304 ();
 sg13g2_decap_8 FILLER_77_2345 ();
 sg13g2_decap_8 FILLER_77_2352 ();
 sg13g2_decap_8 FILLER_77_2359 ();
 sg13g2_fill_1 FILLER_77_2366 ();
 sg13g2_decap_8 FILLER_77_2397 ();
 sg13g2_decap_8 FILLER_77_2408 ();
 sg13g2_decap_8 FILLER_77_2436 ();
 sg13g2_decap_8 FILLER_77_2443 ();
 sg13g2_decap_8 FILLER_77_2450 ();
 sg13g2_decap_8 FILLER_77_2457 ();
 sg13g2_decap_8 FILLER_77_2464 ();
 sg13g2_decap_8 FILLER_77_2471 ();
 sg13g2_decap_8 FILLER_77_2478 ();
 sg13g2_decap_8 FILLER_77_2485 ();
 sg13g2_decap_8 FILLER_77_2492 ();
 sg13g2_decap_8 FILLER_77_2499 ();
 sg13g2_decap_8 FILLER_77_2506 ();
 sg13g2_decap_8 FILLER_77_2513 ();
 sg13g2_decap_8 FILLER_77_2520 ();
 sg13g2_decap_8 FILLER_77_2527 ();
 sg13g2_decap_8 FILLER_77_2534 ();
 sg13g2_decap_8 FILLER_77_2541 ();
 sg13g2_decap_8 FILLER_77_2548 ();
 sg13g2_decap_8 FILLER_77_2555 ();
 sg13g2_decap_8 FILLER_77_2562 ();
 sg13g2_decap_8 FILLER_77_2569 ();
 sg13g2_decap_8 FILLER_77_2576 ();
 sg13g2_decap_8 FILLER_77_2583 ();
 sg13g2_decap_8 FILLER_77_2590 ();
 sg13g2_decap_8 FILLER_77_2597 ();
 sg13g2_decap_8 FILLER_77_2604 ();
 sg13g2_decap_8 FILLER_77_2611 ();
 sg13g2_decap_8 FILLER_77_2618 ();
 sg13g2_decap_8 FILLER_77_2625 ();
 sg13g2_decap_8 FILLER_77_2632 ();
 sg13g2_decap_8 FILLER_77_2639 ();
 sg13g2_decap_8 FILLER_77_2646 ();
 sg13g2_decap_8 FILLER_77_2653 ();
 sg13g2_decap_8 FILLER_77_2660 ();
 sg13g2_fill_2 FILLER_77_2667 ();
 sg13g2_fill_1 FILLER_77_2669 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_68 ();
 sg13g2_decap_8 FILLER_78_75 ();
 sg13g2_decap_8 FILLER_78_82 ();
 sg13g2_decap_8 FILLER_78_89 ();
 sg13g2_decap_8 FILLER_78_96 ();
 sg13g2_decap_8 FILLER_78_103 ();
 sg13g2_decap_8 FILLER_78_110 ();
 sg13g2_decap_4 FILLER_78_117 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_4 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_156 ();
 sg13g2_fill_2 FILLER_78_167 ();
 sg13g2_fill_1 FILLER_78_169 ();
 sg13g2_decap_4 FILLER_78_179 ();
 sg13g2_fill_2 FILLER_78_183 ();
 sg13g2_fill_1 FILLER_78_207 ();
 sg13g2_decap_4 FILLER_78_228 ();
 sg13g2_fill_2 FILLER_78_232 ();
 sg13g2_fill_1 FILLER_78_276 ();
 sg13g2_decap_4 FILLER_78_320 ();
 sg13g2_decap_8 FILLER_78_328 ();
 sg13g2_fill_2 FILLER_78_335 ();
 sg13g2_fill_2 FILLER_78_363 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_4 FILLER_78_441 ();
 sg13g2_fill_1 FILLER_78_445 ();
 sg13g2_decap_4 FILLER_78_452 ();
 sg13g2_fill_2 FILLER_78_456 ();
 sg13g2_fill_2 FILLER_78_475 ();
 sg13g2_decap_8 FILLER_78_516 ();
 sg13g2_fill_2 FILLER_78_523 ();
 sg13g2_fill_1 FILLER_78_525 ();
 sg13g2_fill_1 FILLER_78_530 ();
 sg13g2_decap_8 FILLER_78_578 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_fill_2 FILLER_78_623 ();
 sg13g2_fill_1 FILLER_78_625 ();
 sg13g2_fill_1 FILLER_78_652 ();
 sg13g2_fill_1 FILLER_78_670 ();
 sg13g2_fill_2 FILLER_78_710 ();
 sg13g2_fill_1 FILLER_78_712 ();
 sg13g2_fill_2 FILLER_78_743 ();
 sg13g2_fill_1 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_883 ();
 sg13g2_decap_8 FILLER_78_890 ();
 sg13g2_decap_8 FILLER_78_897 ();
 sg13g2_fill_2 FILLER_78_934 ();
 sg13g2_fill_1 FILLER_78_936 ();
 sg13g2_fill_1 FILLER_78_1090 ();
 sg13g2_fill_1 FILLER_78_1100 ();
 sg13g2_decap_4 FILLER_78_1132 ();
 sg13g2_fill_1 FILLER_78_1170 ();
 sg13g2_decap_4 FILLER_78_1201 ();
 sg13g2_fill_2 FILLER_78_1209 ();
 sg13g2_decap_8 FILLER_78_1245 ();
 sg13g2_decap_4 FILLER_78_1252 ();
 sg13g2_fill_2 FILLER_78_1256 ();
 sg13g2_fill_2 FILLER_78_1288 ();
 sg13g2_fill_2 FILLER_78_1324 ();
 sg13g2_fill_1 FILLER_78_1326 ();
 sg13g2_fill_1 FILLER_78_1440 ();
 sg13g2_decap_8 FILLER_78_1468 ();
 sg13g2_decap_8 FILLER_78_1475 ();
 sg13g2_decap_8 FILLER_78_1482 ();
 sg13g2_decap_8 FILLER_78_1489 ();
 sg13g2_decap_8 FILLER_78_1496 ();
 sg13g2_decap_4 FILLER_78_1503 ();
 sg13g2_fill_1 FILLER_78_1507 ();
 sg13g2_decap_8 FILLER_78_1518 ();
 sg13g2_fill_2 FILLER_78_1525 ();
 sg13g2_fill_1 FILLER_78_1527 ();
 sg13g2_decap_4 FILLER_78_1559 ();
 sg13g2_decap_8 FILLER_78_1598 ();
 sg13g2_decap_4 FILLER_78_1605 ();
 sg13g2_fill_2 FILLER_78_1661 ();
 sg13g2_fill_1 FILLER_78_1663 ();
 sg13g2_decap_8 FILLER_78_1669 ();
 sg13g2_fill_1 FILLER_78_1685 ();
 sg13g2_fill_2 FILLER_78_1690 ();
 sg13g2_fill_2 FILLER_78_1731 ();
 sg13g2_fill_1 FILLER_78_1733 ();
 sg13g2_fill_2 FILLER_78_1791 ();
 sg13g2_fill_1 FILLER_78_1793 ();
 sg13g2_decap_4 FILLER_78_1861 ();
 sg13g2_decap_4 FILLER_78_1894 ();
 sg13g2_fill_2 FILLER_78_1929 ();
 sg13g2_fill_1 FILLER_78_1931 ();
 sg13g2_decap_8 FILLER_78_1936 ();
 sg13g2_decap_4 FILLER_78_1943 ();
 sg13g2_fill_1 FILLER_78_1952 ();
 sg13g2_fill_2 FILLER_78_1988 ();
 sg13g2_decap_8 FILLER_78_2016 ();
 sg13g2_decap_4 FILLER_78_2023 ();
 sg13g2_decap_4 FILLER_78_2061 ();
 sg13g2_fill_1 FILLER_78_2065 ();
 sg13g2_decap_8 FILLER_78_2069 ();
 sg13g2_decap_8 FILLER_78_2076 ();
 sg13g2_decap_4 FILLER_78_2083 ();
 sg13g2_decap_8 FILLER_78_2123 ();
 sg13g2_decap_4 FILLER_78_2130 ();
 sg13g2_fill_1 FILLER_78_2134 ();
 sg13g2_fill_2 FILLER_78_2169 ();
 sg13g2_fill_1 FILLER_78_2171 ();
 sg13g2_fill_1 FILLER_78_2177 ();
 sg13g2_fill_2 FILLER_78_2191 ();
 sg13g2_decap_4 FILLER_78_2201 ();
 sg13g2_fill_2 FILLER_78_2210 ();
 sg13g2_fill_1 FILLER_78_2212 ();
 sg13g2_fill_2 FILLER_78_2247 ();
 sg13g2_decap_4 FILLER_78_2254 ();
 sg13g2_fill_1 FILLER_78_2258 ();
 sg13g2_fill_1 FILLER_78_2268 ();
 sg13g2_fill_1 FILLER_78_2273 ();
 sg13g2_fill_2 FILLER_78_2313 ();
 sg13g2_decap_8 FILLER_78_2341 ();
 sg13g2_decap_8 FILLER_78_2348 ();
 sg13g2_decap_8 FILLER_78_2355 ();
 sg13g2_decap_4 FILLER_78_2362 ();
 sg13g2_fill_1 FILLER_78_2366 ();
 sg13g2_fill_2 FILLER_78_2423 ();
 sg13g2_decap_8 FILLER_78_2451 ();
 sg13g2_decap_8 FILLER_78_2458 ();
 sg13g2_decap_8 FILLER_78_2465 ();
 sg13g2_decap_8 FILLER_78_2472 ();
 sg13g2_decap_8 FILLER_78_2479 ();
 sg13g2_decap_8 FILLER_78_2486 ();
 sg13g2_decap_8 FILLER_78_2493 ();
 sg13g2_decap_8 FILLER_78_2500 ();
 sg13g2_decap_8 FILLER_78_2507 ();
 sg13g2_decap_8 FILLER_78_2514 ();
 sg13g2_decap_8 FILLER_78_2521 ();
 sg13g2_decap_8 FILLER_78_2528 ();
 sg13g2_decap_8 FILLER_78_2535 ();
 sg13g2_decap_8 FILLER_78_2542 ();
 sg13g2_decap_8 FILLER_78_2549 ();
 sg13g2_decap_8 FILLER_78_2556 ();
 sg13g2_decap_8 FILLER_78_2563 ();
 sg13g2_decap_8 FILLER_78_2570 ();
 sg13g2_decap_8 FILLER_78_2577 ();
 sg13g2_decap_8 FILLER_78_2584 ();
 sg13g2_decap_8 FILLER_78_2591 ();
 sg13g2_decap_8 FILLER_78_2598 ();
 sg13g2_decap_8 FILLER_78_2605 ();
 sg13g2_decap_8 FILLER_78_2612 ();
 sg13g2_decap_8 FILLER_78_2619 ();
 sg13g2_decap_8 FILLER_78_2626 ();
 sg13g2_decap_8 FILLER_78_2633 ();
 sg13g2_decap_8 FILLER_78_2640 ();
 sg13g2_decap_8 FILLER_78_2647 ();
 sg13g2_decap_8 FILLER_78_2654 ();
 sg13g2_decap_8 FILLER_78_2661 ();
 sg13g2_fill_2 FILLER_78_2668 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_fill_2 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_86 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_4 FILLER_79_165 ();
 sg13g2_fill_1 FILLER_79_177 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_4 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_219 ();
 sg13g2_fill_2 FILLER_79_226 ();
 sg13g2_fill_2 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_307 ();
 sg13g2_decap_4 FILLER_79_339 ();
 sg13g2_fill_2 FILLER_79_343 ();
 sg13g2_fill_2 FILLER_79_371 ();
 sg13g2_fill_1 FILLER_79_380 ();
 sg13g2_fill_1 FILLER_79_386 ();
 sg13g2_fill_1 FILLER_79_395 ();
 sg13g2_decap_4 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_486 ();
 sg13g2_decap_8 FILLER_79_493 ();
 sg13g2_decap_4 FILLER_79_500 ();
 sg13g2_fill_1 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_531 ();
 sg13g2_fill_1 FILLER_79_538 ();
 sg13g2_decap_8 FILLER_79_547 ();
 sg13g2_fill_1 FILLER_79_554 ();
 sg13g2_fill_1 FILLER_79_581 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_4 FILLER_79_613 ();
 sg13g2_fill_2 FILLER_79_617 ();
 sg13g2_decap_4 FILLER_79_645 ();
 sg13g2_fill_2 FILLER_79_653 ();
 sg13g2_decap_8 FILLER_79_663 ();
 sg13g2_decap_8 FILLER_79_670 ();
 sg13g2_fill_2 FILLER_79_681 ();
 sg13g2_fill_2 FILLER_79_709 ();
 sg13g2_fill_1 FILLER_79_711 ();
 sg13g2_fill_2 FILLER_79_738 ();
 sg13g2_fill_1 FILLER_79_740 ();
 sg13g2_decap_4 FILLER_79_780 ();
 sg13g2_fill_1 FILLER_79_814 ();
 sg13g2_fill_2 FILLER_79_901 ();
 sg13g2_fill_2 FILLER_79_942 ();
 sg13g2_fill_1 FILLER_79_944 ();
 sg13g2_fill_2 FILLER_79_971 ();
 sg13g2_fill_1 FILLER_79_973 ();
 sg13g2_decap_8 FILLER_79_978 ();
 sg13g2_decap_8 FILLER_79_985 ();
 sg13g2_decap_4 FILLER_79_992 ();
 sg13g2_decap_8 FILLER_79_1000 ();
 sg13g2_decap_4 FILLER_79_1007 ();
 sg13g2_fill_1 FILLER_79_1011 ();
 sg13g2_fill_2 FILLER_79_1038 ();
 sg13g2_fill_1 FILLER_79_1040 ();
 sg13g2_fill_1 FILLER_79_1059 ();
 sg13g2_fill_1 FILLER_79_1090 ();
 sg13g2_fill_1 FILLER_79_1143 ();
 sg13g2_decap_4 FILLER_79_1174 ();
 sg13g2_fill_1 FILLER_79_1178 ();
 sg13g2_decap_4 FILLER_79_1252 ();
 sg13g2_fill_2 FILLER_79_1256 ();
 sg13g2_decap_8 FILLER_79_1292 ();
 sg13g2_decap_4 FILLER_79_1299 ();
 sg13g2_fill_2 FILLER_79_1354 ();
 sg13g2_fill_1 FILLER_79_1382 ();
 sg13g2_fill_2 FILLER_79_1391 ();
 sg13g2_decap_8 FILLER_79_1419 ();
 sg13g2_decap_4 FILLER_79_1426 ();
 sg13g2_fill_1 FILLER_79_1430 ();
 sg13g2_fill_2 FILLER_79_1486 ();
 sg13g2_fill_1 FILLER_79_1488 ();
 sg13g2_fill_1 FILLER_79_1515 ();
 sg13g2_decap_8 FILLER_79_1546 ();
 sg13g2_fill_1 FILLER_79_1571 ();
 sg13g2_decap_8 FILLER_79_1598 ();
 sg13g2_fill_1 FILLER_79_1610 ();
 sg13g2_fill_2 FILLER_79_1659 ();
 sg13g2_fill_2 FILLER_79_1713 ();
 sg13g2_fill_2 FILLER_79_1741 ();
 sg13g2_fill_2 FILLER_79_1769 ();
 sg13g2_fill_1 FILLER_79_1771 ();
 sg13g2_decap_4 FILLER_79_1777 ();
 sg13g2_fill_1 FILLER_79_1781 ();
 sg13g2_decap_4 FILLER_79_1808 ();
 sg13g2_fill_2 FILLER_79_1812 ();
 sg13g2_fill_2 FILLER_79_1818 ();
 sg13g2_decap_8 FILLER_79_1824 ();
 sg13g2_decap_8 FILLER_79_1831 ();
 sg13g2_decap_8 FILLER_79_1842 ();
 sg13g2_decap_4 FILLER_79_1849 ();
 sg13g2_fill_2 FILLER_79_1863 ();
 sg13g2_decap_4 FILLER_79_1901 ();
 sg13g2_fill_1 FILLER_79_1905 ();
 sg13g2_fill_2 FILLER_79_1911 ();
 sg13g2_fill_1 FILLER_79_1913 ();
 sg13g2_decap_4 FILLER_79_1918 ();
 sg13g2_fill_1 FILLER_79_1922 ();
 sg13g2_decap_8 FILLER_79_1949 ();
 sg13g2_decap_8 FILLER_79_1956 ();
 sg13g2_fill_2 FILLER_79_1963 ();
 sg13g2_decap_4 FILLER_79_1970 ();
 sg13g2_fill_1 FILLER_79_1974 ();
 sg13g2_decap_8 FILLER_79_1979 ();
 sg13g2_decap_8 FILLER_79_1986 ();
 sg13g2_decap_4 FILLER_79_1993 ();
 sg13g2_fill_1 FILLER_79_1997 ();
 sg13g2_decap_8 FILLER_79_2028 ();
 sg13g2_decap_8 FILLER_79_2035 ();
 sg13g2_decap_8 FILLER_79_2042 ();
 sg13g2_decap_8 FILLER_79_2049 ();
 sg13g2_decap_4 FILLER_79_2056 ();
 sg13g2_fill_1 FILLER_79_2065 ();
 sg13g2_fill_2 FILLER_79_2071 ();
 sg13g2_decap_8 FILLER_79_2099 ();
 sg13g2_decap_8 FILLER_79_2106 ();
 sg13g2_decap_4 FILLER_79_2113 ();
 sg13g2_decap_8 FILLER_79_2144 ();
 sg13g2_fill_2 FILLER_79_2156 ();
 sg13g2_fill_2 FILLER_79_2188 ();
 sg13g2_decap_4 FILLER_79_2195 ();
 sg13g2_decap_4 FILLER_79_2225 ();
 sg13g2_fill_2 FILLER_79_2234 ();
 sg13g2_fill_1 FILLER_79_2262 ();
 sg13g2_decap_8 FILLER_79_2289 ();
 sg13g2_fill_2 FILLER_79_2296 ();
 sg13g2_fill_1 FILLER_79_2298 ();
 sg13g2_decap_4 FILLER_79_2307 ();
 sg13g2_fill_1 FILLER_79_2311 ();
 sg13g2_decap_8 FILLER_79_2346 ();
 sg13g2_decap_8 FILLER_79_2353 ();
 sg13g2_decap_8 FILLER_79_2360 ();
 sg13g2_decap_8 FILLER_79_2367 ();
 sg13g2_decap_4 FILLER_79_2374 ();
 sg13g2_decap_4 FILLER_79_2386 ();
 sg13g2_fill_2 FILLER_79_2420 ();
 sg13g2_decap_8 FILLER_79_2448 ();
 sg13g2_decap_8 FILLER_79_2455 ();
 sg13g2_decap_8 FILLER_79_2462 ();
 sg13g2_decap_8 FILLER_79_2469 ();
 sg13g2_decap_8 FILLER_79_2476 ();
 sg13g2_decap_8 FILLER_79_2483 ();
 sg13g2_decap_8 FILLER_79_2490 ();
 sg13g2_decap_8 FILLER_79_2497 ();
 sg13g2_decap_8 FILLER_79_2504 ();
 sg13g2_decap_8 FILLER_79_2511 ();
 sg13g2_decap_8 FILLER_79_2518 ();
 sg13g2_decap_8 FILLER_79_2525 ();
 sg13g2_decap_8 FILLER_79_2532 ();
 sg13g2_decap_8 FILLER_79_2539 ();
 sg13g2_decap_8 FILLER_79_2546 ();
 sg13g2_decap_8 FILLER_79_2553 ();
 sg13g2_decap_8 FILLER_79_2560 ();
 sg13g2_decap_8 FILLER_79_2567 ();
 sg13g2_decap_8 FILLER_79_2574 ();
 sg13g2_decap_8 FILLER_79_2581 ();
 sg13g2_decap_8 FILLER_79_2588 ();
 sg13g2_decap_8 FILLER_79_2595 ();
 sg13g2_decap_8 FILLER_79_2602 ();
 sg13g2_decap_8 FILLER_79_2609 ();
 sg13g2_decap_8 FILLER_79_2616 ();
 sg13g2_decap_8 FILLER_79_2623 ();
 sg13g2_decap_8 FILLER_79_2630 ();
 sg13g2_decap_8 FILLER_79_2637 ();
 sg13g2_decap_8 FILLER_79_2644 ();
 sg13g2_decap_8 FILLER_79_2651 ();
 sg13g2_decap_8 FILLER_79_2658 ();
 sg13g2_decap_4 FILLER_79_2665 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_1 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_2 FILLER_80_88 ();
 sg13g2_fill_1 FILLER_80_94 ();
 sg13g2_fill_2 FILLER_80_115 ();
 sg13g2_fill_2 FILLER_80_129 ();
 sg13g2_decap_8 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_146 ();
 sg13g2_decap_8 FILLER_80_153 ();
 sg13g2_decap_8 FILLER_80_172 ();
 sg13g2_fill_1 FILLER_80_179 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_fill_2 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_fill_1 FILLER_80_237 ();
 sg13g2_decap_4 FILLER_80_250 ();
 sg13g2_fill_1 FILLER_80_254 ();
 sg13g2_fill_1 FILLER_80_259 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_275 ();
 sg13g2_decap_8 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_decap_8 FILLER_80_317 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_fill_2 FILLER_80_328 ();
 sg13g2_fill_2 FILLER_80_334 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_fill_1 FILLER_80_354 ();
 sg13g2_decap_4 FILLER_80_359 ();
 sg13g2_fill_1 FILLER_80_363 ();
 sg13g2_fill_1 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_8 FILLER_80_404 ();
 sg13g2_decap_8 FILLER_80_411 ();
 sg13g2_decap_8 FILLER_80_418 ();
 sg13g2_decap_8 FILLER_80_425 ();
 sg13g2_fill_2 FILLER_80_432 ();
 sg13g2_fill_1 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_708 ();
 sg13g2_decap_4 FILLER_80_715 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_fill_1 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_fill_2 FILLER_80_767 ();
 sg13g2_fill_1 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_fill_1 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_4 FILLER_80_821 ();
 sg13g2_fill_2 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_fill_1 FILLER_80_852 ();
 sg13g2_decap_8 FILLER_80_865 ();
 sg13g2_decap_4 FILLER_80_872 ();
 sg13g2_fill_2 FILLER_80_876 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_fill_2 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_913 ();
 sg13g2_decap_8 FILLER_80_920 ();
 sg13g2_decap_4 FILLER_80_927 ();
 sg13g2_fill_2 FILLER_80_935 ();
 sg13g2_fill_1 FILLER_80_937 ();
 sg13g2_fill_2 FILLER_80_942 ();
 sg13g2_decap_4 FILLER_80_948 ();
 sg13g2_fill_2 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_958 ();
 sg13g2_decap_8 FILLER_80_965 ();
 sg13g2_decap_8 FILLER_80_972 ();
 sg13g2_decap_8 FILLER_80_979 ();
 sg13g2_decap_4 FILLER_80_986 ();
 sg13g2_decap_4 FILLER_80_1032 ();
 sg13g2_fill_2 FILLER_80_1036 ();
 sg13g2_decap_8 FILLER_80_1042 ();
 sg13g2_fill_1 FILLER_80_1049 ();
 sg13g2_decap_8 FILLER_80_1054 ();
 sg13g2_fill_2 FILLER_80_1061 ();
 sg13g2_fill_1 FILLER_80_1063 ();
 sg13g2_decap_8 FILLER_80_1072 ();
 sg13g2_decap_8 FILLER_80_1079 ();
 sg13g2_decap_8 FILLER_80_1086 ();
 sg13g2_decap_8 FILLER_80_1093 ();
 sg13g2_decap_8 FILLER_80_1100 ();
 sg13g2_decap_8 FILLER_80_1107 ();
 sg13g2_decap_8 FILLER_80_1114 ();
 sg13g2_decap_8 FILLER_80_1121 ();
 sg13g2_decap_4 FILLER_80_1128 ();
 sg13g2_fill_2 FILLER_80_1132 ();
 sg13g2_decap_8 FILLER_80_1139 ();
 sg13g2_fill_2 FILLER_80_1146 ();
 sg13g2_fill_1 FILLER_80_1148 ();
 sg13g2_decap_4 FILLER_80_1157 ();
 sg13g2_decap_8 FILLER_80_1165 ();
 sg13g2_decap_8 FILLER_80_1172 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_4 FILLER_80_1186 ();
 sg13g2_fill_2 FILLER_80_1190 ();
 sg13g2_decap_8 FILLER_80_1196 ();
 sg13g2_decap_4 FILLER_80_1233 ();
 sg13g2_fill_2 FILLER_80_1237 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_fill_2 FILLER_80_1250 ();
 sg13g2_fill_1 FILLER_80_1252 ();
 sg13g2_decap_8 FILLER_80_1283 ();
 sg13g2_decap_8 FILLER_80_1290 ();
 sg13g2_decap_8 FILLER_80_1297 ();
 sg13g2_decap_8 FILLER_80_1304 ();
 sg13g2_fill_2 FILLER_80_1315 ();
 sg13g2_fill_1 FILLER_80_1317 ();
 sg13g2_decap_8 FILLER_80_1322 ();
 sg13g2_decap_8 FILLER_80_1329 ();
 sg13g2_fill_1 FILLER_80_1336 ();
 sg13g2_decap_4 FILLER_80_1341 ();
 sg13g2_decap_8 FILLER_80_1349 ();
 sg13g2_decap_8 FILLER_80_1356 ();
 sg13g2_decap_8 FILLER_80_1367 ();
 sg13g2_decap_8 FILLER_80_1374 ();
 sg13g2_decap_8 FILLER_80_1381 ();
 sg13g2_fill_1 FILLER_80_1388 ();
 sg13g2_fill_1 FILLER_80_1393 ();
 sg13g2_decap_8 FILLER_80_1398 ();
 sg13g2_decap_8 FILLER_80_1405 ();
 sg13g2_decap_8 FILLER_80_1412 ();
 sg13g2_decap_8 FILLER_80_1419 ();
 sg13g2_decap_8 FILLER_80_1426 ();
 sg13g2_decap_8 FILLER_80_1433 ();
 sg13g2_decap_8 FILLER_80_1444 ();
 sg13g2_decap_8 FILLER_80_1451 ();
 sg13g2_decap_8 FILLER_80_1458 ();
 sg13g2_fill_1 FILLER_80_1465 ();
 sg13g2_decap_4 FILLER_80_1478 ();
 sg13g2_fill_1 FILLER_80_1482 ();
 sg13g2_decap_8 FILLER_80_1488 ();
 sg13g2_decap_8 FILLER_80_1495 ();
 sg13g2_decap_8 FILLER_80_1502 ();
 sg13g2_decap_8 FILLER_80_1509 ();
 sg13g2_decap_8 FILLER_80_1516 ();
 sg13g2_fill_1 FILLER_80_1523 ();
 sg13g2_decap_8 FILLER_80_1528 ();
 sg13g2_decap_8 FILLER_80_1535 ();
 sg13g2_decap_8 FILLER_80_1542 ();
 sg13g2_decap_8 FILLER_80_1549 ();
 sg13g2_fill_1 FILLER_80_1556 ();
 sg13g2_decap_4 FILLER_80_1561 ();
 sg13g2_fill_2 FILLER_80_1565 ();
 sg13g2_fill_2 FILLER_80_1571 ();
 sg13g2_fill_1 FILLER_80_1573 ();
 sg13g2_decap_8 FILLER_80_1582 ();
 sg13g2_decap_8 FILLER_80_1589 ();
 sg13g2_decap_8 FILLER_80_1596 ();
 sg13g2_decap_8 FILLER_80_1603 ();
 sg13g2_decap_8 FILLER_80_1610 ();
 sg13g2_decap_8 FILLER_80_1617 ();
 sg13g2_decap_8 FILLER_80_1624 ();
 sg13g2_decap_8 FILLER_80_1631 ();
 sg13g2_decap_8 FILLER_80_1638 ();
 sg13g2_decap_8 FILLER_80_1645 ();
 sg13g2_fill_2 FILLER_80_1652 ();
 sg13g2_decap_8 FILLER_80_1659 ();
 sg13g2_decap_8 FILLER_80_1666 ();
 sg13g2_decap_8 FILLER_80_1673 ();
 sg13g2_decap_8 FILLER_80_1680 ();
 sg13g2_decap_8 FILLER_80_1687 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_decap_4 FILLER_80_1701 ();
 sg13g2_fill_1 FILLER_80_1705 ();
 sg13g2_decap_4 FILLER_80_1711 ();
 sg13g2_fill_1 FILLER_80_1715 ();
 sg13g2_decap_8 FILLER_80_1724 ();
 sg13g2_decap_8 FILLER_80_1731 ();
 sg13g2_decap_4 FILLER_80_1738 ();
 sg13g2_fill_1 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 sg13g2_decap_8 FILLER_80_1768 ();
 sg13g2_decap_8 FILLER_80_1775 ();
 sg13g2_decap_8 FILLER_80_1782 ();
 sg13g2_decap_8 FILLER_80_1789 ();
 sg13g2_decap_8 FILLER_80_1796 ();
 sg13g2_decap_8 FILLER_80_1803 ();
 sg13g2_decap_8 FILLER_80_1810 ();
 sg13g2_decap_8 FILLER_80_1817 ();
 sg13g2_decap_8 FILLER_80_1824 ();
 sg13g2_decap_8 FILLER_80_1831 ();
 sg13g2_decap_8 FILLER_80_1838 ();
 sg13g2_decap_8 FILLER_80_1845 ();
 sg13g2_fill_1 FILLER_80_1852 ();
 sg13g2_fill_1 FILLER_80_1866 ();
 sg13g2_decap_8 FILLER_80_1889 ();
 sg13g2_decap_8 FILLER_80_1896 ();
 sg13g2_decap_8 FILLER_80_1903 ();
 sg13g2_decap_8 FILLER_80_1910 ();
 sg13g2_decap_8 FILLER_80_1925 ();
 sg13g2_decap_8 FILLER_80_1932 ();
 sg13g2_decap_8 FILLER_80_1939 ();
 sg13g2_decap_8 FILLER_80_1946 ();
 sg13g2_decap_8 FILLER_80_1953 ();
 sg13g2_decap_8 FILLER_80_1960 ();
 sg13g2_decap_4 FILLER_80_1967 ();
 sg13g2_fill_2 FILLER_80_1971 ();
 sg13g2_fill_2 FILLER_80_1999 ();
 sg13g2_decap_4 FILLER_80_2019 ();
 sg13g2_fill_1 FILLER_80_2023 ();
 sg13g2_decap_8 FILLER_80_2032 ();
 sg13g2_decap_8 FILLER_80_2039 ();
 sg13g2_decap_8 FILLER_80_2046 ();
 sg13g2_decap_8 FILLER_80_2053 ();
 sg13g2_decap_8 FILLER_80_2060 ();
 sg13g2_decap_8 FILLER_80_2067 ();
 sg13g2_decap_8 FILLER_80_2074 ();
 sg13g2_decap_8 FILLER_80_2081 ();
 sg13g2_decap_8 FILLER_80_2088 ();
 sg13g2_decap_8 FILLER_80_2095 ();
 sg13g2_decap_8 FILLER_80_2102 ();
 sg13g2_decap_8 FILLER_80_2109 ();
 sg13g2_decap_8 FILLER_80_2116 ();
 sg13g2_decap_8 FILLER_80_2123 ();
 sg13g2_decap_8 FILLER_80_2130 ();
 sg13g2_decap_8 FILLER_80_2137 ();
 sg13g2_decap_8 FILLER_80_2144 ();
 sg13g2_decap_8 FILLER_80_2151 ();
 sg13g2_fill_2 FILLER_80_2158 ();
 sg13g2_decap_8 FILLER_80_2168 ();
 sg13g2_decap_8 FILLER_80_2175 ();
 sg13g2_decap_8 FILLER_80_2182 ();
 sg13g2_decap_4 FILLER_80_2189 ();
 sg13g2_fill_2 FILLER_80_2193 ();
 sg13g2_decap_8 FILLER_80_2200 ();
 sg13g2_decap_8 FILLER_80_2207 ();
 sg13g2_decap_8 FILLER_80_2214 ();
 sg13g2_decap_8 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2228 ();
 sg13g2_fill_1 FILLER_80_2235 ();
 sg13g2_decap_8 FILLER_80_2241 ();
 sg13g2_decap_8 FILLER_80_2248 ();
 sg13g2_decap_8 FILLER_80_2255 ();
 sg13g2_decap_8 FILLER_80_2262 ();
 sg13g2_decap_8 FILLER_80_2269 ();
 sg13g2_decap_8 FILLER_80_2276 ();
 sg13g2_decap_8 FILLER_80_2283 ();
 sg13g2_decap_8 FILLER_80_2290 ();
 sg13g2_decap_8 FILLER_80_2297 ();
 sg13g2_decap_8 FILLER_80_2304 ();
 sg13g2_decap_8 FILLER_80_2311 ();
 sg13g2_decap_8 FILLER_80_2318 ();
 sg13g2_decap_8 FILLER_80_2325 ();
 sg13g2_decap_8 FILLER_80_2332 ();
 sg13g2_decap_8 FILLER_80_2339 ();
 sg13g2_decap_8 FILLER_80_2346 ();
 sg13g2_decap_8 FILLER_80_2353 ();
 sg13g2_decap_8 FILLER_80_2360 ();
 sg13g2_decap_8 FILLER_80_2367 ();
 sg13g2_decap_8 FILLER_80_2374 ();
 sg13g2_decap_8 FILLER_80_2381 ();
 sg13g2_decap_8 FILLER_80_2388 ();
 sg13g2_decap_4 FILLER_80_2399 ();
 sg13g2_fill_2 FILLER_80_2403 ();
 sg13g2_decap_8 FILLER_80_2409 ();
 sg13g2_decap_8 FILLER_80_2416 ();
 sg13g2_fill_2 FILLER_80_2423 ();
 sg13g2_fill_1 FILLER_80_2425 ();
 sg13g2_fill_2 FILLER_80_2430 ();
 sg13g2_fill_1 FILLER_80_2432 ();
 sg13g2_decap_8 FILLER_80_2437 ();
 sg13g2_decap_8 FILLER_80_2444 ();
 sg13g2_decap_8 FILLER_80_2451 ();
 sg13g2_decap_8 FILLER_80_2458 ();
 sg13g2_decap_8 FILLER_80_2465 ();
 sg13g2_decap_8 FILLER_80_2472 ();
 sg13g2_decap_8 FILLER_80_2479 ();
 sg13g2_decap_8 FILLER_80_2486 ();
 sg13g2_decap_8 FILLER_80_2493 ();
 sg13g2_decap_8 FILLER_80_2500 ();
 sg13g2_decap_8 FILLER_80_2507 ();
 sg13g2_decap_8 FILLER_80_2514 ();
 sg13g2_decap_8 FILLER_80_2521 ();
 sg13g2_decap_8 FILLER_80_2528 ();
 sg13g2_decap_8 FILLER_80_2535 ();
 sg13g2_decap_8 FILLER_80_2542 ();
 sg13g2_decap_8 FILLER_80_2549 ();
 sg13g2_decap_8 FILLER_80_2556 ();
 sg13g2_decap_8 FILLER_80_2563 ();
 sg13g2_decap_8 FILLER_80_2570 ();
 sg13g2_decap_8 FILLER_80_2577 ();
 sg13g2_decap_8 FILLER_80_2584 ();
 sg13g2_decap_8 FILLER_80_2591 ();
 sg13g2_decap_8 FILLER_80_2598 ();
 sg13g2_decap_8 FILLER_80_2605 ();
 sg13g2_decap_8 FILLER_80_2612 ();
 sg13g2_decap_8 FILLER_80_2619 ();
 sg13g2_decap_8 FILLER_80_2626 ();
 sg13g2_decap_8 FILLER_80_2633 ();
 sg13g2_decap_8 FILLER_80_2640 ();
 sg13g2_decap_8 FILLER_80_2647 ();
 sg13g2_decap_8 FILLER_80_2654 ();
 sg13g2_decap_8 FILLER_80_2661 ();
 sg13g2_fill_2 FILLER_80_2668 ();
endmodule
