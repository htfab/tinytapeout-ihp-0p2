module tt_um_multi_bit_puf_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire clknet_0_clk;
 wire net108;
 wire \puf_instance.puf_loop[0].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[0].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[100].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[100].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[101].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[101].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[102].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[102].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[103].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[103].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[104].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[104].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[105].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[105].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[106].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[106].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[107].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[107].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[108].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[108].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[109].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[109].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[10].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[10].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[110].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[110].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[111].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[111].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[112].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[112].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[113].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[113].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[114].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[114].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[115].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[115].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[116].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[116].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[117].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[117].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[118].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[118].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[119].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[119].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[11].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[11].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[120].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[120].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[121].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[121].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[122].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[122].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[123].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[123].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[124].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[124].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[125].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[125].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[126].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[126].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[127].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[127].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[12].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[12].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[13].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[13].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[14].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[14].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[15].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[15].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[16].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[16].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[17].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[17].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[18].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[18].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[19].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[19].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[1].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[1].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[20].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[20].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[21].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[21].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[22].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[22].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[23].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[23].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[24].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[24].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[25].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[25].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[26].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[26].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[27].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[27].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[28].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[28].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[29].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[29].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[2].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[2].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[30].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[30].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[31].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[31].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[32].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[32].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[33].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[33].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[34].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[34].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[35].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[35].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[36].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[36].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[37].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[37].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[38].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[38].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[39].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[39].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[3].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[3].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[40].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[40].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[41].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[41].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[42].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[42].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[43].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[43].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[44].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[44].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[45].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[45].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[46].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[46].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[47].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[47].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[48].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[48].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[49].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[49].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[4].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[4].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[50].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[50].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[51].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[51].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[52].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[52].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[53].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[53].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[54].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[54].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[55].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[55].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[56].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[56].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[57].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[57].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[58].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[58].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[59].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[59].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[5].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[5].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[60].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[60].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[61].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[61].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[62].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[62].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[63].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[63].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[64].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[64].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[65].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[65].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[66].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[66].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[67].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[67].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[68].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[68].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[69].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[69].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[6].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[6].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[70].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[70].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[71].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[71].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[72].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[72].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[73].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[73].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[74].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[74].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[75].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[75].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[76].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[76].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[77].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[77].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[78].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[78].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[79].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[79].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[7].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[7].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[80].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[80].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[81].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[81].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[82].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[82].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[83].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[83].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[84].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[84].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[85].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[85].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[86].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[86].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[87].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[87].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[88].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[88].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[89].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[89].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[8].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[8].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[90].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[90].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[91].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[91].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[92].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[92].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[93].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[93].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[94].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[94].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[95].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[95].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[96].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[96].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[97].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[97].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[98].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[98].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[99].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[99].puf_inst.Q1 ;
 wire \puf_instance.puf_loop[9].puf_inst.Q0 ;
 wire \puf_instance.puf_loop[9].puf_inst.Q1 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sg13g2_buf_8 _367_ (.A(ui_in[1]),
    .X(_265_));
 sg13g2_buf_8 _368_ (.A(_265_),
    .X(_266_));
 sg13g2_buf_8 _369_ (.A(ui_in[0]),
    .X(_267_));
 sg13g2_buf_1 _370_ (.A(_267_),
    .X(_268_));
 sg13g2_mux4_1 _371_ (.S0(net90),
    .A0(\puf_instance.puf_loop[64].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[80].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[72].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[88].puf_inst.Q1 ),
    .S1(net89),
    .X(_269_));
 sg13g2_nor2b_1 _372_ (.A(net2),
    .B_N(net3),
    .Y(_270_));
 sg13g2_buf_2 _373_ (.A(_270_),
    .X(_271_));
 sg13g2_buf_8 _374_ (.A(_267_),
    .X(_272_));
 sg13g2_buf_1 _375_ (.A(_265_),
    .X(_273_));
 sg13g2_mux4_1 _376_ (.S0(net88),
    .A0(\puf_instance.puf_loop[96].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[104].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[112].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[120].puf_inst.Q1 ),
    .S1(net87),
    .X(_274_));
 sg13g2_and2_1 _377_ (.A(net2),
    .B(net3),
    .X(_275_));
 sg13g2_buf_2 _378_ (.A(_275_),
    .X(_276_));
 sg13g2_a22oi_1 _379_ (.Y(_277_),
    .B1(_274_),
    .B2(_276_),
    .A2(_271_),
    .A1(_269_));
 sg13g2_mux4_1 _380_ (.S0(net90),
    .A0(\puf_instance.puf_loop[0].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[16].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[8].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[24].puf_inst.Q1 ),
    .S1(net89),
    .X(_278_));
 sg13g2_nor2_2 _381_ (.A(net2),
    .B(net3),
    .Y(_279_));
 sg13g2_buf_8 _382_ (.A(_265_),
    .X(_280_));
 sg13g2_buf_1 _383_ (.A(_267_),
    .X(_281_));
 sg13g2_mux4_1 _384_ (.S0(net86),
    .A0(\puf_instance.puf_loop[32].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[48].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[40].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[56].puf_inst.Q1 ),
    .S1(net85),
    .X(_282_));
 sg13g2_nor2b_1 _385_ (.A(net3),
    .B_N(net2),
    .Y(_283_));
 sg13g2_buf_2 _386_ (.A(_283_),
    .X(_284_));
 sg13g2_a22oi_1 _387_ (.Y(_285_),
    .B1(_282_),
    .B2(_284_),
    .A2(_279_),
    .A1(_278_));
 sg13g2_and2_1 _388_ (.A(_277_),
    .B(_285_),
    .X(_257_));
 sg13g2_mux4_1 _389_ (.S0(_266_),
    .A0(\puf_instance.puf_loop[65].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[81].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[73].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[89].puf_inst.Q1 ),
    .S1(_268_),
    .X(_286_));
 sg13g2_mux4_1 _390_ (.S0(net88),
    .A0(\puf_instance.puf_loop[97].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[105].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[113].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[121].puf_inst.Q1 ),
    .S1(net87),
    .X(_287_));
 sg13g2_a22oi_1 _391_ (.Y(_288_),
    .B1(_287_),
    .B2(_276_),
    .A2(_286_),
    .A1(_271_));
 sg13g2_mux4_1 _392_ (.S0(_265_),
    .A0(\puf_instance.puf_loop[1].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[17].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[9].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[25].puf_inst.Q1 ),
    .S1(net88),
    .X(_289_));
 sg13g2_mux4_1 _393_ (.S0(net86),
    .A0(\puf_instance.puf_loop[33].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[49].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[41].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[57].puf_inst.Q1 ),
    .S1(net85),
    .X(_290_));
 sg13g2_a22oi_1 _394_ (.Y(_291_),
    .B1(_290_),
    .B2(_284_),
    .A2(_289_),
    .A1(_279_));
 sg13g2_and2_1 _395_ (.A(_288_),
    .B(_291_),
    .X(_258_));
 sg13g2_mux4_1 _396_ (.S0(_266_),
    .A0(\puf_instance.puf_loop[66].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[82].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[74].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[90].puf_inst.Q1 ),
    .S1(_268_),
    .X(_292_));
 sg13g2_mux4_1 _397_ (.S0(net88),
    .A0(\puf_instance.puf_loop[98].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[106].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[114].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[122].puf_inst.Q1 ),
    .S1(net87),
    .X(_293_));
 sg13g2_a22oi_1 _398_ (.Y(_294_),
    .B1(_293_),
    .B2(_276_),
    .A2(_292_),
    .A1(_271_));
 sg13g2_mux4_1 _399_ (.S0(net88),
    .A0(\puf_instance.puf_loop[2].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[10].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[18].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[26].puf_inst.Q1 ),
    .S1(net87),
    .X(_295_));
 sg13g2_mux4_1 _400_ (.S0(net86),
    .A0(\puf_instance.puf_loop[34].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[50].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[42].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[58].puf_inst.Q1 ),
    .S1(net85),
    .X(_296_));
 sg13g2_a22oi_1 _401_ (.Y(_297_),
    .B1(_296_),
    .B2(_284_),
    .A2(_295_),
    .A1(_279_));
 sg13g2_and2_1 _402_ (.A(_294_),
    .B(_297_),
    .X(_259_));
 sg13g2_mux4_1 _403_ (.S0(net90),
    .A0(\puf_instance.puf_loop[67].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[83].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[75].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[91].puf_inst.Q1 ),
    .S1(net89),
    .X(_298_));
 sg13g2_mux4_1 _404_ (.S0(net88),
    .A0(\puf_instance.puf_loop[99].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[107].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[115].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[123].puf_inst.Q1 ),
    .S1(net87),
    .X(_299_));
 sg13g2_a22oi_1 _405_ (.Y(_300_),
    .B1(_299_),
    .B2(_276_),
    .A2(_298_),
    .A1(_271_));
 sg13g2_mux4_1 _406_ (.S0(net88),
    .A0(\puf_instance.puf_loop[3].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[11].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[19].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[27].puf_inst.Q1 ),
    .S1(net87),
    .X(_301_));
 sg13g2_mux4_1 _407_ (.S0(net86),
    .A0(\puf_instance.puf_loop[35].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[51].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[43].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[59].puf_inst.Q1 ),
    .S1(net85),
    .X(_302_));
 sg13g2_a22oi_1 _408_ (.Y(_303_),
    .B1(_302_),
    .B2(_284_),
    .A2(_301_),
    .A1(_279_));
 sg13g2_and2_1 _409_ (.A(_300_),
    .B(_303_),
    .X(_260_));
 sg13g2_mux4_1 _410_ (.S0(net90),
    .A0(\puf_instance.puf_loop[68].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[84].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[76].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[92].puf_inst.Q1 ),
    .S1(net89),
    .X(_304_));
 sg13g2_mux4_1 _411_ (.S0(net86),
    .A0(\puf_instance.puf_loop[100].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[116].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[108].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[124].puf_inst.Q1 ),
    .S1(net85),
    .X(_305_));
 sg13g2_a22oi_1 _412_ (.Y(_306_),
    .B1(_305_),
    .B2(_276_),
    .A2(_304_),
    .A1(_271_));
 sg13g2_mux4_1 _413_ (.S0(_272_),
    .A0(\puf_instance.puf_loop[4].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[12].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[20].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[28].puf_inst.Q1 ),
    .S1(_273_),
    .X(_307_));
 sg13g2_mux4_1 _414_ (.S0(net86),
    .A0(\puf_instance.puf_loop[36].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[52].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[44].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[60].puf_inst.Q1 ),
    .S1(net85),
    .X(_308_));
 sg13g2_a22oi_1 _415_ (.Y(_309_),
    .B1(_308_),
    .B2(_284_),
    .A2(_307_),
    .A1(_279_));
 sg13g2_and2_1 _416_ (.A(_306_),
    .B(_309_),
    .X(_261_));
 sg13g2_mux4_1 _417_ (.S0(net90),
    .A0(\puf_instance.puf_loop[69].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[85].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[77].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[93].puf_inst.Q1 ),
    .S1(net89),
    .X(_310_));
 sg13g2_mux4_1 _418_ (.S0(net86),
    .A0(\puf_instance.puf_loop[101].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[117].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[109].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[125].puf_inst.Q1 ),
    .S1(net85),
    .X(_311_));
 sg13g2_a22oi_1 _419_ (.Y(_312_),
    .B1(_311_),
    .B2(_276_),
    .A2(_310_),
    .A1(_271_));
 sg13g2_mux4_1 _420_ (.S0(_272_),
    .A0(\puf_instance.puf_loop[5].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[13].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[21].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[29].puf_inst.Q1 ),
    .S1(_273_),
    .X(_313_));
 sg13g2_mux4_1 _421_ (.S0(net86),
    .A0(\puf_instance.puf_loop[37].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[53].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[45].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[61].puf_inst.Q1 ),
    .S1(net85),
    .X(_314_));
 sg13g2_a22oi_1 _422_ (.Y(_315_),
    .B1(_314_),
    .B2(_284_),
    .A2(_313_),
    .A1(_279_));
 sg13g2_and2_1 _423_ (.A(_312_),
    .B(_315_),
    .X(_262_));
 sg13g2_mux4_1 _424_ (.S0(net90),
    .A0(\puf_instance.puf_loop[70].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[86].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[78].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[94].puf_inst.Q1 ),
    .S1(net89),
    .X(_316_));
 sg13g2_mux4_1 _425_ (.S0(_280_),
    .A0(\puf_instance.puf_loop[102].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[118].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[110].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[126].puf_inst.Q1 ),
    .S1(_281_),
    .X(_317_));
 sg13g2_a22oi_1 _426_ (.Y(_318_),
    .B1(_317_),
    .B2(_276_),
    .A2(_316_),
    .A1(_271_));
 sg13g2_mux4_1 _427_ (.S0(_267_),
    .A0(\puf_instance.puf_loop[6].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[14].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[22].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[30].puf_inst.Q1 ),
    .S1(net87),
    .X(_319_));
 sg13g2_mux4_1 _428_ (.S0(net90),
    .A0(\puf_instance.puf_loop[38].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[54].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[46].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[62].puf_inst.Q1 ),
    .S1(net89),
    .X(_320_));
 sg13g2_a22oi_1 _429_ (.Y(_321_),
    .B1(_320_),
    .B2(_284_),
    .A2(_319_),
    .A1(_279_));
 sg13g2_and2_1 _430_ (.A(_318_),
    .B(_321_),
    .X(_263_));
 sg13g2_mux4_1 _431_ (.S0(_265_),
    .A0(\puf_instance.puf_loop[71].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[87].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[79].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[95].puf_inst.Q1 ),
    .S1(net88),
    .X(_322_));
 sg13g2_mux4_1 _432_ (.S0(_280_),
    .A0(\puf_instance.puf_loop[103].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[119].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[111].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[127].puf_inst.Q1 ),
    .S1(_281_),
    .X(_323_));
 sg13g2_a22oi_1 _433_ (.Y(_324_),
    .B1(_323_),
    .B2(_276_),
    .A2(_322_),
    .A1(_271_));
 sg13g2_mux4_1 _434_ (.S0(_267_),
    .A0(\puf_instance.puf_loop[7].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[15].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[23].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[31].puf_inst.Q1 ),
    .S1(net87),
    .X(_325_));
 sg13g2_mux4_1 _435_ (.S0(net90),
    .A0(\puf_instance.puf_loop[39].puf_inst.Q1 ),
    .A1(\puf_instance.puf_loop[55].puf_inst.Q1 ),
    .A2(\puf_instance.puf_loop[47].puf_inst.Q1 ),
    .A3(\puf_instance.puf_loop[63].puf_inst.Q1 ),
    .S1(net89),
    .X(_326_));
 sg13g2_a22oi_1 _436_ (.Y(_327_),
    .B1(_326_),
    .B2(_284_),
    .A2(_325_),
    .A1(_279_));
 sg13g2_and2_1 _437_ (.A(_324_),
    .B(_327_),
    .X(_264_));
 sg13g2_buf_1 _438_ (.A(net91),
    .X(_328_));
 sg13g2_buf_1 _439_ (.A(_328_),
    .X(_329_));
 sg13g2_buf_1 _440_ (.A(net84),
    .X(_330_));
 sg13g2_nor2b_1 _441_ (.A(\puf_instance.puf_loop[9].puf_inst.Q1 ),
    .B_N(net79),
    .Y(_255_));
 sg13g2_nor2b_1 _442_ (.A(\puf_instance.puf_loop[9].puf_inst.Q0 ),
    .B_N(net79),
    .Y(_256_));
 sg13g2_nor2b_1 _443_ (.A(\puf_instance.puf_loop[99].puf_inst.Q1 ),
    .B_N(_330_),
    .Y(_253_));
 sg13g2_nor2b_1 _444_ (.A(\puf_instance.puf_loop[99].puf_inst.Q0 ),
    .B_N(_330_),
    .Y(_254_));
 sg13g2_nor2b_1 _445_ (.A(\puf_instance.puf_loop[98].puf_inst.Q1 ),
    .B_N(net79),
    .Y(_251_));
 sg13g2_nor2b_1 _446_ (.A(\puf_instance.puf_loop[98].puf_inst.Q0 ),
    .B_N(net79),
    .Y(_252_));
 sg13g2_nor2b_1 _447_ (.A(\puf_instance.puf_loop[97].puf_inst.Q1 ),
    .B_N(net79),
    .Y(_249_));
 sg13g2_nor2b_1 _448_ (.A(\puf_instance.puf_loop[97].puf_inst.Q0 ),
    .B_N(net79),
    .Y(_250_));
 sg13g2_nor2b_1 _449_ (.A(\puf_instance.puf_loop[96].puf_inst.Q1 ),
    .B_N(net79),
    .Y(_247_));
 sg13g2_nor2b_1 _450_ (.A(\puf_instance.puf_loop[96].puf_inst.Q0 ),
    .B_N(net79),
    .Y(_248_));
 sg13g2_buf_1 _451_ (.A(net84),
    .X(_331_));
 sg13g2_nor2b_1 _452_ (.A(\puf_instance.puf_loop[95].puf_inst.Q1 ),
    .B_N(_331_),
    .Y(_245_));
 sg13g2_nor2b_1 _453_ (.A(\puf_instance.puf_loop[95].puf_inst.Q0 ),
    .B_N(_331_),
    .Y(_246_));
 sg13g2_nor2b_1 _454_ (.A(\puf_instance.puf_loop[94].puf_inst.Q1 ),
    .B_N(net78),
    .Y(_243_));
 sg13g2_nor2b_1 _455_ (.A(\puf_instance.puf_loop[94].puf_inst.Q0 ),
    .B_N(net78),
    .Y(_244_));
 sg13g2_nor2b_1 _456_ (.A(\puf_instance.puf_loop[93].puf_inst.Q1 ),
    .B_N(net78),
    .Y(_241_));
 sg13g2_nor2b_1 _457_ (.A(\puf_instance.puf_loop[93].puf_inst.Q0 ),
    .B_N(net78),
    .Y(_242_));
 sg13g2_nor2b_1 _458_ (.A(\puf_instance.puf_loop[92].puf_inst.Q1 ),
    .B_N(net78),
    .Y(_239_));
 sg13g2_nor2b_1 _459_ (.A(\puf_instance.puf_loop[92].puf_inst.Q0 ),
    .B_N(net78),
    .Y(_240_));
 sg13g2_nor2b_1 _460_ (.A(\puf_instance.puf_loop[91].puf_inst.Q1 ),
    .B_N(net78),
    .Y(_237_));
 sg13g2_nor2b_1 _461_ (.A(\puf_instance.puf_loop[91].puf_inst.Q0 ),
    .B_N(net78),
    .Y(_238_));
 sg13g2_buf_1 _462_ (.A(net84),
    .X(_332_));
 sg13g2_nor2b_1 _463_ (.A(\puf_instance.puf_loop[90].puf_inst.Q1 ),
    .B_N(net77),
    .Y(_235_));
 sg13g2_nor2b_1 _464_ (.A(\puf_instance.puf_loop[90].puf_inst.Q0 ),
    .B_N(net77),
    .Y(_236_));
 sg13g2_nor2b_1 _465_ (.A(\puf_instance.puf_loop[8].puf_inst.Q1 ),
    .B_N(_332_),
    .Y(_233_));
 sg13g2_nor2b_1 _466_ (.A(\puf_instance.puf_loop[8].puf_inst.Q0 ),
    .B_N(net77),
    .Y(_234_));
 sg13g2_nor2b_1 _467_ (.A(\puf_instance.puf_loop[89].puf_inst.Q1 ),
    .B_N(net77),
    .Y(_231_));
 sg13g2_nor2b_1 _468_ (.A(\puf_instance.puf_loop[89].puf_inst.Q0 ),
    .B_N(net77),
    .Y(_232_));
 sg13g2_nor2b_1 _469_ (.A(\puf_instance.puf_loop[88].puf_inst.Q1 ),
    .B_N(net77),
    .Y(_229_));
 sg13g2_nor2b_1 _470_ (.A(\puf_instance.puf_loop[88].puf_inst.Q0 ),
    .B_N(net77),
    .Y(_230_));
 sg13g2_nor2b_1 _471_ (.A(\puf_instance.puf_loop[87].puf_inst.Q1 ),
    .B_N(_332_),
    .Y(_227_));
 sg13g2_nor2b_1 _472_ (.A(\puf_instance.puf_loop[87].puf_inst.Q0 ),
    .B_N(net77),
    .Y(_228_));
 sg13g2_buf_1 _473_ (.A(_328_),
    .X(_333_));
 sg13g2_buf_1 _474_ (.A(net83),
    .X(_334_));
 sg13g2_nor2b_1 _475_ (.A(\puf_instance.puf_loop[86].puf_inst.Q1 ),
    .B_N(_334_),
    .Y(_225_));
 sg13g2_nor2b_1 _476_ (.A(\puf_instance.puf_loop[86].puf_inst.Q0 ),
    .B_N(_334_),
    .Y(_226_));
 sg13g2_nor2b_1 _477_ (.A(\puf_instance.puf_loop[85].puf_inst.Q1 ),
    .B_N(net76),
    .Y(_223_));
 sg13g2_nor2b_1 _478_ (.A(\puf_instance.puf_loop[85].puf_inst.Q0 ),
    .B_N(net76),
    .Y(_224_));
 sg13g2_nor2b_1 _479_ (.A(\puf_instance.puf_loop[84].puf_inst.Q1 ),
    .B_N(net76),
    .Y(_221_));
 sg13g2_nor2b_1 _480_ (.A(\puf_instance.puf_loop[84].puf_inst.Q0 ),
    .B_N(net76),
    .Y(_222_));
 sg13g2_nor2b_1 _481_ (.A(\puf_instance.puf_loop[83].puf_inst.Q1 ),
    .B_N(net76),
    .Y(_219_));
 sg13g2_nor2b_1 _482_ (.A(\puf_instance.puf_loop[83].puf_inst.Q0 ),
    .B_N(net76),
    .Y(_220_));
 sg13g2_nor2b_1 _483_ (.A(\puf_instance.puf_loop[82].puf_inst.Q1 ),
    .B_N(net76),
    .Y(_217_));
 sg13g2_nor2b_1 _484_ (.A(\puf_instance.puf_loop[82].puf_inst.Q0 ),
    .B_N(net76),
    .Y(_218_));
 sg13g2_buf_1 _485_ (.A(net83),
    .X(_335_));
 sg13g2_nor2b_1 _486_ (.A(\puf_instance.puf_loop[81].puf_inst.Q1 ),
    .B_N(net75),
    .Y(_215_));
 sg13g2_nor2b_1 _487_ (.A(\puf_instance.puf_loop[81].puf_inst.Q0 ),
    .B_N(net75),
    .Y(_216_));
 sg13g2_nor2b_1 _488_ (.A(\puf_instance.puf_loop[80].puf_inst.Q1 ),
    .B_N(net75),
    .Y(_213_));
 sg13g2_nor2b_1 _489_ (.A(\puf_instance.puf_loop[80].puf_inst.Q0 ),
    .B_N(net75),
    .Y(_214_));
 sg13g2_nor2b_1 _490_ (.A(\puf_instance.puf_loop[7].puf_inst.Q1 ),
    .B_N(_335_),
    .Y(_211_));
 sg13g2_nor2b_1 _491_ (.A(\puf_instance.puf_loop[7].puf_inst.Q0 ),
    .B_N(net75),
    .Y(_212_));
 sg13g2_nor2b_1 _492_ (.A(\puf_instance.puf_loop[79].puf_inst.Q1 ),
    .B_N(_335_),
    .Y(_209_));
 sg13g2_nor2b_1 _493_ (.A(\puf_instance.puf_loop[79].puf_inst.Q0 ),
    .B_N(net75),
    .Y(_210_));
 sg13g2_nor2b_1 _494_ (.A(\puf_instance.puf_loop[78].puf_inst.Q1 ),
    .B_N(net75),
    .Y(_207_));
 sg13g2_nor2b_1 _495_ (.A(\puf_instance.puf_loop[78].puf_inst.Q0 ),
    .B_N(net75),
    .Y(_208_));
 sg13g2_buf_1 _496_ (.A(net83),
    .X(_336_));
 sg13g2_nor2b_1 _497_ (.A(\puf_instance.puf_loop[77].puf_inst.Q1 ),
    .B_N(net74),
    .Y(_205_));
 sg13g2_nor2b_1 _498_ (.A(\puf_instance.puf_loop[77].puf_inst.Q0 ),
    .B_N(net74),
    .Y(_206_));
 sg13g2_nor2b_1 _499_ (.A(\puf_instance.puf_loop[76].puf_inst.Q1 ),
    .B_N(net74),
    .Y(_203_));
 sg13g2_nor2b_1 _500_ (.A(\puf_instance.puf_loop[76].puf_inst.Q0 ),
    .B_N(net74),
    .Y(_204_));
 sg13g2_nor2b_1 _501_ (.A(\puf_instance.puf_loop[75].puf_inst.Q1 ),
    .B_N(net74),
    .Y(_201_));
 sg13g2_nor2b_1 _502_ (.A(\puf_instance.puf_loop[75].puf_inst.Q0 ),
    .B_N(net74),
    .Y(_202_));
 sg13g2_nor2b_1 _503_ (.A(\puf_instance.puf_loop[74].puf_inst.Q1 ),
    .B_N(net74),
    .Y(_199_));
 sg13g2_nor2b_1 _504_ (.A(\puf_instance.puf_loop[74].puf_inst.Q0 ),
    .B_N(net74),
    .Y(_200_));
 sg13g2_nor2b_1 _505_ (.A(\puf_instance.puf_loop[73].puf_inst.Q1 ),
    .B_N(_336_),
    .Y(_197_));
 sg13g2_nor2b_1 _506_ (.A(\puf_instance.puf_loop[73].puf_inst.Q0 ),
    .B_N(_336_),
    .Y(_198_));
 sg13g2_buf_1 _507_ (.A(_333_),
    .X(_337_));
 sg13g2_nor2b_1 _508_ (.A(\puf_instance.puf_loop[72].puf_inst.Q1 ),
    .B_N(net73),
    .Y(_195_));
 sg13g2_nor2b_1 _509_ (.A(\puf_instance.puf_loop[72].puf_inst.Q0 ),
    .B_N(net73),
    .Y(_196_));
 sg13g2_nor2b_1 _510_ (.A(\puf_instance.puf_loop[71].puf_inst.Q1 ),
    .B_N(_337_),
    .Y(_193_));
 sg13g2_nor2b_1 _511_ (.A(\puf_instance.puf_loop[71].puf_inst.Q0 ),
    .B_N(_337_),
    .Y(_194_));
 sg13g2_nor2b_1 _512_ (.A(\puf_instance.puf_loop[70].puf_inst.Q1 ),
    .B_N(net73),
    .Y(_191_));
 sg13g2_nor2b_1 _513_ (.A(\puf_instance.puf_loop[70].puf_inst.Q0 ),
    .B_N(net73),
    .Y(_192_));
 sg13g2_nor2b_1 _514_ (.A(\puf_instance.puf_loop[6].puf_inst.Q1 ),
    .B_N(net73),
    .Y(_189_));
 sg13g2_nor2b_1 _515_ (.A(\puf_instance.puf_loop[6].puf_inst.Q0 ),
    .B_N(net73),
    .Y(_190_));
 sg13g2_nor2b_1 _516_ (.A(\puf_instance.puf_loop[69].puf_inst.Q1 ),
    .B_N(net73),
    .Y(_187_));
 sg13g2_nor2b_1 _517_ (.A(\puf_instance.puf_loop[69].puf_inst.Q0 ),
    .B_N(net73),
    .Y(_188_));
 sg13g2_buf_1 _518_ (.A(_333_),
    .X(_338_));
 sg13g2_nor2b_1 _519_ (.A(\puf_instance.puf_loop[68].puf_inst.Q1 ),
    .B_N(net72),
    .Y(_185_));
 sg13g2_nor2b_1 _520_ (.A(\puf_instance.puf_loop[68].puf_inst.Q0 ),
    .B_N(net72),
    .Y(_186_));
 sg13g2_nor2b_1 _521_ (.A(\puf_instance.puf_loop[67].puf_inst.Q1 ),
    .B_N(net72),
    .Y(_183_));
 sg13g2_nor2b_1 _522_ (.A(\puf_instance.puf_loop[67].puf_inst.Q0 ),
    .B_N(net72),
    .Y(_184_));
 sg13g2_nor2b_1 _523_ (.A(\puf_instance.puf_loop[66].puf_inst.Q1 ),
    .B_N(net72),
    .Y(_181_));
 sg13g2_nor2b_1 _524_ (.A(\puf_instance.puf_loop[66].puf_inst.Q0 ),
    .B_N(net72),
    .Y(_182_));
 sg13g2_nor2b_1 _525_ (.A(\puf_instance.puf_loop[65].puf_inst.Q1 ),
    .B_N(net72),
    .Y(_179_));
 sg13g2_nor2b_1 _526_ (.A(\puf_instance.puf_loop[65].puf_inst.Q0 ),
    .B_N(net72),
    .Y(_180_));
 sg13g2_nor2b_1 _527_ (.A(\puf_instance.puf_loop[64].puf_inst.Q1 ),
    .B_N(_338_),
    .Y(_177_));
 sg13g2_nor2b_1 _528_ (.A(\puf_instance.puf_loop[64].puf_inst.Q0 ),
    .B_N(_338_),
    .Y(_178_));
 sg13g2_buf_1 _529_ (.A(net83),
    .X(_339_));
 sg13g2_nor2b_1 _530_ (.A(\puf_instance.puf_loop[63].puf_inst.Q1 ),
    .B_N(net71),
    .Y(_175_));
 sg13g2_nor2b_1 _531_ (.A(\puf_instance.puf_loop[63].puf_inst.Q0 ),
    .B_N(net71),
    .Y(_176_));
 sg13g2_nor2b_1 _532_ (.A(\puf_instance.puf_loop[62].puf_inst.Q1 ),
    .B_N(net71),
    .Y(_173_));
 sg13g2_nor2b_1 _533_ (.A(\puf_instance.puf_loop[62].puf_inst.Q0 ),
    .B_N(net71),
    .Y(_174_));
 sg13g2_nor2b_1 _534_ (.A(\puf_instance.puf_loop[61].puf_inst.Q1 ),
    .B_N(net71),
    .Y(_171_));
 sg13g2_nor2b_1 _535_ (.A(\puf_instance.puf_loop[61].puf_inst.Q0 ),
    .B_N(net71),
    .Y(_172_));
 sg13g2_nor2b_1 _536_ (.A(\puf_instance.puf_loop[60].puf_inst.Q1 ),
    .B_N(net71),
    .Y(_169_));
 sg13g2_nor2b_1 _537_ (.A(\puf_instance.puf_loop[60].puf_inst.Q0 ),
    .B_N(net71),
    .Y(_170_));
 sg13g2_nor2b_1 _538_ (.A(\puf_instance.puf_loop[5].puf_inst.Q1 ),
    .B_N(_339_),
    .Y(_167_));
 sg13g2_nor2b_1 _539_ (.A(\puf_instance.puf_loop[5].puf_inst.Q0 ),
    .B_N(_339_),
    .Y(_168_));
 sg13g2_buf_1 _540_ (.A(net83),
    .X(_340_));
 sg13g2_nor2b_1 _541_ (.A(\puf_instance.puf_loop[59].puf_inst.Q1 ),
    .B_N(net70),
    .Y(_165_));
 sg13g2_nor2b_1 _542_ (.A(\puf_instance.puf_loop[59].puf_inst.Q0 ),
    .B_N(net70),
    .Y(_166_));
 sg13g2_nor2b_1 _543_ (.A(\puf_instance.puf_loop[58].puf_inst.Q1 ),
    .B_N(_340_),
    .Y(_163_));
 sg13g2_nor2b_1 _544_ (.A(\puf_instance.puf_loop[58].puf_inst.Q0 ),
    .B_N(_340_),
    .Y(_164_));
 sg13g2_nor2b_1 _545_ (.A(\puf_instance.puf_loop[57].puf_inst.Q1 ),
    .B_N(net70),
    .Y(_161_));
 sg13g2_nor2b_1 _546_ (.A(\puf_instance.puf_loop[57].puf_inst.Q0 ),
    .B_N(net70),
    .Y(_162_));
 sg13g2_nor2b_1 _547_ (.A(\puf_instance.puf_loop[56].puf_inst.Q1 ),
    .B_N(net70),
    .Y(_159_));
 sg13g2_nor2b_1 _548_ (.A(\puf_instance.puf_loop[56].puf_inst.Q0 ),
    .B_N(net70),
    .Y(_160_));
 sg13g2_nor2b_1 _549_ (.A(\puf_instance.puf_loop[55].puf_inst.Q1 ),
    .B_N(net70),
    .Y(_157_));
 sg13g2_nor2b_1 _550_ (.A(\puf_instance.puf_loop[55].puf_inst.Q0 ),
    .B_N(net70),
    .Y(_158_));
 sg13g2_buf_1 _551_ (.A(net83),
    .X(_341_));
 sg13g2_nor2b_1 _552_ (.A(\puf_instance.puf_loop[54].puf_inst.Q1 ),
    .B_N(net69),
    .Y(_155_));
 sg13g2_nor2b_1 _553_ (.A(\puf_instance.puf_loop[54].puf_inst.Q0 ),
    .B_N(net69),
    .Y(_156_));
 sg13g2_nor2b_1 _554_ (.A(\puf_instance.puf_loop[53].puf_inst.Q1 ),
    .B_N(net69),
    .Y(_153_));
 sg13g2_nor2b_1 _555_ (.A(\puf_instance.puf_loop[53].puf_inst.Q0 ),
    .B_N(net69),
    .Y(_154_));
 sg13g2_nor2b_1 _556_ (.A(\puf_instance.puf_loop[52].puf_inst.Q1 ),
    .B_N(net69),
    .Y(_151_));
 sg13g2_nor2b_1 _557_ (.A(\puf_instance.puf_loop[52].puf_inst.Q0 ),
    .B_N(net69),
    .Y(_152_));
 sg13g2_nor2b_1 _558_ (.A(\puf_instance.puf_loop[51].puf_inst.Q1 ),
    .B_N(net69),
    .Y(_149_));
 sg13g2_nor2b_1 _559_ (.A(\puf_instance.puf_loop[51].puf_inst.Q0 ),
    .B_N(net69),
    .Y(_150_));
 sg13g2_nor2b_1 _560_ (.A(\puf_instance.puf_loop[50].puf_inst.Q1 ),
    .B_N(_341_),
    .Y(_147_));
 sg13g2_nor2b_1 _561_ (.A(\puf_instance.puf_loop[50].puf_inst.Q0 ),
    .B_N(_341_),
    .Y(_148_));
 sg13g2_buf_1 _562_ (.A(net83),
    .X(_342_));
 sg13g2_nor2b_1 _563_ (.A(\puf_instance.puf_loop[4].puf_inst.Q1 ),
    .B_N(_342_),
    .Y(_145_));
 sg13g2_nor2b_1 _564_ (.A(\puf_instance.puf_loop[4].puf_inst.Q0 ),
    .B_N(_342_),
    .Y(_146_));
 sg13g2_nor2b_1 _565_ (.A(\puf_instance.puf_loop[49].puf_inst.Q1 ),
    .B_N(net68),
    .Y(_143_));
 sg13g2_nor2b_1 _566_ (.A(\puf_instance.puf_loop[49].puf_inst.Q0 ),
    .B_N(net68),
    .Y(_144_));
 sg13g2_nor2b_1 _567_ (.A(\puf_instance.puf_loop[48].puf_inst.Q1 ),
    .B_N(net68),
    .Y(_141_));
 sg13g2_nor2b_1 _568_ (.A(\puf_instance.puf_loop[48].puf_inst.Q0 ),
    .B_N(net68),
    .Y(_142_));
 sg13g2_nor2b_1 _569_ (.A(\puf_instance.puf_loop[47].puf_inst.Q1 ),
    .B_N(net68),
    .Y(_139_));
 sg13g2_nor2b_1 _570_ (.A(\puf_instance.puf_loop[47].puf_inst.Q0 ),
    .B_N(net68),
    .Y(_140_));
 sg13g2_nor2b_1 _571_ (.A(\puf_instance.puf_loop[46].puf_inst.Q1 ),
    .B_N(net68),
    .Y(_137_));
 sg13g2_nor2b_1 _572_ (.A(\puf_instance.puf_loop[46].puf_inst.Q0 ),
    .B_N(net68),
    .Y(_138_));
 sg13g2_buf_1 _573_ (.A(net83),
    .X(_343_));
 sg13g2_nor2b_1 _574_ (.A(\puf_instance.puf_loop[45].puf_inst.Q1 ),
    .B_N(net67),
    .Y(_135_));
 sg13g2_nor2b_1 _575_ (.A(\puf_instance.puf_loop[45].puf_inst.Q0 ),
    .B_N(net67),
    .Y(_136_));
 sg13g2_nor2b_1 _576_ (.A(\puf_instance.puf_loop[44].puf_inst.Q1 ),
    .B_N(net67),
    .Y(_133_));
 sg13g2_nor2b_1 _577_ (.A(\puf_instance.puf_loop[44].puf_inst.Q0 ),
    .B_N(net67),
    .Y(_134_));
 sg13g2_nor2b_1 _578_ (.A(\puf_instance.puf_loop[43].puf_inst.Q1 ),
    .B_N(net67),
    .Y(_131_));
 sg13g2_nor2b_1 _579_ (.A(\puf_instance.puf_loop[43].puf_inst.Q0 ),
    .B_N(net67),
    .Y(_132_));
 sg13g2_nor2b_1 _580_ (.A(\puf_instance.puf_loop[42].puf_inst.Q1 ),
    .B_N(_343_),
    .Y(_129_));
 sg13g2_nor2b_1 _581_ (.A(\puf_instance.puf_loop[42].puf_inst.Q0 ),
    .B_N(_343_),
    .Y(_130_));
 sg13g2_nor2b_1 _582_ (.A(\puf_instance.puf_loop[41].puf_inst.Q1 ),
    .B_N(net67),
    .Y(_127_));
 sg13g2_nor2b_1 _583_ (.A(\puf_instance.puf_loop[41].puf_inst.Q0 ),
    .B_N(net67),
    .Y(_128_));
 sg13g2_buf_1 _584_ (.A(_328_),
    .X(_344_));
 sg13g2_buf_1 _585_ (.A(net82),
    .X(_345_));
 sg13g2_nor2b_1 _586_ (.A(\puf_instance.puf_loop[40].puf_inst.Q1 ),
    .B_N(net66),
    .Y(_125_));
 sg13g2_nor2b_1 _587_ (.A(\puf_instance.puf_loop[40].puf_inst.Q0 ),
    .B_N(net66),
    .Y(_126_));
 sg13g2_nor2b_1 _588_ (.A(\puf_instance.puf_loop[3].puf_inst.Q1 ),
    .B_N(_345_),
    .Y(_123_));
 sg13g2_nor2b_1 _589_ (.A(\puf_instance.puf_loop[3].puf_inst.Q0 ),
    .B_N(_345_),
    .Y(_124_));
 sg13g2_nor2b_1 _590_ (.A(\puf_instance.puf_loop[39].puf_inst.Q1 ),
    .B_N(net66),
    .Y(_121_));
 sg13g2_nor2b_1 _591_ (.A(\puf_instance.puf_loop[39].puf_inst.Q0 ),
    .B_N(net66),
    .Y(_122_));
 sg13g2_nor2b_1 _592_ (.A(\puf_instance.puf_loop[38].puf_inst.Q1 ),
    .B_N(net66),
    .Y(_119_));
 sg13g2_nor2b_1 _593_ (.A(\puf_instance.puf_loop[38].puf_inst.Q0 ),
    .B_N(net66),
    .Y(_120_));
 sg13g2_nor2b_1 _594_ (.A(\puf_instance.puf_loop[37].puf_inst.Q1 ),
    .B_N(net66),
    .Y(_117_));
 sg13g2_nor2b_1 _595_ (.A(\puf_instance.puf_loop[37].puf_inst.Q0 ),
    .B_N(net66),
    .Y(_118_));
 sg13g2_buf_1 _596_ (.A(net82),
    .X(_346_));
 sg13g2_nor2b_1 _597_ (.A(\puf_instance.puf_loop[36].puf_inst.Q1 ),
    .B_N(net65),
    .Y(_115_));
 sg13g2_nor2b_1 _598_ (.A(\puf_instance.puf_loop[36].puf_inst.Q0 ),
    .B_N(net65),
    .Y(_116_));
 sg13g2_nor2b_1 _599_ (.A(\puf_instance.puf_loop[35].puf_inst.Q1 ),
    .B_N(net65),
    .Y(_113_));
 sg13g2_nor2b_1 _600_ (.A(\puf_instance.puf_loop[35].puf_inst.Q0 ),
    .B_N(net65),
    .Y(_114_));
 sg13g2_nor2b_1 _601_ (.A(\puf_instance.puf_loop[34].puf_inst.Q1 ),
    .B_N(_346_),
    .Y(_111_));
 sg13g2_nor2b_1 _602_ (.A(\puf_instance.puf_loop[34].puf_inst.Q0 ),
    .B_N(_346_),
    .Y(_112_));
 sg13g2_nor2b_1 _603_ (.A(\puf_instance.puf_loop[33].puf_inst.Q1 ),
    .B_N(net65),
    .Y(_109_));
 sg13g2_nor2b_1 _604_ (.A(\puf_instance.puf_loop[33].puf_inst.Q0 ),
    .B_N(net65),
    .Y(_110_));
 sg13g2_nor2b_1 _605_ (.A(\puf_instance.puf_loop[32].puf_inst.Q1 ),
    .B_N(net65),
    .Y(_107_));
 sg13g2_nor2b_1 _606_ (.A(\puf_instance.puf_loop[32].puf_inst.Q0 ),
    .B_N(net65),
    .Y(_108_));
 sg13g2_buf_1 _607_ (.A(net82),
    .X(_347_));
 sg13g2_nor2b_1 _608_ (.A(\puf_instance.puf_loop[31].puf_inst.Q1 ),
    .B_N(net64),
    .Y(_105_));
 sg13g2_nor2b_1 _609_ (.A(\puf_instance.puf_loop[31].puf_inst.Q0 ),
    .B_N(net64),
    .Y(_106_));
 sg13g2_nor2b_1 _610_ (.A(\puf_instance.puf_loop[30].puf_inst.Q1 ),
    .B_N(net64),
    .Y(_103_));
 sg13g2_nor2b_1 _611_ (.A(\puf_instance.puf_loop[30].puf_inst.Q0 ),
    .B_N(net64),
    .Y(_104_));
 sg13g2_nor2b_1 _612_ (.A(\puf_instance.puf_loop[2].puf_inst.Q1 ),
    .B_N(_347_),
    .Y(_101_));
 sg13g2_nor2b_1 _613_ (.A(\puf_instance.puf_loop[2].puf_inst.Q0 ),
    .B_N(_347_),
    .Y(_102_));
 sg13g2_nor2b_1 _614_ (.A(\puf_instance.puf_loop[29].puf_inst.Q1 ),
    .B_N(net64),
    .Y(_099_));
 sg13g2_nor2b_1 _615_ (.A(\puf_instance.puf_loop[29].puf_inst.Q0 ),
    .B_N(net64),
    .Y(_100_));
 sg13g2_nor2b_1 _616_ (.A(\puf_instance.puf_loop[28].puf_inst.Q1 ),
    .B_N(net64),
    .Y(_097_));
 sg13g2_nor2b_1 _617_ (.A(\puf_instance.puf_loop[28].puf_inst.Q0 ),
    .B_N(net64),
    .Y(_098_));
 sg13g2_buf_1 _618_ (.A(net82),
    .X(_348_));
 sg13g2_nor2b_1 _619_ (.A(\puf_instance.puf_loop[27].puf_inst.Q1 ),
    .B_N(net63),
    .Y(_095_));
 sg13g2_nor2b_1 _620_ (.A(\puf_instance.puf_loop[27].puf_inst.Q0 ),
    .B_N(net63),
    .Y(_096_));
 sg13g2_nor2b_1 _621_ (.A(\puf_instance.puf_loop[26].puf_inst.Q1 ),
    .B_N(net63),
    .Y(_093_));
 sg13g2_nor2b_1 _622_ (.A(\puf_instance.puf_loop[26].puf_inst.Q0 ),
    .B_N(net63),
    .Y(_094_));
 sg13g2_nor2b_1 _623_ (.A(\puf_instance.puf_loop[25].puf_inst.Q1 ),
    .B_N(net63),
    .Y(_091_));
 sg13g2_nor2b_1 _624_ (.A(\puf_instance.puf_loop[25].puf_inst.Q0 ),
    .B_N(net63),
    .Y(_092_));
 sg13g2_nor2b_1 _625_ (.A(\puf_instance.puf_loop[24].puf_inst.Q1 ),
    .B_N(net63),
    .Y(_089_));
 sg13g2_nor2b_1 _626_ (.A(\puf_instance.puf_loop[24].puf_inst.Q0 ),
    .B_N(net63),
    .Y(_090_));
 sg13g2_nor2b_1 _627_ (.A(\puf_instance.puf_loop[23].puf_inst.Q1 ),
    .B_N(_348_),
    .Y(_087_));
 sg13g2_nor2b_1 _628_ (.A(\puf_instance.puf_loop[23].puf_inst.Q0 ),
    .B_N(_348_),
    .Y(_088_));
 sg13g2_buf_1 _629_ (.A(net82),
    .X(_349_));
 sg13g2_nor2b_1 _630_ (.A(\puf_instance.puf_loop[22].puf_inst.Q1 ),
    .B_N(net62),
    .Y(_085_));
 sg13g2_nor2b_1 _631_ (.A(\puf_instance.puf_loop[22].puf_inst.Q0 ),
    .B_N(net62),
    .Y(_086_));
 sg13g2_nor2b_1 _632_ (.A(\puf_instance.puf_loop[21].puf_inst.Q1 ),
    .B_N(net62),
    .Y(_083_));
 sg13g2_nor2b_1 _633_ (.A(\puf_instance.puf_loop[21].puf_inst.Q0 ),
    .B_N(net62),
    .Y(_084_));
 sg13g2_nor2b_1 _634_ (.A(\puf_instance.puf_loop[20].puf_inst.Q1 ),
    .B_N(net62),
    .Y(_081_));
 sg13g2_nor2b_1 _635_ (.A(\puf_instance.puf_loop[20].puf_inst.Q0 ),
    .B_N(net62),
    .Y(_082_));
 sg13g2_nor2b_1 _636_ (.A(\puf_instance.puf_loop[1].puf_inst.Q1 ),
    .B_N(_349_),
    .Y(_079_));
 sg13g2_nor2b_1 _637_ (.A(\puf_instance.puf_loop[1].puf_inst.Q0 ),
    .B_N(_349_),
    .Y(_080_));
 sg13g2_nor2b_1 _638_ (.A(\puf_instance.puf_loop[19].puf_inst.Q1 ),
    .B_N(net62),
    .Y(_077_));
 sg13g2_nor2b_1 _639_ (.A(\puf_instance.puf_loop[19].puf_inst.Q0 ),
    .B_N(net62),
    .Y(_078_));
 sg13g2_buf_1 _640_ (.A(net82),
    .X(_350_));
 sg13g2_nor2b_1 _641_ (.A(\puf_instance.puf_loop[18].puf_inst.Q1 ),
    .B_N(_350_),
    .Y(_075_));
 sg13g2_nor2b_1 _642_ (.A(\puf_instance.puf_loop[18].puf_inst.Q0 ),
    .B_N(_350_),
    .Y(_076_));
 sg13g2_nor2b_1 _643_ (.A(\puf_instance.puf_loop[17].puf_inst.Q1 ),
    .B_N(net61),
    .Y(_073_));
 sg13g2_nor2b_1 _644_ (.A(\puf_instance.puf_loop[17].puf_inst.Q0 ),
    .B_N(net61),
    .Y(_074_));
 sg13g2_nor2b_1 _645_ (.A(\puf_instance.puf_loop[16].puf_inst.Q1 ),
    .B_N(net61),
    .Y(_071_));
 sg13g2_nor2b_1 _646_ (.A(\puf_instance.puf_loop[16].puf_inst.Q0 ),
    .B_N(net61),
    .Y(_072_));
 sg13g2_nor2b_1 _647_ (.A(\puf_instance.puf_loop[15].puf_inst.Q1 ),
    .B_N(net61),
    .Y(_069_));
 sg13g2_nor2b_1 _648_ (.A(\puf_instance.puf_loop[15].puf_inst.Q0 ),
    .B_N(net61),
    .Y(_070_));
 sg13g2_nor2b_1 _649_ (.A(\puf_instance.puf_loop[14].puf_inst.Q1 ),
    .B_N(net61),
    .Y(_067_));
 sg13g2_nor2b_1 _650_ (.A(\puf_instance.puf_loop[14].puf_inst.Q0 ),
    .B_N(net61),
    .Y(_068_));
 sg13g2_buf_1 _651_ (.A(net82),
    .X(_351_));
 sg13g2_nor2b_1 _652_ (.A(\puf_instance.puf_loop[13].puf_inst.Q1 ),
    .B_N(net60),
    .Y(_065_));
 sg13g2_nor2b_1 _653_ (.A(\puf_instance.puf_loop[13].puf_inst.Q0 ),
    .B_N(net60),
    .Y(_066_));
 sg13g2_nor2b_1 _654_ (.A(\puf_instance.puf_loop[12].puf_inst.Q1 ),
    .B_N(net60),
    .Y(_063_));
 sg13g2_nor2b_1 _655_ (.A(\puf_instance.puf_loop[12].puf_inst.Q0 ),
    .B_N(net60),
    .Y(_064_));
 sg13g2_nor2b_1 _656_ (.A(\puf_instance.puf_loop[127].puf_inst.Q1 ),
    .B_N(net60),
    .Y(_061_));
 sg13g2_nor2b_1 _657_ (.A(\puf_instance.puf_loop[127].puf_inst.Q0 ),
    .B_N(net60),
    .Y(_062_));
 sg13g2_nor2b_1 _658_ (.A(\puf_instance.puf_loop[126].puf_inst.Q1 ),
    .B_N(net60),
    .Y(_059_));
 sg13g2_nor2b_1 _659_ (.A(\puf_instance.puf_loop[126].puf_inst.Q0 ),
    .B_N(net60),
    .Y(_060_));
 sg13g2_nor2b_1 _660_ (.A(\puf_instance.puf_loop[125].puf_inst.Q1 ),
    .B_N(_351_),
    .Y(_057_));
 sg13g2_nor2b_1 _661_ (.A(\puf_instance.puf_loop[125].puf_inst.Q0 ),
    .B_N(_351_),
    .Y(_058_));
 sg13g2_buf_1 _662_ (.A(_344_),
    .X(_352_));
 sg13g2_nor2b_1 _663_ (.A(\puf_instance.puf_loop[124].puf_inst.Q1 ),
    .B_N(net59),
    .Y(_055_));
 sg13g2_nor2b_1 _664_ (.A(\puf_instance.puf_loop[124].puf_inst.Q0 ),
    .B_N(net59),
    .Y(_056_));
 sg13g2_nor2b_1 _665_ (.A(\puf_instance.puf_loop[123].puf_inst.Q1 ),
    .B_N(net59),
    .Y(_053_));
 sg13g2_nor2b_1 _666_ (.A(\puf_instance.puf_loop[123].puf_inst.Q0 ),
    .B_N(net59),
    .Y(_054_));
 sg13g2_nor2b_1 _667_ (.A(\puf_instance.puf_loop[122].puf_inst.Q1 ),
    .B_N(net59),
    .Y(_051_));
 sg13g2_nor2b_1 _668_ (.A(\puf_instance.puf_loop[122].puf_inst.Q0 ),
    .B_N(net59),
    .Y(_052_));
 sg13g2_nor2b_1 _669_ (.A(\puf_instance.puf_loop[121].puf_inst.Q1 ),
    .B_N(net59),
    .Y(_049_));
 sg13g2_nor2b_1 _670_ (.A(\puf_instance.puf_loop[121].puf_inst.Q0 ),
    .B_N(net59),
    .Y(_050_));
 sg13g2_nor2b_1 _671_ (.A(\puf_instance.puf_loop[120].puf_inst.Q1 ),
    .B_N(_352_),
    .Y(_047_));
 sg13g2_nor2b_1 _672_ (.A(\puf_instance.puf_loop[120].puf_inst.Q0 ),
    .B_N(_352_),
    .Y(_048_));
 sg13g2_buf_1 _673_ (.A(net82),
    .X(_353_));
 sg13g2_nor2b_1 _674_ (.A(\puf_instance.puf_loop[11].puf_inst.Q1 ),
    .B_N(_353_),
    .Y(_045_));
 sg13g2_nor2b_1 _675_ (.A(\puf_instance.puf_loop[11].puf_inst.Q0 ),
    .B_N(_353_),
    .Y(_046_));
 sg13g2_nor2b_1 _676_ (.A(\puf_instance.puf_loop[119].puf_inst.Q1 ),
    .B_N(net58),
    .Y(_043_));
 sg13g2_nor2b_1 _677_ (.A(\puf_instance.puf_loop[119].puf_inst.Q0 ),
    .B_N(net58),
    .Y(_044_));
 sg13g2_nor2b_1 _678_ (.A(\puf_instance.puf_loop[118].puf_inst.Q1 ),
    .B_N(net58),
    .Y(_041_));
 sg13g2_nor2b_1 _679_ (.A(\puf_instance.puf_loop[118].puf_inst.Q0 ),
    .B_N(net58),
    .Y(_042_));
 sg13g2_nor2b_1 _680_ (.A(\puf_instance.puf_loop[117].puf_inst.Q1 ),
    .B_N(net58),
    .Y(_039_));
 sg13g2_nor2b_1 _681_ (.A(\puf_instance.puf_loop[117].puf_inst.Q0 ),
    .B_N(net58),
    .Y(_040_));
 sg13g2_nor2b_1 _682_ (.A(\puf_instance.puf_loop[116].puf_inst.Q1 ),
    .B_N(net58),
    .Y(_037_));
 sg13g2_nor2b_1 _683_ (.A(\puf_instance.puf_loop[116].puf_inst.Q0 ),
    .B_N(net58),
    .Y(_038_));
 sg13g2_buf_1 _684_ (.A(_344_),
    .X(_354_));
 sg13g2_nor2b_1 _685_ (.A(\puf_instance.puf_loop[115].puf_inst.Q1 ),
    .B_N(net57),
    .Y(_035_));
 sg13g2_nor2b_1 _686_ (.A(\puf_instance.puf_loop[115].puf_inst.Q0 ),
    .B_N(net57),
    .Y(_036_));
 sg13g2_nor2b_1 _687_ (.A(\puf_instance.puf_loop[114].puf_inst.Q1 ),
    .B_N(net57),
    .Y(_033_));
 sg13g2_nor2b_1 _688_ (.A(\puf_instance.puf_loop[114].puf_inst.Q0 ),
    .B_N(net57),
    .Y(_034_));
 sg13g2_nor2b_1 _689_ (.A(\puf_instance.puf_loop[113].puf_inst.Q1 ),
    .B_N(net57),
    .Y(_031_));
 sg13g2_nor2b_1 _690_ (.A(\puf_instance.puf_loop[113].puf_inst.Q0 ),
    .B_N(net57),
    .Y(_032_));
 sg13g2_nor2b_1 _691_ (.A(\puf_instance.puf_loop[112].puf_inst.Q1 ),
    .B_N(net57),
    .Y(_029_));
 sg13g2_nor2b_1 _692_ (.A(\puf_instance.puf_loop[112].puf_inst.Q0 ),
    .B_N(net57),
    .Y(_030_));
 sg13g2_nor2b_1 _693_ (.A(\puf_instance.puf_loop[111].puf_inst.Q1 ),
    .B_N(_354_),
    .Y(_027_));
 sg13g2_nor2b_1 _694_ (.A(\puf_instance.puf_loop[111].puf_inst.Q0 ),
    .B_N(_354_),
    .Y(_028_));
 sg13g2_buf_1 _695_ (.A(_328_),
    .X(_355_));
 sg13g2_nor2b_1 _696_ (.A(\puf_instance.puf_loop[110].puf_inst.Q1 ),
    .B_N(net81),
    .Y(_025_));
 sg13g2_nor2b_1 _697_ (.A(\puf_instance.puf_loop[110].puf_inst.Q0 ),
    .B_N(net81),
    .Y(_026_));
 sg13g2_nor2b_1 _698_ (.A(\puf_instance.puf_loop[10].puf_inst.Q1 ),
    .B_N(net81),
    .Y(_023_));
 sg13g2_nor2b_1 _699_ (.A(\puf_instance.puf_loop[10].puf_inst.Q0 ),
    .B_N(net81),
    .Y(_024_));
 sg13g2_nor2b_1 _700_ (.A(\puf_instance.puf_loop[109].puf_inst.Q1 ),
    .B_N(net81),
    .Y(_021_));
 sg13g2_nor2b_1 _701_ (.A(\puf_instance.puf_loop[109].puf_inst.Q0 ),
    .B_N(net81),
    .Y(_022_));
 sg13g2_nor2b_1 _702_ (.A(\puf_instance.puf_loop[108].puf_inst.Q1 ),
    .B_N(net81),
    .Y(_019_));
 sg13g2_nor2b_1 _703_ (.A(\puf_instance.puf_loop[108].puf_inst.Q0 ),
    .B_N(net81),
    .Y(_020_));
 sg13g2_nor2b_1 _704_ (.A(\puf_instance.puf_loop[107].puf_inst.Q1 ),
    .B_N(_355_),
    .Y(_017_));
 sg13g2_nor2b_1 _705_ (.A(\puf_instance.puf_loop[107].puf_inst.Q0 ),
    .B_N(_355_),
    .Y(_018_));
 sg13g2_buf_1 _706_ (.A(_328_),
    .X(_356_));
 sg13g2_nor2b_1 _707_ (.A(\puf_instance.puf_loop[106].puf_inst.Q1 ),
    .B_N(net80),
    .Y(_015_));
 sg13g2_nor2b_1 _708_ (.A(\puf_instance.puf_loop[106].puf_inst.Q0 ),
    .B_N(net80),
    .Y(_016_));
 sg13g2_nor2b_1 _709_ (.A(\puf_instance.puf_loop[105].puf_inst.Q1 ),
    .B_N(net80),
    .Y(_013_));
 sg13g2_nor2b_1 _710_ (.A(\puf_instance.puf_loop[105].puf_inst.Q0 ),
    .B_N(net80),
    .Y(_014_));
 sg13g2_nor2b_1 _711_ (.A(\puf_instance.puf_loop[104].puf_inst.Q1 ),
    .B_N(_356_),
    .Y(_011_));
 sg13g2_nor2b_1 _712_ (.A(\puf_instance.puf_loop[104].puf_inst.Q0 ),
    .B_N(_356_),
    .Y(_012_));
 sg13g2_nor2b_1 _713_ (.A(\puf_instance.puf_loop[103].puf_inst.Q1 ),
    .B_N(net80),
    .Y(_009_));
 sg13g2_nor2b_1 _714_ (.A(\puf_instance.puf_loop[103].puf_inst.Q0 ),
    .B_N(net80),
    .Y(_010_));
 sg13g2_nor2b_1 _715_ (.A(\puf_instance.puf_loop[102].puf_inst.Q1 ),
    .B_N(net80),
    .Y(_007_));
 sg13g2_nor2b_1 _716_ (.A(\puf_instance.puf_loop[102].puf_inst.Q0 ),
    .B_N(net80),
    .Y(_008_));
 sg13g2_nor2b_1 _717_ (.A(\puf_instance.puf_loop[101].puf_inst.Q1 ),
    .B_N(net84),
    .Y(_005_));
 sg13g2_nor2b_1 _718_ (.A(\puf_instance.puf_loop[101].puf_inst.Q0 ),
    .B_N(net84),
    .Y(_006_));
 sg13g2_nor2b_1 _719_ (.A(\puf_instance.puf_loop[100].puf_inst.Q1 ),
    .B_N(net84),
    .Y(_003_));
 sg13g2_nor2b_1 _720_ (.A(\puf_instance.puf_loop[100].puf_inst.Q0 ),
    .B_N(net84),
    .Y(_004_));
 sg13g2_nor2b_1 _721_ (.A(net4),
    .B_N(_329_),
    .Y(_001_));
 sg13g2_nor2b_1 _722_ (.A(\puf_instance.puf_loop[0].puf_inst.Q1 ),
    .B_N(net84),
    .Y(_000_));
 sg13g2_nor2b_1 _723_ (.A(\puf_instance.puf_loop[0].puf_inst.Q0 ),
    .B_N(_329_),
    .Y(_002_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \puf_instance.puf_loop[0].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_108  (.L_HI(net108));
 sg13g2_buf_1 _726_ (.A(net92),
    .X(uio_oe[0]));
 sg13g2_buf_1 _727_ (.A(net93),
    .X(uio_oe[1]));
 sg13g2_buf_1 _728_ (.A(net94),
    .X(uio_oe[2]));
 sg13g2_buf_1 _729_ (.A(net95),
    .X(uio_oe[3]));
 sg13g2_buf_1 _730_ (.A(net96),
    .X(uio_oe[4]));
 sg13g2_buf_1 _731_ (.A(net97),
    .X(uio_oe[5]));
 sg13g2_buf_1 _732_ (.A(net98),
    .X(uio_oe[6]));
 sg13g2_buf_1 _733_ (.A(net99),
    .X(uio_oe[7]));
 sg13g2_buf_1 _734_ (.A(net100),
    .X(uio_out[0]));
 sg13g2_buf_1 _735_ (.A(net101),
    .X(uio_out[1]));
 sg13g2_buf_1 _736_ (.A(net102),
    .X(uio_out[2]));
 sg13g2_buf_1 _737_ (.A(net103),
    .X(uio_out[3]));
 sg13g2_buf_1 _738_ (.A(net104),
    .X(uio_out[4]));
 sg13g2_buf_1 _739_ (.A(net105),
    .X(uio_out[5]));
 sg13g2_buf_1 _740_ (.A(net106),
    .X(uio_out[6]));
 sg13g2_buf_1 _741_ (.A(net107),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[0]$_DFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net91),
    .D(_257_),
    .Q_N(_358_),
    .Q(net5));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[1]$_DFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net91),
    .D(_258_),
    .Q_N(_359_),
    .Q(net6));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[2]$_DFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net91),
    .D(_259_),
    .Q_N(_360_),
    .Q(net7));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[3]$_DFF_PN0_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net91),
    .D(_260_),
    .Q_N(_361_),
    .Q(net8));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[4]$_DFF_PN0_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net91),
    .D(_261_),
    .Q_N(_362_),
    .Q(net9));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[5]$_DFF_PN0_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net1),
    .D(_262_),
    .Q_N(_363_),
    .Q(net10));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[6]$_DFF_PN0_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net91),
    .D(_263_),
    .Q_N(_364_),
    .Q(net11));
 sg13g2_dfrbp_1 \puf_instance.OUT_reg[7]$_DFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net91),
    .D(_264_),
    .Q_N(_357_),
    .Q(net12));
 sg13g2_dllrq_1 \puf_instance.puf_loop[0].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_000_),
    .GATE_N(net48),
    .RESET_B(net108),
    .Q(\puf_instance.puf_loop[0].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[0].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_002_),
    .GATE_N(net48),
    .RESET_B(net109),
    .Q(\puf_instance.puf_loop[0].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[100].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_003_),
    .GATE_N(net18),
    .RESET_B(net110),
    .Q(\puf_instance.puf_loop[100].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[100].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_004_),
    .GATE_N(net20),
    .RESET_B(net111),
    .Q(\puf_instance.puf_loop[100].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[101].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_005_),
    .GATE_N(net32),
    .RESET_B(net112),
    .Q(\puf_instance.puf_loop[101].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[101].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_006_),
    .GATE_N(net32),
    .RESET_B(net113),
    .Q(\puf_instance.puf_loop[101].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[102].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_007_),
    .GATE_N(net37),
    .RESET_B(net114),
    .Q(\puf_instance.puf_loop[102].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[102].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_008_),
    .GATE_N(net18),
    .RESET_B(net115),
    .Q(\puf_instance.puf_loop[102].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[103].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_009_),
    .GATE_N(net37),
    .RESET_B(net116),
    .Q(\puf_instance.puf_loop[103].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[103].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_010_),
    .GATE_N(net37),
    .RESET_B(net117),
    .Q(\puf_instance.puf_loop[103].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[104].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_011_),
    .GATE_N(net42),
    .RESET_B(net118),
    .Q(\puf_instance.puf_loop[104].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[104].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_012_),
    .GATE_N(net42),
    .RESET_B(net119),
    .Q(\puf_instance.puf_loop[104].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[105].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_013_),
    .GATE_N(net44),
    .RESET_B(net120),
    .Q(\puf_instance.puf_loop[105].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[105].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_014_),
    .GATE_N(net44),
    .RESET_B(net121),
    .Q(\puf_instance.puf_loop[105].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[106].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_015_),
    .GATE_N(net42),
    .RESET_B(net122),
    .Q(\puf_instance.puf_loop[106].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[106].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_016_),
    .GATE_N(net42),
    .RESET_B(net123),
    .Q(\puf_instance.puf_loop[106].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[107].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_017_),
    .GATE_N(net43),
    .RESET_B(net124),
    .Q(\puf_instance.puf_loop[107].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[107].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_018_),
    .GATE_N(net43),
    .RESET_B(net125),
    .Q(\puf_instance.puf_loop[107].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[108].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_019_),
    .GATE_N(net18),
    .RESET_B(net126),
    .Q(\puf_instance.puf_loop[108].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[108].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_020_),
    .GATE_N(net18),
    .RESET_B(net127),
    .Q(\puf_instance.puf_loop[108].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[109].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_021_),
    .GATE_N(net32),
    .RESET_B(net128),
    .Q(\puf_instance.puf_loop[109].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[109].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_022_),
    .GATE_N(net32),
    .RESET_B(net129),
    .Q(\puf_instance.puf_loop[109].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[10].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_023_),
    .GATE_N(net51),
    .RESET_B(net130),
    .Q(\puf_instance.puf_loop[10].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[10].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_024_),
    .GATE_N(net51),
    .RESET_B(net131),
    .Q(\puf_instance.puf_loop[10].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[110].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_025_),
    .GATE_N(net30),
    .RESET_B(net132),
    .Q(\puf_instance.puf_loop[110].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[110].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_026_),
    .GATE_N(net29),
    .RESET_B(net133),
    .Q(\puf_instance.puf_loop[110].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[111].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_027_),
    .GATE_N(net44),
    .RESET_B(net134),
    .Q(\puf_instance.puf_loop[111].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[111].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_028_),
    .GATE_N(net44),
    .RESET_B(net135),
    .Q(\puf_instance.puf_loop[111].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[112].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_029_),
    .GATE_N(net41),
    .RESET_B(net136),
    .Q(\puf_instance.puf_loop[112].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[112].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_030_),
    .GATE_N(net41),
    .RESET_B(net137),
    .Q(\puf_instance.puf_loop[112].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[113].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_031_),
    .GATE_N(net40),
    .RESET_B(net138),
    .Q(\puf_instance.puf_loop[113].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[113].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_032_),
    .GATE_N(net40),
    .RESET_B(net139),
    .Q(\puf_instance.puf_loop[113].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[114].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_033_),
    .GATE_N(net41),
    .RESET_B(net140),
    .Q(\puf_instance.puf_loop[114].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[114].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_034_),
    .GATE_N(net41),
    .RESET_B(net141),
    .Q(\puf_instance.puf_loop[114].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[115].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_035_),
    .GATE_N(net43),
    .RESET_B(net142),
    .Q(\puf_instance.puf_loop[115].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[115].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_036_),
    .GATE_N(net43),
    .RESET_B(net143),
    .Q(\puf_instance.puf_loop[115].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[116].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_037_),
    .GATE_N(net20),
    .RESET_B(net144),
    .Q(\puf_instance.puf_loop[116].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[116].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_038_),
    .GATE_N(net20),
    .RESET_B(net145),
    .Q(\puf_instance.puf_loop[116].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[117].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_039_),
    .GATE_N(net32),
    .RESET_B(net146),
    .Q(\puf_instance.puf_loop[117].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[117].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_040_),
    .GATE_N(net32),
    .RESET_B(net147),
    .Q(\puf_instance.puf_loop[117].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[118].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_041_),
    .GATE_N(net30),
    .RESET_B(net148),
    .Q(\puf_instance.puf_loop[118].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[118].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_042_),
    .GATE_N(net30),
    .RESET_B(net149),
    .Q(\puf_instance.puf_loop[118].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[119].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_043_),
    .GATE_N(net48),
    .RESET_B(net150),
    .Q(\puf_instance.puf_loop[119].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[119].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_044_),
    .GATE_N(net48),
    .RESET_B(net151),
    .Q(\puf_instance.puf_loop[119].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[11].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_045_),
    .GATE_N(net46),
    .RESET_B(net152),
    .Q(\puf_instance.puf_loop[11].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[11].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_046_),
    .GATE_N(net46),
    .RESET_B(net153),
    .Q(\puf_instance.puf_loop[11].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[120].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_047_),
    .GATE_N(net42),
    .RESET_B(net154),
    .Q(\puf_instance.puf_loop[120].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[120].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_048_),
    .GATE_N(net42),
    .RESET_B(net155),
    .Q(\puf_instance.puf_loop[120].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[121].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_049_),
    .GATE_N(net40),
    .RESET_B(net156),
    .Q(\puf_instance.puf_loop[121].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[121].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_050_),
    .GATE_N(net40),
    .RESET_B(net157),
    .Q(\puf_instance.puf_loop[121].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[122].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_051_),
    .GATE_N(net40),
    .RESET_B(net158),
    .Q(\puf_instance.puf_loop[122].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[122].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_052_),
    .GATE_N(net40),
    .RESET_B(net159),
    .Q(\puf_instance.puf_loop[122].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[123].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_053_),
    .GATE_N(net43),
    .RESET_B(net160),
    .Q(\puf_instance.puf_loop[123].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[123].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_054_),
    .GATE_N(net43),
    .RESET_B(net161),
    .Q(\puf_instance.puf_loop[123].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[124].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_055_),
    .GATE_N(net44),
    .RESET_B(net162),
    .Q(\puf_instance.puf_loop[124].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[124].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_056_),
    .GATE_N(net44),
    .RESET_B(net163),
    .Q(\puf_instance.puf_loop[124].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[125].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_057_),
    .GATE_N(net33),
    .RESET_B(net164),
    .Q(\puf_instance.puf_loop[125].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[125].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_058_),
    .GATE_N(net33),
    .RESET_B(net165),
    .Q(\puf_instance.puf_loop[125].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[126].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_059_),
    .GATE_N(net29),
    .RESET_B(net166),
    .Q(\puf_instance.puf_loop[126].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[126].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_060_),
    .GATE_N(net30),
    .RESET_B(net167),
    .Q(\puf_instance.puf_loop[126].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[127].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_061_),
    .GATE_N(net48),
    .RESET_B(net168),
    .Q(\puf_instance.puf_loop[127].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[127].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_062_),
    .GATE_N(net48),
    .RESET_B(net169),
    .Q(\puf_instance.puf_loop[127].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[12].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_063_),
    .GATE_N(net46),
    .RESET_B(net170),
    .Q(\puf_instance.puf_loop[12].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[12].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_064_),
    .GATE_N(net46),
    .RESET_B(net171),
    .Q(\puf_instance.puf_loop[12].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[13].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_065_),
    .GATE_N(net46),
    .RESET_B(net172),
    .Q(\puf_instance.puf_loop[13].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[13].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_066_),
    .GATE_N(net46),
    .RESET_B(net173),
    .Q(\puf_instance.puf_loop[13].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[14].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_067_),
    .GATE_N(net52),
    .RESET_B(net174),
    .Q(\puf_instance.puf_loop[14].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[14].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_068_),
    .GATE_N(net52),
    .RESET_B(net175),
    .Q(\puf_instance.puf_loop[14].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[15].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_069_),
    .GATE_N(net51),
    .RESET_B(net176),
    .Q(\puf_instance.puf_loop[15].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[15].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_070_),
    .GATE_N(net51),
    .RESET_B(net177),
    .Q(\puf_instance.puf_loop[15].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[16].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_071_),
    .GATE_N(net50),
    .RESET_B(net178),
    .Q(\puf_instance.puf_loop[16].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[16].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_072_),
    .GATE_N(net50),
    .RESET_B(net179),
    .Q(\puf_instance.puf_loop[16].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[17].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_073_),
    .GATE_N(net50),
    .RESET_B(net180),
    .Q(\puf_instance.puf_loop[17].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[17].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_074_),
    .GATE_N(net50),
    .RESET_B(net181),
    .Q(\puf_instance.puf_loop[17].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[18].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_075_),
    .GATE_N(net52),
    .RESET_B(net182),
    .Q(\puf_instance.puf_loop[18].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[18].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_076_),
    .GATE_N(net52),
    .RESET_B(net183),
    .Q(\puf_instance.puf_loop[18].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[19].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_077_),
    .GATE_N(net47),
    .RESET_B(net184),
    .Q(\puf_instance.puf_loop[19].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[19].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_078_),
    .GATE_N(net47),
    .RESET_B(net185),
    .Q(\puf_instance.puf_loop[19].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[1].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_079_),
    .GATE_N(net49),
    .RESET_B(net186),
    .Q(\puf_instance.puf_loop[1].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[1].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_080_),
    .GATE_N(net49),
    .RESET_B(net187),
    .Q(\puf_instance.puf_loop[1].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[20].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_081_),
    .GATE_N(net46),
    .RESET_B(net188),
    .Q(\puf_instance.puf_loop[20].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[20].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_082_),
    .GATE_N(net47),
    .RESET_B(net189),
    .Q(\puf_instance.puf_loop[20].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[21].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_083_),
    .GATE_N(net46),
    .RESET_B(net190),
    .Q(\puf_instance.puf_loop[21].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[21].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_084_),
    .GATE_N(net47),
    .RESET_B(net191),
    .Q(\puf_instance.puf_loop[21].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[22].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_085_),
    .GATE_N(net53),
    .RESET_B(net192),
    .Q(\puf_instance.puf_loop[22].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[22].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_086_),
    .GATE_N(net53),
    .RESET_B(net193),
    .Q(\puf_instance.puf_loop[22].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[23].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_087_),
    .GATE_N(net51),
    .RESET_B(net194),
    .Q(\puf_instance.puf_loop[23].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[23].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_088_),
    .GATE_N(net51),
    .RESET_B(net195),
    .Q(\puf_instance.puf_loop[23].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[24].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_089_),
    .GATE_N(net49),
    .RESET_B(net196),
    .Q(\puf_instance.puf_loop[24].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[24].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_090_),
    .GATE_N(net50),
    .RESET_B(net197),
    .Q(\puf_instance.puf_loop[24].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[25].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_091_),
    .GATE_N(net50),
    .RESET_B(net198),
    .Q(\puf_instance.puf_loop[25].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[25].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_092_),
    .GATE_N(net50),
    .RESET_B(net199),
    .Q(\puf_instance.puf_loop[25].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[26].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_093_),
    .GATE_N(net51),
    .RESET_B(net200),
    .Q(\puf_instance.puf_loop[26].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[26].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_094_),
    .GATE_N(net51),
    .RESET_B(net201),
    .Q(\puf_instance.puf_loop[26].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[27].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_095_),
    .GATE_N(net47),
    .RESET_B(net202),
    .Q(\puf_instance.puf_loop[27].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[27].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_096_),
    .GATE_N(net47),
    .RESET_B(net203),
    .Q(\puf_instance.puf_loop[27].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[28].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_097_),
    .GATE_N(net53),
    .RESET_B(net204),
    .Q(\puf_instance.puf_loop[28].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[28].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_098_),
    .GATE_N(net53),
    .RESET_B(net205),
    .Q(\puf_instance.puf_loop[28].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[29].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_099_),
    .GATE_N(net53),
    .RESET_B(net206),
    .Q(\puf_instance.puf_loop[29].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[29].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_100_),
    .GATE_N(net53),
    .RESET_B(net207),
    .Q(\puf_instance.puf_loop[29].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[2].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_101_),
    .GATE_N(net52),
    .RESET_B(net208),
    .Q(\puf_instance.puf_loop[2].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[2].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_102_),
    .GATE_N(net52),
    .RESET_B(net209),
    .Q(\puf_instance.puf_loop[2].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[30].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_103_),
    .GATE_N(net53),
    .RESET_B(net210),
    .Q(\puf_instance.puf_loop[30].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[30].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_104_),
    .GATE_N(net53),
    .RESET_B(net211),
    .Q(\puf_instance.puf_loop[30].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[31].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_105_),
    .GATE_N(net52),
    .RESET_B(net212),
    .Q(\puf_instance.puf_loop[31].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[31].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_106_),
    .GATE_N(net52),
    .RESET_B(net213),
    .Q(\puf_instance.puf_loop[31].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[32].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_107_),
    .GATE_N(net13),
    .RESET_B(net214),
    .Q(\puf_instance.puf_loop[32].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[32].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_108_),
    .GATE_N(net13),
    .RESET_B(net215),
    .Q(\puf_instance.puf_loop[32].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[33].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_109_),
    .GATE_N(net13),
    .RESET_B(net216),
    .Q(\puf_instance.puf_loop[33].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[33].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_110_),
    .GATE_N(net13),
    .RESET_B(net217),
    .Q(\puf_instance.puf_loop[33].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[34].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_111_),
    .GATE_N(net26),
    .RESET_B(net218),
    .Q(\puf_instance.puf_loop[34].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[34].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_112_),
    .GATE_N(net26),
    .RESET_B(net219),
    .Q(\puf_instance.puf_loop[34].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[35].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_113_),
    .GATE_N(net23),
    .RESET_B(net220),
    .Q(\puf_instance.puf_loop[35].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[35].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_114_),
    .GATE_N(net23),
    .RESET_B(net221),
    .Q(\puf_instance.puf_loop[35].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[36].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_115_),
    .GATE_N(net25),
    .RESET_B(net222),
    .Q(\puf_instance.puf_loop[36].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[36].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_116_),
    .GATE_N(net25),
    .RESET_B(net223),
    .Q(\puf_instance.puf_loop[36].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[37].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_117_),
    .GATE_N(net27),
    .RESET_B(net224),
    .Q(\puf_instance.puf_loop[37].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[37].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_118_),
    .GATE_N(net27),
    .RESET_B(net225),
    .Q(\puf_instance.puf_loop[37].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[38].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_119_),
    .GATE_N(net29),
    .RESET_B(net226),
    .Q(\puf_instance.puf_loop[38].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[38].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_120_),
    .GATE_N(net29),
    .RESET_B(net227),
    .Q(\puf_instance.puf_loop[38].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[39].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_121_),
    .GATE_N(net19),
    .RESET_B(net228),
    .Q(\puf_instance.puf_loop[39].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[39].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_122_),
    .GATE_N(net19),
    .RESET_B(net229),
    .Q(\puf_instance.puf_loop[39].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[3].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_123_),
    .GATE_N(net31),
    .RESET_B(net230),
    .Q(\puf_instance.puf_loop[3].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[3].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_124_),
    .GATE_N(net31),
    .RESET_B(net231),
    .Q(\puf_instance.puf_loop[3].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[40].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_125_),
    .GATE_N(net24),
    .RESET_B(net232),
    .Q(\puf_instance.puf_loop[40].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[40].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_126_),
    .GATE_N(net24),
    .RESET_B(net233),
    .Q(\puf_instance.puf_loop[40].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[41].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_127_),
    .GATE_N(net23),
    .RESET_B(net234),
    .Q(\puf_instance.puf_loop[41].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[41].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_128_),
    .GATE_N(net23),
    .RESET_B(net235),
    .Q(\puf_instance.puf_loop[41].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[42].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_129_),
    .GATE_N(net26),
    .RESET_B(net236),
    .Q(\puf_instance.puf_loop[42].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[42].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_130_),
    .GATE_N(net26),
    .RESET_B(net237),
    .Q(\puf_instance.puf_loop[42].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[43].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_131_),
    .GATE_N(net23),
    .RESET_B(net238),
    .Q(\puf_instance.puf_loop[43].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[43].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_132_),
    .GATE_N(net23),
    .RESET_B(net239),
    .Q(\puf_instance.puf_loop[43].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[44].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_133_),
    .GATE_N(net25),
    .RESET_B(net240),
    .Q(\puf_instance.puf_loop[44].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[44].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_134_),
    .GATE_N(net25),
    .RESET_B(net241),
    .Q(\puf_instance.puf_loop[44].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[45].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_135_),
    .GATE_N(net25),
    .RESET_B(net242),
    .Q(\puf_instance.puf_loop[45].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[45].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_136_),
    .GATE_N(net25),
    .RESET_B(net243),
    .Q(\puf_instance.puf_loop[45].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[46].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_137_),
    .GATE_N(net31),
    .RESET_B(net244),
    .Q(\puf_instance.puf_loop[46].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[46].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_138_),
    .GATE_N(net31),
    .RESET_B(net245),
    .Q(\puf_instance.puf_loop[46].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[47].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_139_),
    .GATE_N(net19),
    .RESET_B(net246),
    .Q(\puf_instance.puf_loop[47].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[47].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_140_),
    .GATE_N(net19),
    .RESET_B(net247),
    .Q(\puf_instance.puf_loop[47].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[48].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_141_),
    .GATE_N(net24),
    .RESET_B(net248),
    .Q(\puf_instance.puf_loop[48].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[48].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_142_),
    .GATE_N(net24),
    .RESET_B(net249),
    .Q(\puf_instance.puf_loop[48].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[49].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_143_),
    .GATE_N(net13),
    .RESET_B(net250),
    .Q(\puf_instance.puf_loop[49].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[49].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_144_),
    .GATE_N(net13),
    .RESET_B(net251),
    .Q(\puf_instance.puf_loop[49].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[4].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_145_),
    .GATE_N(net31),
    .RESET_B(net252),
    .Q(\puf_instance.puf_loop[4].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[4].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_146_),
    .GATE_N(net31),
    .RESET_B(net253),
    .Q(\puf_instance.puf_loop[4].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[50].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_147_),
    .GATE_N(net26),
    .RESET_B(net254),
    .Q(\puf_instance.puf_loop[50].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[50].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_148_),
    .GATE_N(net26),
    .RESET_B(net255),
    .Q(\puf_instance.puf_loop[50].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[51].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_149_),
    .GATE_N(net23),
    .RESET_B(net256),
    .Q(\puf_instance.puf_loop[51].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[51].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_150_),
    .GATE_N(net23),
    .RESET_B(net257),
    .Q(\puf_instance.puf_loop[51].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[52].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_151_),
    .GATE_N(net27),
    .RESET_B(net258),
    .Q(\puf_instance.puf_loop[52].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[52].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_152_),
    .GATE_N(net25),
    .RESET_B(net259),
    .Q(\puf_instance.puf_loop[52].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[53].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_153_),
    .GATE_N(net27),
    .RESET_B(net260),
    .Q(\puf_instance.puf_loop[53].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[53].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_154_),
    .GATE_N(net27),
    .RESET_B(net261),
    .Q(\puf_instance.puf_loop[53].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[54].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_155_),
    .GATE_N(net24),
    .RESET_B(net262),
    .Q(\puf_instance.puf_loop[54].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[54].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_156_),
    .GATE_N(net24),
    .RESET_B(net263),
    .Q(\puf_instance.puf_loop[54].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[55].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_157_),
    .GATE_N(net14),
    .RESET_B(net264),
    .Q(\puf_instance.puf_loop[55].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[55].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_158_),
    .GATE_N(net14),
    .RESET_B(net265),
    .Q(\puf_instance.puf_loop[55].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[56].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_159_),
    .GATE_N(net14),
    .RESET_B(net266),
    .Q(\puf_instance.puf_loop[56].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[56].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_160_),
    .GATE_N(net14),
    .RESET_B(net267),
    .Q(\puf_instance.puf_loop[56].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[57].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_161_),
    .GATE_N(net13),
    .RESET_B(net268),
    .Q(\puf_instance.puf_loop[57].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[57].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_162_),
    .GATE_N(net13),
    .RESET_B(net269),
    .Q(\puf_instance.puf_loop[57].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[58].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_163_),
    .GATE_N(net26),
    .RESET_B(net270),
    .Q(\puf_instance.puf_loop[58].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[58].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_164_),
    .GATE_N(net28),
    .RESET_B(net271),
    .Q(\puf_instance.puf_loop[58].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[59].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_165_),
    .GATE_N(net24),
    .RESET_B(net272),
    .Q(\puf_instance.puf_loop[59].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[59].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_166_),
    .GATE_N(net24),
    .RESET_B(net273),
    .Q(\puf_instance.puf_loop[59].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[5].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_167_),
    .GATE_N(net31),
    .RESET_B(net274),
    .Q(\puf_instance.puf_loop[5].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[5].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_168_),
    .GATE_N(net31),
    .RESET_B(net275),
    .Q(\puf_instance.puf_loop[5].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[60].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_169_),
    .GATE_N(net25),
    .RESET_B(net276),
    .Q(\puf_instance.puf_loop[60].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[60].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_170_),
    .GATE_N(net27),
    .RESET_B(net277),
    .Q(\puf_instance.puf_loop[60].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[61].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_171_),
    .GATE_N(net27),
    .RESET_B(net278),
    .Q(\puf_instance.puf_loop[61].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[61].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_172_),
    .GATE_N(net32),
    .RESET_B(net279),
    .Q(\puf_instance.puf_loop[61].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[62].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_173_),
    .GATE_N(net29),
    .RESET_B(net280),
    .Q(\puf_instance.puf_loop[62].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[62].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_174_),
    .GATE_N(net29),
    .RESET_B(net281),
    .Q(\puf_instance.puf_loop[62].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[63].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_175_),
    .GATE_N(net29),
    .RESET_B(net282),
    .Q(\puf_instance.puf_loop[63].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[63].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_176_),
    .GATE_N(net29),
    .RESET_B(net283),
    .Q(\puf_instance.puf_loop[63].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[64].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_177_),
    .GATE_N(net34),
    .RESET_B(net284),
    .Q(\puf_instance.puf_loop[64].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[64].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_178_),
    .GATE_N(net34),
    .RESET_B(net285),
    .Q(\puf_instance.puf_loop[64].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[65].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_179_),
    .GATE_N(net34),
    .RESET_B(net286),
    .Q(\puf_instance.puf_loop[65].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[65].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_180_),
    .GATE_N(net34),
    .RESET_B(net287),
    .Q(\puf_instance.puf_loop[65].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[66].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_181_),
    .GATE_N(net35),
    .RESET_B(net288),
    .Q(\puf_instance.puf_loop[66].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[66].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_182_),
    .GATE_N(net35),
    .RESET_B(net289),
    .Q(\puf_instance.puf_loop[66].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[67].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_183_),
    .GATE_N(net17),
    .RESET_B(net290),
    .Q(\puf_instance.puf_loop[67].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[67].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_184_),
    .GATE_N(net17),
    .RESET_B(net291),
    .Q(\puf_instance.puf_loop[67].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[68].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_185_),
    .GATE_N(net17),
    .RESET_B(net292),
    .Q(\puf_instance.puf_loop[68].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[68].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_186_),
    .GATE_N(net17),
    .RESET_B(net293),
    .Q(\puf_instance.puf_loop[68].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[69].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_187_),
    .GATE_N(net19),
    .RESET_B(net294),
    .Q(\puf_instance.puf_loop[69].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[69].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_188_),
    .GATE_N(net19),
    .RESET_B(net295),
    .Q(\puf_instance.puf_loop[69].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[6].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_189_),
    .GATE_N(net44),
    .RESET_B(net296),
    .Q(\puf_instance.puf_loop[6].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[6].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_190_),
    .GATE_N(net49),
    .RESET_B(net297),
    .Q(\puf_instance.puf_loop[6].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[70].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_191_),
    .GATE_N(net19),
    .RESET_B(net298),
    .Q(\puf_instance.puf_loop[70].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[70].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_192_),
    .GATE_N(net19),
    .RESET_B(net299),
    .Q(\puf_instance.puf_loop[70].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[71].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_193_),
    .GATE_N(net37),
    .RESET_B(net300),
    .Q(\puf_instance.puf_loop[71].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[71].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_194_),
    .GATE_N(net37),
    .RESET_B(net301),
    .Q(\puf_instance.puf_loop[71].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[72].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_195_),
    .GATE_N(net38),
    .RESET_B(net302),
    .Q(\puf_instance.puf_loop[72].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[72].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_196_),
    .GATE_N(net38),
    .RESET_B(net303),
    .Q(\puf_instance.puf_loop[72].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[73].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_197_),
    .GATE_N(net35),
    .RESET_B(net304),
    .Q(\puf_instance.puf_loop[73].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[73].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_198_),
    .GATE_N(net35),
    .RESET_B(net305),
    .Q(\puf_instance.puf_loop[73].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[74].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_199_),
    .GATE_N(net35),
    .RESET_B(net306),
    .Q(\puf_instance.puf_loop[74].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[74].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_200_),
    .GATE_N(net35),
    .RESET_B(net307),
    .Q(\puf_instance.puf_loop[74].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[75].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_201_),
    .GATE_N(net17),
    .RESET_B(net308),
    .Q(\puf_instance.puf_loop[75].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[75].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_202_),
    .GATE_N(net17),
    .RESET_B(net309),
    .Q(\puf_instance.puf_loop[75].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[76].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_203_),
    .GATE_N(net16),
    .RESET_B(net310),
    .Q(\puf_instance.puf_loop[76].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[76].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_204_),
    .GATE_N(net16),
    .RESET_B(net311),
    .Q(\puf_instance.puf_loop[76].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[77].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_205_),
    .GATE_N(net16),
    .RESET_B(net312),
    .Q(\puf_instance.puf_loop[77].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[77].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_206_),
    .GATE_N(net16),
    .RESET_B(net313),
    .Q(\puf_instance.puf_loop[77].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[78].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_207_),
    .GATE_N(net18),
    .RESET_B(net314),
    .Q(\puf_instance.puf_loop[78].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[78].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_208_),
    .GATE_N(net18),
    .RESET_B(net315),
    .Q(\puf_instance.puf_loop[78].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[79].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_209_),
    .GATE_N(net38),
    .RESET_B(net316),
    .Q(\puf_instance.puf_loop[79].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[79].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_210_),
    .GATE_N(net38),
    .RESET_B(net317),
    .Q(\puf_instance.puf_loop[79].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[7].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_211_),
    .GATE_N(net49),
    .RESET_B(net318),
    .Q(\puf_instance.puf_loop[7].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[7].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_212_),
    .GATE_N(net49),
    .RESET_B(net319),
    .Q(\puf_instance.puf_loop[7].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[80].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_213_),
    .GATE_N(net37),
    .RESET_B(net320),
    .Q(\puf_instance.puf_loop[80].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[80].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_214_),
    .GATE_N(net36),
    .RESET_B(net321),
    .Q(\puf_instance.puf_loop[80].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[81].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_215_),
    .GATE_N(net35),
    .RESET_B(net322),
    .Q(\puf_instance.puf_loop[81].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[81].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_216_),
    .GATE_N(net35),
    .RESET_B(net323),
    .Q(\puf_instance.puf_loop[81].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[82].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_217_),
    .GATE_N(net15),
    .RESET_B(net324),
    .Q(\puf_instance.puf_loop[82].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[82].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_218_),
    .GATE_N(net15),
    .RESET_B(net325),
    .Q(\puf_instance.puf_loop[82].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[83].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_219_),
    .GATE_N(net15),
    .RESET_B(net326),
    .Q(\puf_instance.puf_loop[83].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[83].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_220_),
    .GATE_N(net15),
    .RESET_B(net327),
    .Q(\puf_instance.puf_loop[83].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[84].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_221_),
    .GATE_N(net15),
    .RESET_B(net328),
    .Q(\puf_instance.puf_loop[84].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[84].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_222_),
    .GATE_N(net15),
    .RESET_B(net329),
    .Q(\puf_instance.puf_loop[84].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[85].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_223_),
    .GATE_N(net15),
    .RESET_B(net330),
    .Q(\puf_instance.puf_loop[85].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[85].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_224_),
    .GATE_N(net15),
    .RESET_B(net331),
    .Q(\puf_instance.puf_loop[85].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[86].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_225_),
    .GATE_N(net14),
    .RESET_B(net332),
    .Q(\puf_instance.puf_loop[86].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[86].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_226_),
    .GATE_N(net14),
    .RESET_B(net333),
    .Q(\puf_instance.puf_loop[86].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[87].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_227_),
    .GATE_N(net38),
    .RESET_B(net334),
    .Q(\puf_instance.puf_loop[87].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[87].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_228_),
    .GATE_N(net38),
    .RESET_B(net335),
    .Q(\puf_instance.puf_loop[87].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[88].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_229_),
    .GATE_N(net36),
    .RESET_B(net336),
    .Q(\puf_instance.puf_loop[88].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[88].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_230_),
    .GATE_N(net36),
    .RESET_B(net337),
    .Q(\puf_instance.puf_loop[88].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[89].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_231_),
    .GATE_N(net34),
    .RESET_B(net338),
    .Q(\puf_instance.puf_loop[89].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[89].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_232_),
    .GATE_N(net34),
    .RESET_B(net339),
    .Q(\puf_instance.puf_loop[89].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[8].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_233_),
    .GATE_N(net38),
    .RESET_B(net340),
    .Q(\puf_instance.puf_loop[8].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[8].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_234_),
    .GATE_N(net38),
    .RESET_B(net341),
    .Q(\puf_instance.puf_loop[8].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[90].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_235_),
    .GATE_N(net34),
    .RESET_B(net342),
    .Q(\puf_instance.puf_loop[90].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[90].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_236_),
    .GATE_N(net34),
    .RESET_B(net343),
    .Q(\puf_instance.puf_loop[90].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[91].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_237_),
    .GATE_N(net17),
    .RESET_B(net344),
    .Q(\puf_instance.puf_loop[91].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[91].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_238_),
    .GATE_N(net17),
    .RESET_B(net345),
    .Q(\puf_instance.puf_loop[91].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[92].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_239_),
    .GATE_N(net16),
    .RESET_B(net346),
    .Q(\puf_instance.puf_loop[92].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[92].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_240_),
    .GATE_N(net16),
    .RESET_B(net347),
    .Q(\puf_instance.puf_loop[92].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[93].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_241_),
    .GATE_N(net16),
    .RESET_B(net348),
    .Q(\puf_instance.puf_loop[93].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[93].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_242_),
    .GATE_N(net16),
    .RESET_B(net349),
    .Q(\puf_instance.puf_loop[93].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[94].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_243_),
    .GATE_N(net18),
    .RESET_B(net350),
    .Q(\puf_instance.puf_loop[94].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[94].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_244_),
    .GATE_N(net18),
    .RESET_B(net351),
    .Q(\puf_instance.puf_loop[94].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[95].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_245_),
    .GATE_N(net37),
    .RESET_B(net352),
    .Q(\puf_instance.puf_loop[95].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[95].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_246_),
    .GATE_N(net37),
    .RESET_B(net353),
    .Q(\puf_instance.puf_loop[95].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[96].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_247_),
    .GATE_N(net42),
    .RESET_B(net354),
    .Q(\puf_instance.puf_loop[96].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[96].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_248_),
    .GATE_N(net42),
    .RESET_B(net355),
    .Q(\puf_instance.puf_loop[96].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[97].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_249_),
    .GATE_N(net40),
    .RESET_B(net356),
    .Q(\puf_instance.puf_loop[97].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[97].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_250_),
    .GATE_N(net40),
    .RESET_B(net357),
    .Q(\puf_instance.puf_loop[97].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[98].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_251_),
    .GATE_N(net41),
    .RESET_B(net358),
    .Q(\puf_instance.puf_loop[98].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[98].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_252_),
    .GATE_N(net41),
    .RESET_B(net359),
    .Q(\puf_instance.puf_loop[98].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[99].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_253_),
    .GATE_N(net43),
    .RESET_B(net360),
    .Q(\puf_instance.puf_loop[99].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[99].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_254_),
    .GATE_N(net43),
    .RESET_B(net361),
    .Q(\puf_instance.puf_loop[99].puf_inst.Q1 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[9].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_255_),
    .GATE_N(net49),
    .RESET_B(net362),
    .Q(\puf_instance.puf_loop[9].puf_inst.Q0 ));
 sg13g2_dllrq_1 \puf_instance.puf_loop[9].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_256_),
    .GATE_N(net49),
    .RESET_B(net363),
    .Q(\puf_instance.puf_loop[9].puf_inst.Q1 ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[2]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[4]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[7]));
 sg13g2_buf_1 fanout13 (.A(net22),
    .X(net13));
 sg13g2_buf_1 fanout14 (.A(net22),
    .X(net14));
 sg13g2_buf_1 fanout15 (.A(net22),
    .X(net15));
 sg13g2_buf_1 fanout16 (.A(net21),
    .X(net16));
 sg13g2_buf_1 fanout17 (.A(net21),
    .X(net17));
 sg13g2_buf_1 fanout18 (.A(net20),
    .X(net18));
 sg13g2_buf_1 fanout19 (.A(net21),
    .X(net19));
 sg13g2_buf_1 fanout20 (.A(net21),
    .X(net20));
 sg13g2_buf_1 fanout21 (.A(net22),
    .X(net21));
 sg13g2_buf_1 fanout22 (.A(net56),
    .X(net22));
 sg13g2_buf_1 fanout23 (.A(net28),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(net28),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(net26),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(net56),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(net33),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net33),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net33),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net56),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net36),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net39),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(net39),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(net39),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net55),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net45),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net45),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net45),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net55),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net48),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(net55),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net54),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(net54),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net54),
    .X(net52));
 sg13g2_buf_1 fanout53 (.A(net54),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(net56),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(_001_),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(_354_),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(_353_),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(_352_),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(_351_),
    .X(net60));
 sg13g2_buf_1 fanout61 (.A(_350_),
    .X(net61));
 sg13g2_buf_1 fanout62 (.A(_349_),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(_348_),
    .X(net63));
 sg13g2_buf_1 fanout64 (.A(_347_),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(_346_),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(_345_),
    .X(net66));
 sg13g2_buf_1 fanout67 (.A(_343_),
    .X(net67));
 sg13g2_buf_1 fanout68 (.A(_342_),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(_341_),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(_340_),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(_339_),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(_338_),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(_337_),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(_336_),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(_335_),
    .X(net75));
 sg13g2_buf_1 fanout76 (.A(_334_),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(_332_),
    .X(net77));
 sg13g2_buf_1 fanout78 (.A(_331_),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(_330_),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(_356_),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(_355_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_344_),
    .X(net82));
 sg13g2_buf_1 fanout83 (.A(_333_),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(_329_),
    .X(net84));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_281_));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_280_));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(_273_));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_272_));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(_268_));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(_266_));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net1));
 sg13g2_tielo _726__92 (.L_LO(net92));
 sg13g2_tielo _727__93 (.L_LO(net93));
 sg13g2_tielo _728__94 (.L_LO(net94));
 sg13g2_tielo _729__95 (.L_LO(net95));
 sg13g2_tielo _730__96 (.L_LO(net96));
 sg13g2_tielo _731__97 (.L_LO(net97));
 sg13g2_tielo _732__98 (.L_LO(net98));
 sg13g2_tielo _733__99 (.L_LO(net99));
 sg13g2_tielo _734__100 (.L_LO(net100));
 sg13g2_tielo _735__101 (.L_LO(net101));
 sg13g2_tielo _736__102 (.L_LO(net102));
 sg13g2_tielo _737__103 (.L_LO(net103));
 sg13g2_tielo _738__104 (.L_LO(net104));
 sg13g2_tielo _739__105 (.L_LO(net105));
 sg13g2_tielo _740__106 (.L_LO(net106));
 sg13g2_tielo _741__107 (.L_LO(net107));
 sg13g2_tiehi \puf_instance.puf_loop[0].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_109  (.L_HI(net109));
 sg13g2_tiehi \puf_instance.puf_loop[100].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_110  (.L_HI(net110));
 sg13g2_tiehi \puf_instance.puf_loop[100].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_111  (.L_HI(net111));
 sg13g2_tiehi \puf_instance.puf_loop[101].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_112  (.L_HI(net112));
 sg13g2_tiehi \puf_instance.puf_loop[101].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_113  (.L_HI(net113));
 sg13g2_tiehi \puf_instance.puf_loop[102].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_114  (.L_HI(net114));
 sg13g2_tiehi \puf_instance.puf_loop[102].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_115  (.L_HI(net115));
 sg13g2_tiehi \puf_instance.puf_loop[103].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_116  (.L_HI(net116));
 sg13g2_tiehi \puf_instance.puf_loop[103].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_117  (.L_HI(net117));
 sg13g2_tiehi \puf_instance.puf_loop[104].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_118  (.L_HI(net118));
 sg13g2_tiehi \puf_instance.puf_loop[104].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_119  (.L_HI(net119));
 sg13g2_tiehi \puf_instance.puf_loop[105].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_120  (.L_HI(net120));
 sg13g2_tiehi \puf_instance.puf_loop[105].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_121  (.L_HI(net121));
 sg13g2_tiehi \puf_instance.puf_loop[106].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_122  (.L_HI(net122));
 sg13g2_tiehi \puf_instance.puf_loop[106].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_123  (.L_HI(net123));
 sg13g2_tiehi \puf_instance.puf_loop[107].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_124  (.L_HI(net124));
 sg13g2_tiehi \puf_instance.puf_loop[107].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_125  (.L_HI(net125));
 sg13g2_tiehi \puf_instance.puf_loop[108].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_126  (.L_HI(net126));
 sg13g2_tiehi \puf_instance.puf_loop[108].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_127  (.L_HI(net127));
 sg13g2_tiehi \puf_instance.puf_loop[109].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_128  (.L_HI(net128));
 sg13g2_tiehi \puf_instance.puf_loop[109].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_129  (.L_HI(net129));
 sg13g2_tiehi \puf_instance.puf_loop[10].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_130  (.L_HI(net130));
 sg13g2_tiehi \puf_instance.puf_loop[10].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_131  (.L_HI(net131));
 sg13g2_tiehi \puf_instance.puf_loop[110].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_132  (.L_HI(net132));
 sg13g2_tiehi \puf_instance.puf_loop[110].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_133  (.L_HI(net133));
 sg13g2_tiehi \puf_instance.puf_loop[111].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_134  (.L_HI(net134));
 sg13g2_tiehi \puf_instance.puf_loop[111].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_135  (.L_HI(net135));
 sg13g2_tiehi \puf_instance.puf_loop[112].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_136  (.L_HI(net136));
 sg13g2_tiehi \puf_instance.puf_loop[112].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_137  (.L_HI(net137));
 sg13g2_tiehi \puf_instance.puf_loop[113].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_138  (.L_HI(net138));
 sg13g2_tiehi \puf_instance.puf_loop[113].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_139  (.L_HI(net139));
 sg13g2_tiehi \puf_instance.puf_loop[114].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_140  (.L_HI(net140));
 sg13g2_tiehi \puf_instance.puf_loop[114].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_141  (.L_HI(net141));
 sg13g2_tiehi \puf_instance.puf_loop[115].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_142  (.L_HI(net142));
 sg13g2_tiehi \puf_instance.puf_loop[115].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_143  (.L_HI(net143));
 sg13g2_tiehi \puf_instance.puf_loop[116].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_144  (.L_HI(net144));
 sg13g2_tiehi \puf_instance.puf_loop[116].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_145  (.L_HI(net145));
 sg13g2_tiehi \puf_instance.puf_loop[117].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_146  (.L_HI(net146));
 sg13g2_tiehi \puf_instance.puf_loop[117].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_147  (.L_HI(net147));
 sg13g2_tiehi \puf_instance.puf_loop[118].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_148  (.L_HI(net148));
 sg13g2_tiehi \puf_instance.puf_loop[118].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_149  (.L_HI(net149));
 sg13g2_tiehi \puf_instance.puf_loop[119].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_150  (.L_HI(net150));
 sg13g2_tiehi \puf_instance.puf_loop[119].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_151  (.L_HI(net151));
 sg13g2_tiehi \puf_instance.puf_loop[11].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_152  (.L_HI(net152));
 sg13g2_tiehi \puf_instance.puf_loop[11].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_153  (.L_HI(net153));
 sg13g2_tiehi \puf_instance.puf_loop[120].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_154  (.L_HI(net154));
 sg13g2_tiehi \puf_instance.puf_loop[120].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_155  (.L_HI(net155));
 sg13g2_tiehi \puf_instance.puf_loop[121].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_156  (.L_HI(net156));
 sg13g2_tiehi \puf_instance.puf_loop[121].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_157  (.L_HI(net157));
 sg13g2_tiehi \puf_instance.puf_loop[122].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_158  (.L_HI(net158));
 sg13g2_tiehi \puf_instance.puf_loop[122].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_159  (.L_HI(net159));
 sg13g2_tiehi \puf_instance.puf_loop[123].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_160  (.L_HI(net160));
 sg13g2_tiehi \puf_instance.puf_loop[123].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_161  (.L_HI(net161));
 sg13g2_tiehi \puf_instance.puf_loop[124].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_162  (.L_HI(net162));
 sg13g2_tiehi \puf_instance.puf_loop[124].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_163  (.L_HI(net163));
 sg13g2_tiehi \puf_instance.puf_loop[125].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_164  (.L_HI(net164));
 sg13g2_tiehi \puf_instance.puf_loop[125].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_165  (.L_HI(net165));
 sg13g2_tiehi \puf_instance.puf_loop[126].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_166  (.L_HI(net166));
 sg13g2_tiehi \puf_instance.puf_loop[126].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_167  (.L_HI(net167));
 sg13g2_tiehi \puf_instance.puf_loop[127].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_168  (.L_HI(net168));
 sg13g2_tiehi \puf_instance.puf_loop[127].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_169  (.L_HI(net169));
 sg13g2_tiehi \puf_instance.puf_loop[12].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_170  (.L_HI(net170));
 sg13g2_tiehi \puf_instance.puf_loop[12].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_171  (.L_HI(net171));
 sg13g2_tiehi \puf_instance.puf_loop[13].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_172  (.L_HI(net172));
 sg13g2_tiehi \puf_instance.puf_loop[13].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_173  (.L_HI(net173));
 sg13g2_tiehi \puf_instance.puf_loop[14].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_174  (.L_HI(net174));
 sg13g2_tiehi \puf_instance.puf_loop[14].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_175  (.L_HI(net175));
 sg13g2_tiehi \puf_instance.puf_loop[15].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_176  (.L_HI(net176));
 sg13g2_tiehi \puf_instance.puf_loop[15].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_177  (.L_HI(net177));
 sg13g2_tiehi \puf_instance.puf_loop[16].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_178  (.L_HI(net178));
 sg13g2_tiehi \puf_instance.puf_loop[16].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_179  (.L_HI(net179));
 sg13g2_tiehi \puf_instance.puf_loop[17].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_180  (.L_HI(net180));
 sg13g2_tiehi \puf_instance.puf_loop[17].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_181  (.L_HI(net181));
 sg13g2_tiehi \puf_instance.puf_loop[18].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_182  (.L_HI(net182));
 sg13g2_tiehi \puf_instance.puf_loop[18].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_183  (.L_HI(net183));
 sg13g2_tiehi \puf_instance.puf_loop[19].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_184  (.L_HI(net184));
 sg13g2_tiehi \puf_instance.puf_loop[19].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_185  (.L_HI(net185));
 sg13g2_tiehi \puf_instance.puf_loop[1].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_186  (.L_HI(net186));
 sg13g2_tiehi \puf_instance.puf_loop[1].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_187  (.L_HI(net187));
 sg13g2_tiehi \puf_instance.puf_loop[20].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_188  (.L_HI(net188));
 sg13g2_tiehi \puf_instance.puf_loop[20].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_189  (.L_HI(net189));
 sg13g2_tiehi \puf_instance.puf_loop[21].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_190  (.L_HI(net190));
 sg13g2_tiehi \puf_instance.puf_loop[21].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_191  (.L_HI(net191));
 sg13g2_tiehi \puf_instance.puf_loop[22].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_192  (.L_HI(net192));
 sg13g2_tiehi \puf_instance.puf_loop[22].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_193  (.L_HI(net193));
 sg13g2_tiehi \puf_instance.puf_loop[23].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_194  (.L_HI(net194));
 sg13g2_tiehi \puf_instance.puf_loop[23].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_195  (.L_HI(net195));
 sg13g2_tiehi \puf_instance.puf_loop[24].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_196  (.L_HI(net196));
 sg13g2_tiehi \puf_instance.puf_loop[24].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_197  (.L_HI(net197));
 sg13g2_tiehi \puf_instance.puf_loop[25].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_198  (.L_HI(net198));
 sg13g2_tiehi \puf_instance.puf_loop[25].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_199  (.L_HI(net199));
 sg13g2_tiehi \puf_instance.puf_loop[26].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_200  (.L_HI(net200));
 sg13g2_tiehi \puf_instance.puf_loop[26].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_201  (.L_HI(net201));
 sg13g2_tiehi \puf_instance.puf_loop[27].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_202  (.L_HI(net202));
 sg13g2_tiehi \puf_instance.puf_loop[27].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_203  (.L_HI(net203));
 sg13g2_tiehi \puf_instance.puf_loop[28].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_204  (.L_HI(net204));
 sg13g2_tiehi \puf_instance.puf_loop[28].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_205  (.L_HI(net205));
 sg13g2_tiehi \puf_instance.puf_loop[29].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_206  (.L_HI(net206));
 sg13g2_tiehi \puf_instance.puf_loop[29].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_207  (.L_HI(net207));
 sg13g2_tiehi \puf_instance.puf_loop[2].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_208  (.L_HI(net208));
 sg13g2_tiehi \puf_instance.puf_loop[2].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_209  (.L_HI(net209));
 sg13g2_tiehi \puf_instance.puf_loop[30].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_210  (.L_HI(net210));
 sg13g2_tiehi \puf_instance.puf_loop[30].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_211  (.L_HI(net211));
 sg13g2_tiehi \puf_instance.puf_loop[31].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_212  (.L_HI(net212));
 sg13g2_tiehi \puf_instance.puf_loop[31].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_213  (.L_HI(net213));
 sg13g2_tiehi \puf_instance.puf_loop[32].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_214  (.L_HI(net214));
 sg13g2_tiehi \puf_instance.puf_loop[32].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_215  (.L_HI(net215));
 sg13g2_tiehi \puf_instance.puf_loop[33].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_216  (.L_HI(net216));
 sg13g2_tiehi \puf_instance.puf_loop[33].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_217  (.L_HI(net217));
 sg13g2_tiehi \puf_instance.puf_loop[34].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_218  (.L_HI(net218));
 sg13g2_tiehi \puf_instance.puf_loop[34].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_219  (.L_HI(net219));
 sg13g2_tiehi \puf_instance.puf_loop[35].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_220  (.L_HI(net220));
 sg13g2_tiehi \puf_instance.puf_loop[35].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_221  (.L_HI(net221));
 sg13g2_tiehi \puf_instance.puf_loop[36].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_222  (.L_HI(net222));
 sg13g2_tiehi \puf_instance.puf_loop[36].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_223  (.L_HI(net223));
 sg13g2_tiehi \puf_instance.puf_loop[37].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_224  (.L_HI(net224));
 sg13g2_tiehi \puf_instance.puf_loop[37].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_225  (.L_HI(net225));
 sg13g2_tiehi \puf_instance.puf_loop[38].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_226  (.L_HI(net226));
 sg13g2_tiehi \puf_instance.puf_loop[38].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_227  (.L_HI(net227));
 sg13g2_tiehi \puf_instance.puf_loop[39].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_228  (.L_HI(net228));
 sg13g2_tiehi \puf_instance.puf_loop[39].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_229  (.L_HI(net229));
 sg13g2_tiehi \puf_instance.puf_loop[3].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_230  (.L_HI(net230));
 sg13g2_tiehi \puf_instance.puf_loop[3].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_231  (.L_HI(net231));
 sg13g2_tiehi \puf_instance.puf_loop[40].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_232  (.L_HI(net232));
 sg13g2_tiehi \puf_instance.puf_loop[40].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_233  (.L_HI(net233));
 sg13g2_tiehi \puf_instance.puf_loop[41].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_234  (.L_HI(net234));
 sg13g2_tiehi \puf_instance.puf_loop[41].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_235  (.L_HI(net235));
 sg13g2_tiehi \puf_instance.puf_loop[42].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_236  (.L_HI(net236));
 sg13g2_tiehi \puf_instance.puf_loop[42].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_237  (.L_HI(net237));
 sg13g2_tiehi \puf_instance.puf_loop[43].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_238  (.L_HI(net238));
 sg13g2_tiehi \puf_instance.puf_loop[43].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_239  (.L_HI(net239));
 sg13g2_tiehi \puf_instance.puf_loop[44].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_240  (.L_HI(net240));
 sg13g2_tiehi \puf_instance.puf_loop[44].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_241  (.L_HI(net241));
 sg13g2_tiehi \puf_instance.puf_loop[45].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_242  (.L_HI(net242));
 sg13g2_tiehi \puf_instance.puf_loop[45].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_243  (.L_HI(net243));
 sg13g2_tiehi \puf_instance.puf_loop[46].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_244  (.L_HI(net244));
 sg13g2_tiehi \puf_instance.puf_loop[46].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_245  (.L_HI(net245));
 sg13g2_tiehi \puf_instance.puf_loop[47].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_246  (.L_HI(net246));
 sg13g2_tiehi \puf_instance.puf_loop[47].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_247  (.L_HI(net247));
 sg13g2_tiehi \puf_instance.puf_loop[48].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_248  (.L_HI(net248));
 sg13g2_tiehi \puf_instance.puf_loop[48].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_249  (.L_HI(net249));
 sg13g2_tiehi \puf_instance.puf_loop[49].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_250  (.L_HI(net250));
 sg13g2_tiehi \puf_instance.puf_loop[49].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_251  (.L_HI(net251));
 sg13g2_tiehi \puf_instance.puf_loop[4].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_252  (.L_HI(net252));
 sg13g2_tiehi \puf_instance.puf_loop[4].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_253  (.L_HI(net253));
 sg13g2_tiehi \puf_instance.puf_loop[50].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_254  (.L_HI(net254));
 sg13g2_tiehi \puf_instance.puf_loop[50].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_255  (.L_HI(net255));
 sg13g2_tiehi \puf_instance.puf_loop[51].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_256  (.L_HI(net256));
 sg13g2_tiehi \puf_instance.puf_loop[51].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_257  (.L_HI(net257));
 sg13g2_tiehi \puf_instance.puf_loop[52].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_258  (.L_HI(net258));
 sg13g2_tiehi \puf_instance.puf_loop[52].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_259  (.L_HI(net259));
 sg13g2_tiehi \puf_instance.puf_loop[53].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_260  (.L_HI(net260));
 sg13g2_tiehi \puf_instance.puf_loop[53].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_261  (.L_HI(net261));
 sg13g2_tiehi \puf_instance.puf_loop[54].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_262  (.L_HI(net262));
 sg13g2_tiehi \puf_instance.puf_loop[54].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_263  (.L_HI(net263));
 sg13g2_tiehi \puf_instance.puf_loop[55].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_264  (.L_HI(net264));
 sg13g2_tiehi \puf_instance.puf_loop[55].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_265  (.L_HI(net265));
 sg13g2_tiehi \puf_instance.puf_loop[56].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_266  (.L_HI(net266));
 sg13g2_tiehi \puf_instance.puf_loop[56].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_267  (.L_HI(net267));
 sg13g2_tiehi \puf_instance.puf_loop[57].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_268  (.L_HI(net268));
 sg13g2_tiehi \puf_instance.puf_loop[57].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_269  (.L_HI(net269));
 sg13g2_tiehi \puf_instance.puf_loop[58].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_270  (.L_HI(net270));
 sg13g2_tiehi \puf_instance.puf_loop[58].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_271  (.L_HI(net271));
 sg13g2_tiehi \puf_instance.puf_loop[59].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_272  (.L_HI(net272));
 sg13g2_tiehi \puf_instance.puf_loop[59].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_273  (.L_HI(net273));
 sg13g2_tiehi \puf_instance.puf_loop[5].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_274  (.L_HI(net274));
 sg13g2_tiehi \puf_instance.puf_loop[5].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_275  (.L_HI(net275));
 sg13g2_tiehi \puf_instance.puf_loop[60].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_276  (.L_HI(net276));
 sg13g2_tiehi \puf_instance.puf_loop[60].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_277  (.L_HI(net277));
 sg13g2_tiehi \puf_instance.puf_loop[61].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_278  (.L_HI(net278));
 sg13g2_tiehi \puf_instance.puf_loop[61].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_279  (.L_HI(net279));
 sg13g2_tiehi \puf_instance.puf_loop[62].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_280  (.L_HI(net280));
 sg13g2_tiehi \puf_instance.puf_loop[62].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_281  (.L_HI(net281));
 sg13g2_tiehi \puf_instance.puf_loop[63].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_282  (.L_HI(net282));
 sg13g2_tiehi \puf_instance.puf_loop[63].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_283  (.L_HI(net283));
 sg13g2_tiehi \puf_instance.puf_loop[64].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_284  (.L_HI(net284));
 sg13g2_tiehi \puf_instance.puf_loop[64].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_285  (.L_HI(net285));
 sg13g2_tiehi \puf_instance.puf_loop[65].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_286  (.L_HI(net286));
 sg13g2_tiehi \puf_instance.puf_loop[65].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_287  (.L_HI(net287));
 sg13g2_tiehi \puf_instance.puf_loop[66].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_288  (.L_HI(net288));
 sg13g2_tiehi \puf_instance.puf_loop[66].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_289  (.L_HI(net289));
 sg13g2_tiehi \puf_instance.puf_loop[67].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_290  (.L_HI(net290));
 sg13g2_tiehi \puf_instance.puf_loop[67].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_291  (.L_HI(net291));
 sg13g2_tiehi \puf_instance.puf_loop[68].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_292  (.L_HI(net292));
 sg13g2_tiehi \puf_instance.puf_loop[68].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_293  (.L_HI(net293));
 sg13g2_tiehi \puf_instance.puf_loop[69].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_294  (.L_HI(net294));
 sg13g2_tiehi \puf_instance.puf_loop[69].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_295  (.L_HI(net295));
 sg13g2_tiehi \puf_instance.puf_loop[6].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_296  (.L_HI(net296));
 sg13g2_tiehi \puf_instance.puf_loop[6].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_297  (.L_HI(net297));
 sg13g2_tiehi \puf_instance.puf_loop[70].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_298  (.L_HI(net298));
 sg13g2_tiehi \puf_instance.puf_loop[70].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_299  (.L_HI(net299));
 sg13g2_tiehi \puf_instance.puf_loop[71].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_300  (.L_HI(net300));
 sg13g2_tiehi \puf_instance.puf_loop[71].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_301  (.L_HI(net301));
 sg13g2_tiehi \puf_instance.puf_loop[72].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_302  (.L_HI(net302));
 sg13g2_tiehi \puf_instance.puf_loop[72].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_303  (.L_HI(net303));
 sg13g2_tiehi \puf_instance.puf_loop[73].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_304  (.L_HI(net304));
 sg13g2_tiehi \puf_instance.puf_loop[73].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_305  (.L_HI(net305));
 sg13g2_tiehi \puf_instance.puf_loop[74].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_306  (.L_HI(net306));
 sg13g2_tiehi \puf_instance.puf_loop[74].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_307  (.L_HI(net307));
 sg13g2_tiehi \puf_instance.puf_loop[75].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_308  (.L_HI(net308));
 sg13g2_tiehi \puf_instance.puf_loop[75].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_309  (.L_HI(net309));
 sg13g2_tiehi \puf_instance.puf_loop[76].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_310  (.L_HI(net310));
 sg13g2_tiehi \puf_instance.puf_loop[76].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_311  (.L_HI(net311));
 sg13g2_tiehi \puf_instance.puf_loop[77].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_312  (.L_HI(net312));
 sg13g2_tiehi \puf_instance.puf_loop[77].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_313  (.L_HI(net313));
 sg13g2_tiehi \puf_instance.puf_loop[78].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_314  (.L_HI(net314));
 sg13g2_tiehi \puf_instance.puf_loop[78].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_315  (.L_HI(net315));
 sg13g2_tiehi \puf_instance.puf_loop[79].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_316  (.L_HI(net316));
 sg13g2_tiehi \puf_instance.puf_loop[79].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_317  (.L_HI(net317));
 sg13g2_tiehi \puf_instance.puf_loop[7].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_318  (.L_HI(net318));
 sg13g2_tiehi \puf_instance.puf_loop[7].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_319  (.L_HI(net319));
 sg13g2_tiehi \puf_instance.puf_loop[80].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_320  (.L_HI(net320));
 sg13g2_tiehi \puf_instance.puf_loop[80].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_321  (.L_HI(net321));
 sg13g2_tiehi \puf_instance.puf_loop[81].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_322  (.L_HI(net322));
 sg13g2_tiehi \puf_instance.puf_loop[81].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_323  (.L_HI(net323));
 sg13g2_tiehi \puf_instance.puf_loop[82].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_324  (.L_HI(net324));
 sg13g2_tiehi \puf_instance.puf_loop[82].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_325  (.L_HI(net325));
 sg13g2_tiehi \puf_instance.puf_loop[83].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_326  (.L_HI(net326));
 sg13g2_tiehi \puf_instance.puf_loop[83].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_327  (.L_HI(net327));
 sg13g2_tiehi \puf_instance.puf_loop[84].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_328  (.L_HI(net328));
 sg13g2_tiehi \puf_instance.puf_loop[84].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_329  (.L_HI(net329));
 sg13g2_tiehi \puf_instance.puf_loop[85].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_330  (.L_HI(net330));
 sg13g2_tiehi \puf_instance.puf_loop[85].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_331  (.L_HI(net331));
 sg13g2_tiehi \puf_instance.puf_loop[86].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_332  (.L_HI(net332));
 sg13g2_tiehi \puf_instance.puf_loop[86].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_333  (.L_HI(net333));
 sg13g2_tiehi \puf_instance.puf_loop[87].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_334  (.L_HI(net334));
 sg13g2_tiehi \puf_instance.puf_loop[87].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_335  (.L_HI(net335));
 sg13g2_tiehi \puf_instance.puf_loop[88].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_336  (.L_HI(net336));
 sg13g2_tiehi \puf_instance.puf_loop[88].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_337  (.L_HI(net337));
 sg13g2_tiehi \puf_instance.puf_loop[89].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_338  (.L_HI(net338));
 sg13g2_tiehi \puf_instance.puf_loop[89].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_339  (.L_HI(net339));
 sg13g2_tiehi \puf_instance.puf_loop[8].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_340  (.L_HI(net340));
 sg13g2_tiehi \puf_instance.puf_loop[8].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_341  (.L_HI(net341));
 sg13g2_tiehi \puf_instance.puf_loop[90].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_342  (.L_HI(net342));
 sg13g2_tiehi \puf_instance.puf_loop[90].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_343  (.L_HI(net343));
 sg13g2_tiehi \puf_instance.puf_loop[91].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_344  (.L_HI(net344));
 sg13g2_tiehi \puf_instance.puf_loop[91].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_345  (.L_HI(net345));
 sg13g2_tiehi \puf_instance.puf_loop[92].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_346  (.L_HI(net346));
 sg13g2_tiehi \puf_instance.puf_loop[92].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_347  (.L_HI(net347));
 sg13g2_tiehi \puf_instance.puf_loop[93].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_348  (.L_HI(net348));
 sg13g2_tiehi \puf_instance.puf_loop[93].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_349  (.L_HI(net349));
 sg13g2_tiehi \puf_instance.puf_loop[94].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_350  (.L_HI(net350));
 sg13g2_tiehi \puf_instance.puf_loop[94].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_351  (.L_HI(net351));
 sg13g2_tiehi \puf_instance.puf_loop[95].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_352  (.L_HI(net352));
 sg13g2_tiehi \puf_instance.puf_loop[95].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_353  (.L_HI(net353));
 sg13g2_tiehi \puf_instance.puf_loop[96].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_354  (.L_HI(net354));
 sg13g2_tiehi \puf_instance.puf_loop[96].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_355  (.L_HI(net355));
 sg13g2_tiehi \puf_instance.puf_loop[97].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_356  (.L_HI(net356));
 sg13g2_tiehi \puf_instance.puf_loop[97].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_357  (.L_HI(net357));
 sg13g2_tiehi \puf_instance.puf_loop[98].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_358  (.L_HI(net358));
 sg13g2_tiehi \puf_instance.puf_loop[98].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_359  (.L_HI(net359));
 sg13g2_tiehi \puf_instance.puf_loop[99].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_360  (.L_HI(net360));
 sg13g2_tiehi \puf_instance.puf_loop[99].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_361  (.L_HI(net361));
 sg13g2_tiehi \puf_instance.puf_loop[9].puf_inst.dl0.Q$_DLATCH_N_._TECHMAP_DLATCH_N_362  (.L_HI(net362));
 sg13g2_tiehi \puf_instance.puf_loop[9].puf_inst.dl1.Q$_DLATCH_N_._TECHMAP_DLATCH_N_363  (.L_HI(net363));
 sg13g2_buf_1 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_1 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_fill_1 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_229 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_decap_4 FILLER_9_282 ();
 sg13g2_fill_1 FILLER_9_286 ();
 sg13g2_decap_4 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_8 FILLER_9_404 ();
 sg13g2_decap_8 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_105 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_121 ();
 sg13g2_decap_8 FILLER_11_155 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_decap_8 FILLER_11_211 ();
 sg13g2_decap_4 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_330 ();
 sg13g2_decap_4 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_416 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_4 FILLER_12_123 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_138 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_fill_1 FILLER_12_150 ();
 sg13g2_decap_4 FILLER_12_172 ();
 sg13g2_fill_2 FILLER_12_176 ();
 sg13g2_fill_1 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_4 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_236 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_4 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_371 ();
 sg13g2_decap_4 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_4 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_decap_4 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_4 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_279 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_411 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_4 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_90 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_4 FILLER_14_199 ();
 sg13g2_fill_2 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_decap_4 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_365 ();
 sg13g2_fill_1 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_104 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_115 ();
 sg13g2_decap_8 FILLER_15_122 ();
 sg13g2_decap_8 FILLER_15_129 ();
 sg13g2_decap_4 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_140 ();
 sg13g2_fill_1 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_4 FILLER_15_245 ();
 sg13g2_decap_4 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_350 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_4 FILLER_15_368 ();
 sg13g2_fill_1 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_15_423 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_decap_8 FILLER_16_115 ();
 sg13g2_decap_8 FILLER_16_122 ();
 sg13g2_fill_2 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_131 ();
 sg13g2_fill_2 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_177 ();
 sg13g2_fill_2 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_247 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_345 ();
 sg13g2_fill_1 FILLER_16_347 ();
 sg13g2_decap_4 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_356 ();
 sg13g2_decap_4 FILLER_16_369 ();
 sg13g2_decap_4 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_120 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_decap_8 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_4 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_368 ();
 sg13g2_fill_2 FILLER_17_376 ();
 sg13g2_decap_4 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_decap_4 FILLER_17_426 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_132 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_decap_4 FILLER_18_271 ();
 sg13g2_fill_2 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_395 ();
 sg13g2_fill_1 FILLER_18_397 ();
 sg13g2_fill_2 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_fill_2 FILLER_19_78 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_fill_2 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_decap_8 FILLER_20_150 ();
 sg13g2_decap_4 FILLER_20_157 ();
 sg13g2_decap_4 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_decap_4 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_decap_4 FILLER_21_61 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_86 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_decap_4 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_4 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_396 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_34 ();
 sg13g2_decap_8 FILLER_22_41 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_58 ();
 sg13g2_decap_4 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_fill_2 FILLER_22_87 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_decap_8 FILLER_22_94 ();
 sg13g2_decap_8 FILLER_22_101 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_decap_4 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_4 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_4 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_424 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_17 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_65 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_decap_8 FILLER_23_146 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_234 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_decap_4 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_decap_4 FILLER_24_195 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_24_206 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_decap_4 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_decap_4 FILLER_24_367 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_decap_8 FILLER_24_419 ();
 sg13g2_decap_4 FILLER_24_426 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_20 ();
 sg13g2_fill_1 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_43 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_decap_4 FILLER_25_111 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_decap_4 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_4 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_266 ();
 sg13g2_decap_4 FILLER_25_278 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_decap_4 FILLER_25_395 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_11 ();
 sg13g2_fill_2 FILLER_26_73 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_decap_8 FILLER_26_89 ();
 sg13g2_decap_8 FILLER_26_96 ();
 sg13g2_decap_4 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_107 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_4 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_36 ();
 sg13g2_decap_4 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_decap_8 FILLER_27_86 ();
 sg13g2_decap_8 FILLER_27_93 ();
 sg13g2_decap_8 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_4 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_304 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_decap_4 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_4 FILLER_27_367 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_41 ();
 sg13g2_decap_4 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_139 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_decap_4 FILLER_28_397 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_fill_2 FILLER_28_413 ();
 sg13g2_fill_1 FILLER_28_415 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_44 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_decap_4 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_decap_8 FILLER_29_299 ();
 sg13g2_fill_2 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_4 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_fill_1 FILLER_30_19 ();
 sg13g2_decap_8 FILLER_30_40 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_decap_4 FILLER_30_106 ();
 sg13g2_fill_2 FILLER_30_131 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_4 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_decap_8 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_decap_4 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_349 ();
 sg13g2_decap_4 FILLER_30_381 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_48 ();
 sg13g2_fill_2 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_4 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_358 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_fill_1 FILLER_31_402 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_11 ();
 sg13g2_fill_1 FILLER_32_43 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_71 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_decap_4 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_43 ();
 sg13g2_decap_4 FILLER_33_48 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_decap_4 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_decap_4 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_167 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_311 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_decap_8 FILLER_33_332 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_355 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_24 ();
 sg13g2_decap_4 FILLER_34_31 ();
 sg13g2_decap_4 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_74 ();
 sg13g2_fill_1 FILLER_34_76 ();
 sg13g2_decap_4 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_4 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_4 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_decap_4 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_384 ();
 sg13g2_decap_4 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_55 ();
 sg13g2_fill_1 FILLER_35_57 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_decap_4 FILLER_35_134 ();
 sg13g2_decap_4 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_fill_2 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_424 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_fill_1 FILLER_36_58 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_2 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_87 ();
 sg13g2_fill_2 FILLER_36_92 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_decap_4 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_202 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_422 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_16 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_fill_1 FILLER_37_47 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_fill_1 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_decap_4 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_121 ();
 sg13g2_decap_4 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_fill_2 FILLER_37_201 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_368 ();
 sg13g2_fill_2 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_4 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_53 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_128 ();
 sg13g2_decap_8 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_167 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_4 FILLER_38_259 ();
 sg13g2_fill_2 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_410 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
