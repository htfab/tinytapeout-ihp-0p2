module tt_um_favoritohjs_scroller (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire clknet_0_clk;
 wire net58;
 wire \bd[0] ;
 wire \bd[1] ;
 wire \bd[2] ;
 wire \color_ditherer.dither ;
 wire \color_ditherer.gin[0] ;
 wire \color_ditherer.gin[1] ;
 wire \color_ditherer.gin[2] ;
 wire \count1[0] ;
 wire \count1[1] ;
 wire \count1[2] ;
 wire \count1b[0] ;
 wire \count1b[1] ;
 wire \count1b[2] ;
 wire \count2[0] ;
 wire \count2[1] ;
 wire \count2b[0] ;
 wire \count2b[1] ;
 wire count2low;
 wire \cutoff1[0] ;
 wire \cutoff1[1] ;
 wire \cutoff1[2] ;
 wire \cutoff1[3] ;
 wire \cutoff1[4] ;
 wire \cutoff2[0] ;
 wire \cutoff2[1] ;
 wire \cutoff2[2] ;
 wire \cutoff2[3] ;
 wire \cutoff2[4] ;
 wire \hcount[0] ;
 wire \hcount[1] ;
 wire \hcount[2] ;
 wire \hcount[3] ;
 wire \hcount[4] ;
 wire \hcount[5] ;
 wire \hcount[6] ;
 wire \hcount[7] ;
 wire \hcount[8] ;
 wire \hcount[9] ;
 wire hsync;
 wire \l1[0] ;
 wire \l1[1] ;
 wire \l1[2] ;
 wire \l1[3] ;
 wire \l2[0] ;
 wire \l2[1] ;
 wire \l2[2] ;
 wire \l2[3] ;
 wire \lfsr1[4] ;
 wire \lfsr1[5] ;
 wire \lfsr1[6] ;
 wire \lfsr1[7] ;
 wire \lfsr1[8] ;
 wire \lfsr1[9] ;
 wire \lfsr1b[0] ;
 wire \lfsr1b[1] ;
 wire \lfsr1b[2] ;
 wire \lfsr1b[3] ;
 wire \lfsr1b[4] ;
 wire \lfsr1b[5] ;
 wire \lfsr1b[6] ;
 wire \lfsr1b[7] ;
 wire \lfsr1b[8] ;
 wire \lfsr1b[9] ;
 wire \lfsr2[4] ;
 wire \lfsr2[5] ;
 wire \lfsr2[6] ;
 wire \lfsr2[7] ;
 wire \lfsr2[8] ;
 wire \lfsr2[9] ;
 wire \lfsr2b[0] ;
 wire \lfsr2b[1] ;
 wire \lfsr2b[2] ;
 wire \lfsr2b[3] ;
 wire \lfsr2b[4] ;
 wire \lfsr2b[5] ;
 wire \lfsr2b[6] ;
 wire \lfsr2b[7] ;
 wire \lfsr2b[8] ;
 wire \lfsr2b[9] ;
 wire vborder1;
 wire vborder2;
 wire \vcount[0] ;
 wire \vcount[1] ;
 wire \vcount[2] ;
 wire \vcount[3] ;
 wire \vcount[4] ;
 wire \vcount[5] ;
 wire \vcount[6] ;
 wire \vcount[7] ;
 wire \vcount[8] ;
 wire \vcount[9] ;
 wire \vga_sync.vga_vsync ;
 wire \vga_sync.xvisible ;
 wire \vga_sync.yvisible ;
 wire \vscheudler1.blockline[0] ;
 wire \vscheudler1.blockline[1] ;
 wire \vscheudler1.blockline[2] ;
 wire \vscheudler1.blockline[3] ;
 wire \vscheudler1.blockline[4] ;
 wire \vscheudler1.started ;
 wire \vscheudler2.blockline[0] ;
 wire \vscheudler2.blockline[1] ;
 wire \vscheudler2.blockline[2] ;
 wire \vscheudler2.blockline[3] ;
 wire \vscheudler2.blockline[4] ;
 wire \vscheudler2.started ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _0673_ (.A(net1),
    .X(_0121_));
 sg13g2_and2_1 _0674_ (.A(\vga_sync.yvisible ),
    .B(\vga_sync.xvisible ),
    .X(_0122_));
 sg13g2_buf_1 _0675_ (.A(_0122_),
    .X(_0123_));
 sg13g2_nand2_1 _0676_ (.Y(_0124_),
    .A(net41),
    .B(net35));
 sg13g2_inv_1 _0677_ (.Y(_0125_),
    .A(\cutoff1[1] ));
 sg13g2_nand2b_1 _0678_ (.Y(_0126_),
    .B(\cutoff1[0] ),
    .A_N(\l1[0] ));
 sg13g2_o21ai_1 _0679_ (.B1(_0126_),
    .Y(_0127_),
    .A1(\l1[1] ),
    .A2(_0125_));
 sg13g2_inv_1 _0680_ (.Y(_0128_),
    .A(\cutoff1[2] ));
 sg13g2_a22oi_1 _0681_ (.Y(_0129_),
    .B1(\l1[1] ),
    .B2(_0125_),
    .A2(\l1[2] ),
    .A1(_0128_));
 sg13g2_inv_1 _0682_ (.Y(_0130_),
    .A(\cutoff1[4] ));
 sg13g2_nand2_1 _0683_ (.Y(_0131_),
    .A(\l1[3] ),
    .B(_0130_));
 sg13g2_inv_1 _0684_ (.Y(_0132_),
    .A(\cutoff1[3] ));
 sg13g2_nand2_1 _0685_ (.Y(_0133_),
    .A(_0132_),
    .B(_0130_));
 sg13g2_nor2_1 _0686_ (.A(_0128_),
    .B(\l1[2] ),
    .Y(_0134_));
 sg13g2_a221oi_1 _0687_ (.B2(_0133_),
    .C1(_0134_),
    .B1(_0131_),
    .A1(_0127_),
    .Y(_0135_),
    .A2(_0129_));
 sg13g2_nor2_1 _0688_ (.A(\count1[1] ),
    .B(\count1[2] ),
    .Y(_0136_));
 sg13g2_nor2_1 _0689_ (.A(vborder1),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_and3_1 _0690_ (.X(_0138_),
    .A(_0132_),
    .B(\l1[3] ),
    .C(_0130_));
 sg13g2_or2_1 _0691_ (.X(_0139_),
    .B(_0138_),
    .A(_0137_));
 sg13g2_or3_1 _0692_ (.A(_0124_),
    .B(_0135_),
    .C(_0139_),
    .X(_0140_));
 sg13g2_inv_1 _0693_ (.Y(_0070_),
    .A(_0140_));
 sg13g2_buf_2 _0694_ (.A(\hcount[6] ),
    .X(_0141_));
 sg13g2_inv_1 _0695_ (.Y(_0142_),
    .A(_0141_));
 sg13g2_buf_8 _0696_ (.A(\hcount[1] ),
    .X(_0143_));
 sg13g2_nor3_1 _0697_ (.A(_0143_),
    .B(\hcount[3] ),
    .C(\hcount[2] ),
    .Y(_0144_));
 sg13g2_buf_2 _0698_ (.A(\hcount[0] ),
    .X(_0145_));
 sg13g2_nor2b_1 _0699_ (.A(_0145_),
    .B_N(\hcount[9] ),
    .Y(_0146_));
 sg13g2_and3_1 _0700_ (.X(_0147_),
    .A(_0142_),
    .B(_0144_),
    .C(_0146_));
 sg13g2_buf_2 _0701_ (.A(_0147_),
    .X(_0148_));
 sg13g2_buf_8 _0702_ (.A(\hcount[7] ),
    .X(_0149_));
 sg13g2_inv_1 _0703_ (.Y(_0150_),
    .A(\hcount[8] ));
 sg13g2_nand2b_1 _0704_ (.Y(_0151_),
    .B(\hcount[5] ),
    .A_N(\hcount[4] ));
 sg13g2_nor3_2 _0705_ (.A(_0149_),
    .B(_0150_),
    .C(_0151_),
    .Y(_0152_));
 sg13g2_nand2_2 _0706_ (.Y(_0153_),
    .A(_0148_),
    .B(_0152_));
 sg13g2_nand2_1 _0707_ (.Y(_0154_),
    .A(net41),
    .B(_0153_));
 sg13g2_buf_1 _0708_ (.A(_0154_),
    .X(_0155_));
 sg13g2_or2_1 _0709_ (.X(_0075_),
    .B(net12),
    .A(_0010_));
 sg13g2_xnor2_1 _0710_ (.Y(_0156_),
    .A(_0143_),
    .B(_0145_));
 sg13g2_nor2_1 _0711_ (.A(net12),
    .B(_0156_),
    .Y(_0076_));
 sg13g2_nand2_1 _0712_ (.Y(_0157_),
    .A(_0143_),
    .B(_0145_));
 sg13g2_xor2_1 _0713_ (.B(_0157_),
    .A(\hcount[2] ),
    .X(_0158_));
 sg13g2_nor2_1 _0714_ (.A(net12),
    .B(_0158_),
    .Y(_0077_));
 sg13g2_nand3_1 _0715_ (.B(_0145_),
    .C(\hcount[2] ),
    .A(_0143_),
    .Y(_0159_));
 sg13g2_xor2_1 _0716_ (.B(_0159_),
    .A(\hcount[3] ),
    .X(_0160_));
 sg13g2_nor2_1 _0717_ (.A(net12),
    .B(_0160_),
    .Y(_0078_));
 sg13g2_inv_1 _0718_ (.Y(_0161_),
    .A(\hcount[4] ));
 sg13g2_nand4_1 _0719_ (.B(_0145_),
    .C(\hcount[3] ),
    .A(_0143_),
    .Y(_0162_),
    .D(\hcount[2] ));
 sg13g2_xnor2_1 _0720_ (.Y(_0163_),
    .A(_0161_),
    .B(_0162_));
 sg13g2_nor2_1 _0721_ (.A(net12),
    .B(_0163_),
    .Y(_0079_));
 sg13g2_nor2_1 _0722_ (.A(_0161_),
    .B(_0162_),
    .Y(_0164_));
 sg13g2_xnor2_1 _0723_ (.Y(_0165_),
    .A(\hcount[5] ),
    .B(_0164_));
 sg13g2_nor2_1 _0724_ (.A(net12),
    .B(_0165_),
    .Y(_0080_));
 sg13g2_nand2_1 _0725_ (.Y(_0166_),
    .A(\hcount[5] ),
    .B(\hcount[4] ));
 sg13g2_nor2_2 _0726_ (.A(_0162_),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_xnor2_1 _0727_ (.Y(_0168_),
    .A(_0141_),
    .B(_0167_));
 sg13g2_nor2_1 _0728_ (.A(net12),
    .B(_0168_),
    .Y(_0081_));
 sg13g2_inv_1 _0729_ (.Y(_0169_),
    .A(_0149_));
 sg13g2_nand2_1 _0730_ (.Y(_0170_),
    .A(_0141_),
    .B(_0167_));
 sg13g2_xnor2_1 _0731_ (.Y(_0171_),
    .A(_0169_),
    .B(_0170_));
 sg13g2_nor2_1 _0732_ (.A(net12),
    .B(_0171_),
    .Y(_0082_));
 sg13g2_nand3_1 _0733_ (.B(_0149_),
    .C(_0167_),
    .A(_0141_),
    .Y(_0172_));
 sg13g2_xnor2_1 _0734_ (.Y(_0173_),
    .A(_0150_),
    .B(_0172_));
 sg13g2_nor2_1 _0735_ (.A(_0155_),
    .B(_0173_),
    .Y(_0083_));
 sg13g2_inv_1 _0736_ (.Y(_0174_),
    .A(\hcount[9] ));
 sg13g2_nand4_1 _0737_ (.B(_0149_),
    .C(\hcount[8] ),
    .A(_0141_),
    .Y(_0175_),
    .D(_0167_));
 sg13g2_xnor2_1 _0738_ (.Y(_0176_),
    .A(_0174_),
    .B(_0175_));
 sg13g2_nor2_1 _0739_ (.A(_0155_),
    .B(_0176_),
    .Y(_0084_));
 sg13g2_and2_1 _0740_ (.A(net41),
    .B(\vga_sync.vga_vsync ),
    .X(_0177_));
 sg13g2_buf_1 _0741_ (.A(_0177_),
    .X(_0178_));
 sg13g2_buf_1 _0742_ (.A(\vscheudler1.started ),
    .X(_0179_));
 sg13g2_buf_8 _0743_ (.A(_0148_),
    .X(_0180_));
 sg13g2_nor2b_1 _0744_ (.A(\hcount[8] ),
    .B_N(_0149_),
    .Y(_0181_));
 sg13g2_nor2b_1 _0745_ (.A(\hcount[5] ),
    .B_N(\hcount[4] ),
    .Y(_0182_));
 sg13g2_and2_1 _0746_ (.A(_0181_),
    .B(_0182_),
    .X(_0183_));
 sg13g2_buf_2 _0747_ (.A(_0183_),
    .X(_0184_));
 sg13g2_buf_8 _0748_ (.A(_0184_),
    .X(_0185_));
 sg13g2_nand3_1 _0749_ (.B(net25),
    .C(net24),
    .A(_0179_),
    .Y(_0186_));
 sg13g2_xor2_1 _0750_ (.B(_0186_),
    .A(\vscheudler1.blockline[0] ),
    .X(_0187_));
 sg13g2_nand2_1 _0751_ (.Y(_0097_),
    .A(net34),
    .B(_0187_));
 sg13g2_nor2_1 _0752_ (.A(\vscheudler1.blockline[1] ),
    .B(\vscheudler1.blockline[0] ),
    .Y(_0188_));
 sg13g2_nand4_1 _0753_ (.B(net25),
    .C(net24),
    .A(_0179_),
    .Y(_0189_),
    .D(_0188_));
 sg13g2_o21ai_1 _0754_ (.B1(\vscheudler1.blockline[1] ),
    .Y(_0190_),
    .A1(\vscheudler1.blockline[0] ),
    .A2(_0186_));
 sg13g2_nand3_1 _0755_ (.B(_0189_),
    .C(_0190_),
    .A(net34),
    .Y(_0098_));
 sg13g2_buf_2 _0756_ (.A(\vscheudler1.blockline[2] ),
    .X(_0191_));
 sg13g2_xor2_1 _0757_ (.B(_0189_),
    .A(_0191_),
    .X(_0192_));
 sg13g2_nand2_1 _0758_ (.Y(_0099_),
    .A(net34),
    .B(_0192_));
 sg13g2_nor3_1 _0759_ (.A(\vscheudler1.blockline[3] ),
    .B(_0191_),
    .C(_0189_),
    .Y(_0193_));
 sg13g2_o21ai_1 _0760_ (.B1(\vscheudler1.blockline[3] ),
    .Y(_0194_),
    .A1(_0191_),
    .A2(_0189_));
 sg13g2_nand3b_1 _0761_ (.B(_0194_),
    .C(net34),
    .Y(_0100_),
    .A_N(_0193_));
 sg13g2_nand2_1 _0762_ (.Y(_0195_),
    .A(\vscheudler1.blockline[4] ),
    .B(_0186_));
 sg13g2_nor4_2 _0763_ (.A(\vscheudler1.blockline[1] ),
    .B(\vscheudler1.blockline[0] ),
    .C(\vscheudler1.blockline[3] ),
    .Y(_0196_),
    .D(_0191_));
 sg13g2_or3_1 _0764_ (.A(_0000_),
    .B(_0186_),
    .C(_0196_),
    .X(_0197_));
 sg13g2_nand2_2 _0765_ (.Y(_0198_),
    .A(_0121_),
    .B(\vga_sync.vga_vsync ));
 sg13g2_buf_1 _0766_ (.A(_0198_),
    .X(_0199_));
 sg13g2_a21oi_1 _0767_ (.A1(_0195_),
    .A2(_0197_),
    .Y(_0101_),
    .B1(net33));
 sg13g2_and2_1 _0768_ (.A(_0000_),
    .B(_0196_),
    .X(_0200_));
 sg13g2_nand4_1 _0769_ (.B(net25),
    .C(net24),
    .A(_0179_),
    .Y(_0201_),
    .D(_0200_));
 sg13g2_o21ai_1 _0770_ (.B1(net34),
    .Y(_0202_),
    .A1(_0007_),
    .A2(_0201_));
 sg13g2_nor4_1 _0771_ (.A(\cutoff1[3] ),
    .B(_0130_),
    .C(\cutoff1[2] ),
    .D(\cutoff1[1] ),
    .Y(_0203_));
 sg13g2_inv_1 _0772_ (.Y(_0204_),
    .A(\cutoff1[0] ));
 sg13g2_o21ai_1 _0773_ (.B1(_0204_),
    .Y(_0205_),
    .A1(_0201_),
    .A2(_0203_));
 sg13g2_nor2b_1 _0774_ (.A(_0202_),
    .B_N(_0205_),
    .Y(_0102_));
 sg13g2_o21ai_1 _0775_ (.B1(\cutoff1[1] ),
    .Y(_0206_),
    .A1(_0204_),
    .A2(_0201_));
 sg13g2_and4_1 _0776_ (.A(_0179_),
    .B(net25),
    .C(net24),
    .D(_0200_),
    .X(_0207_));
 sg13g2_nand3_1 _0777_ (.B(\cutoff1[0] ),
    .C(_0207_),
    .A(_0125_),
    .Y(_0208_));
 sg13g2_a21oi_1 _0778_ (.A1(_0206_),
    .A2(_0208_),
    .Y(_0103_),
    .B1(net33));
 sg13g2_nand2_1 _0779_ (.Y(_0209_),
    .A(\cutoff1[1] ),
    .B(\cutoff1[0] ));
 sg13g2_o21ai_1 _0780_ (.B1(\cutoff1[2] ),
    .Y(_0210_),
    .A1(_0209_),
    .A2(_0201_));
 sg13g2_nand4_1 _0781_ (.B(\cutoff1[1] ),
    .C(\cutoff1[0] ),
    .A(_0128_),
    .Y(_0211_),
    .D(_0207_));
 sg13g2_a21oi_1 _0782_ (.A1(_0210_),
    .A2(_0211_),
    .Y(_0104_),
    .B1(net33));
 sg13g2_inv_1 _0783_ (.Y(_0212_),
    .A(_0179_));
 sg13g2_nand3_1 _0784_ (.B(_0144_),
    .C(_0146_),
    .A(_0142_),
    .Y(_0213_));
 sg13g2_buf_1 _0785_ (.A(_0213_),
    .X(_0214_));
 sg13g2_nand2_2 _0786_ (.Y(_0215_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_and2_1 _0787_ (.A(\cutoff1[0] ),
    .B(_0000_),
    .X(_0216_));
 sg13g2_nand4_1 _0788_ (.B(\cutoff1[1] ),
    .C(_0196_),
    .A(\cutoff1[2] ),
    .Y(_0217_),
    .D(_0216_));
 sg13g2_or4_1 _0789_ (.A(_0212_),
    .B(net27),
    .C(_0215_),
    .D(_0217_),
    .X(_0218_));
 sg13g2_xnor2_1 _0790_ (.Y(_0219_),
    .A(_0132_),
    .B(_0218_));
 sg13g2_nor2_1 _0791_ (.A(net33),
    .B(_0219_),
    .Y(_0105_));
 sg13g2_o21ai_1 _0792_ (.B1(\cutoff1[4] ),
    .Y(_0220_),
    .A1(_0132_),
    .A2(_0218_));
 sg13g2_or3_1 _0793_ (.A(_0132_),
    .B(\cutoff1[4] ),
    .C(_0218_),
    .X(_0221_));
 sg13g2_a21oi_1 _0794_ (.A1(_0220_),
    .A2(_0221_),
    .Y(_0106_),
    .B1(net33));
 sg13g2_inv_1 _0795_ (.Y(_0222_),
    .A(vborder1));
 sg13g2_nand4_1 _0796_ (.B(_0000_),
    .C(net25),
    .A(_0179_),
    .Y(_0223_),
    .D(net24));
 sg13g2_or4_1 _0797_ (.A(\vscheudler1.blockline[1] ),
    .B(\vscheudler1.blockline[3] ),
    .C(_0191_),
    .D(_0223_),
    .X(_0224_));
 sg13g2_nand4_1 _0798_ (.B(\vscheudler1.blockline[0] ),
    .C(\vscheudler1.blockline[3] ),
    .A(\vscheudler1.blockline[1] ),
    .Y(_0225_),
    .D(_0191_));
 sg13g2_o21ai_1 _0799_ (.B1(net34),
    .Y(_0226_),
    .A1(_0223_),
    .A2(_0225_));
 sg13g2_a21oi_1 _0800_ (.A1(_0222_),
    .A2(_0224_),
    .Y(_0107_),
    .B1(_0226_));
 sg13g2_buf_1 _0801_ (.A(\vcount[0] ),
    .X(_0227_));
 sg13g2_inv_1 _0802_ (.Y(_0228_),
    .A(net40));
 sg13g2_nor3_1 _0803_ (.A(\vcount[1] ),
    .B(\vcount[9] ),
    .C(\vcount[8] ),
    .Y(_0229_));
 sg13g2_and2_1 _0804_ (.A(\vcount[4] ),
    .B(\vcount[5] ),
    .X(_0230_));
 sg13g2_buf_1 _0805_ (.A(_0230_),
    .X(_0231_));
 sg13g2_and3_1 _0806_ (.X(_0232_),
    .A(_0228_),
    .B(_0229_),
    .C(_0231_));
 sg13g2_buf_2 _0807_ (.A(\vcount[2] ),
    .X(_0233_));
 sg13g2_inv_1 _0808_ (.Y(_0234_),
    .A(_0233_));
 sg13g2_inv_1 _0809_ (.Y(_0235_),
    .A(\vcount[6] ));
 sg13g2_nor4_1 _0810_ (.A(\vcount[3] ),
    .B(_0234_),
    .C(\vcount[7] ),
    .D(_0235_),
    .Y(_0236_));
 sg13g2_a21oi_1 _0811_ (.A1(_0232_),
    .A2(_0236_),
    .Y(_0237_),
    .B1(_0179_));
 sg13g2_nor2_1 _0812_ (.A(net33),
    .B(_0237_),
    .Y(_0108_));
 sg13g2_buf_1 _0813_ (.A(\vscheudler2.started ),
    .X(_0238_));
 sg13g2_inv_1 _0814_ (.Y(_0239_),
    .A(_0238_));
 sg13g2_or4_1 _0815_ (.A(_0239_),
    .B(\vscheudler2.blockline[0] ),
    .C(net27),
    .D(_0215_),
    .X(_0240_));
 sg13g2_nand3_1 _0816_ (.B(_0180_),
    .C(net24),
    .A(_0238_),
    .Y(_0241_));
 sg13g2_nand2_1 _0817_ (.Y(_0242_),
    .A(\vscheudler2.blockline[0] ),
    .B(_0241_));
 sg13g2_nand3_1 _0818_ (.B(_0240_),
    .C(_0242_),
    .A(net34),
    .Y(_0109_));
 sg13g2_buf_8 _0819_ (.A(\vscheudler2.blockline[1] ),
    .X(_0243_));
 sg13g2_xor2_1 _0820_ (.B(_0240_),
    .A(_0243_),
    .X(_0244_));
 sg13g2_nand2_1 _0821_ (.Y(_0110_),
    .A(_0178_),
    .B(_0244_));
 sg13g2_nor3_1 _0822_ (.A(_0243_),
    .B(\vscheudler2.blockline[0] ),
    .C(\vscheudler2.blockline[2] ),
    .Y(_0245_));
 sg13g2_nand4_1 _0823_ (.B(net25),
    .C(net24),
    .A(_0238_),
    .Y(_0246_),
    .D(_0245_));
 sg13g2_o21ai_1 _0824_ (.B1(\vscheudler2.blockline[2] ),
    .Y(_0247_),
    .A1(_0243_),
    .A2(_0240_));
 sg13g2_nand3_1 _0825_ (.B(_0246_),
    .C(_0247_),
    .A(_0178_),
    .Y(_0111_));
 sg13g2_nand2_1 _0826_ (.Y(_0248_),
    .A(\vscheudler2.blockline[3] ),
    .B(_0246_));
 sg13g2_or3_1 _0827_ (.A(\vscheudler2.blockline[3] ),
    .B(_0001_),
    .C(_0246_),
    .X(_0249_));
 sg13g2_a21oi_1 _0828_ (.A1(_0248_),
    .A2(_0249_),
    .Y(_0112_),
    .B1(net33));
 sg13g2_nand2_1 _0829_ (.Y(_0250_),
    .A(\vscheudler2.blockline[4] ),
    .B(_0241_));
 sg13g2_nor4_2 _0830_ (.A(_0243_),
    .B(\vscheudler2.blockline[0] ),
    .C(\vscheudler2.blockline[3] ),
    .Y(_0251_),
    .D(\vscheudler2.blockline[2] ));
 sg13g2_or3_1 _0831_ (.A(_0001_),
    .B(_0241_),
    .C(_0251_),
    .X(_0252_));
 sg13g2_a21oi_1 _0832_ (.A1(_0250_),
    .A2(_0252_),
    .Y(_0113_),
    .B1(_0198_));
 sg13g2_inv_1 _0833_ (.Y(_0253_),
    .A(\cutoff2[1] ));
 sg13g2_buf_1 _0834_ (.A(\cutoff2[2] ),
    .X(_0254_));
 sg13g2_nor4_1 _0835_ (.A(\cutoff2[0] ),
    .B(\cutoff2[3] ),
    .C(_0254_),
    .D(_0002_),
    .Y(_0255_));
 sg13g2_a21oi_1 _0836_ (.A1(_0253_),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0198_));
 sg13g2_and2_1 _0837_ (.A(_0006_),
    .B(_0256_),
    .X(_0257_));
 sg13g2_and2_1 _0838_ (.A(\cutoff2[0] ),
    .B(net34),
    .X(_0258_));
 sg13g2_nor2_2 _0839_ (.A(net27),
    .B(_0215_),
    .Y(_0259_));
 sg13g2_nand4_1 _0840_ (.B(_0001_),
    .C(_0259_),
    .A(_0238_),
    .Y(_0260_),
    .D(_0251_));
 sg13g2_mux2_1 _0841_ (.A0(_0257_),
    .A1(_0258_),
    .S(_0260_),
    .X(_0114_));
 sg13g2_nand4_1 _0842_ (.B(_0001_),
    .C(_0148_),
    .A(_0238_),
    .Y(_0261_),
    .D(_0184_));
 sg13g2_nand2_1 _0843_ (.Y(_0262_),
    .A(\cutoff2[0] ),
    .B(_0251_));
 sg13g2_nor2_1 _0844_ (.A(_0253_),
    .B(_0198_),
    .Y(_0263_));
 sg13g2_o21ai_1 _0845_ (.B1(_0263_),
    .Y(_0264_),
    .A1(_0261_),
    .A2(_0262_));
 sg13g2_or4_1 _0846_ (.A(\cutoff2[1] ),
    .B(_0198_),
    .C(_0261_),
    .D(_0262_),
    .X(_0265_));
 sg13g2_nand2_1 _0847_ (.Y(_0115_),
    .A(_0264_),
    .B(_0265_));
 sg13g2_inv_1 _0848_ (.Y(_0266_),
    .A(_0254_));
 sg13g2_and4_1 _0849_ (.A(_0001_),
    .B(\cutoff2[1] ),
    .C(\cutoff2[0] ),
    .D(_0251_),
    .X(_0267_));
 sg13g2_nand4_1 _0850_ (.B(_0180_),
    .C(_0185_),
    .A(_0238_),
    .Y(_0268_),
    .D(_0267_));
 sg13g2_xnor2_1 _0851_ (.Y(_0269_),
    .A(_0266_),
    .B(_0268_));
 sg13g2_nor2_1 _0852_ (.A(_0199_),
    .B(_0269_),
    .Y(_0116_));
 sg13g2_o21ai_1 _0853_ (.B1(\cutoff2[3] ),
    .Y(_0270_),
    .A1(_0266_),
    .A2(_0268_));
 sg13g2_or3_1 _0854_ (.A(\cutoff2[3] ),
    .B(_0266_),
    .C(_0268_),
    .X(_0271_));
 sg13g2_a21oi_1 _0855_ (.A1(_0270_),
    .A2(_0271_),
    .Y(_0117_),
    .B1(_0198_));
 sg13g2_buf_1 _0856_ (.A(_0214_),
    .X(_0272_));
 sg13g2_buf_1 _0857_ (.A(_0215_),
    .X(_0273_));
 sg13g2_and4_1 _0858_ (.A(_0001_),
    .B(\cutoff2[1] ),
    .C(\cutoff2[3] ),
    .D(_0254_),
    .X(_0274_));
 sg13g2_nand3_1 _0859_ (.B(_0251_),
    .C(_0274_),
    .A(\cutoff2[0] ),
    .Y(_0275_));
 sg13g2_nor4_1 _0860_ (.A(_0239_),
    .B(net23),
    .C(net26),
    .D(_0275_),
    .Y(_0276_));
 sg13g2_xnor2_1 _0861_ (.Y(_0277_),
    .A(\cutoff2[4] ),
    .B(_0276_));
 sg13g2_nor2_1 _0862_ (.A(_0199_),
    .B(_0277_),
    .Y(_0118_));
 sg13g2_inv_1 _0863_ (.Y(_0278_),
    .A(vborder2));
 sg13g2_or4_1 _0864_ (.A(_0243_),
    .B(\vscheudler2.blockline[3] ),
    .C(\vscheudler2.blockline[2] ),
    .D(_0261_),
    .X(_0279_));
 sg13g2_inv_1 _0865_ (.Y(_0280_),
    .A(\vscheudler2.blockline[2] ));
 sg13g2_nand2_1 _0866_ (.Y(_0281_),
    .A(_0243_),
    .B(\vscheudler2.blockline[0] ));
 sg13g2_nor4_1 _0867_ (.A(\vscheudler2.blockline[3] ),
    .B(_0280_),
    .C(\vscheudler2.blockline[4] ),
    .D(_0281_),
    .Y(_0282_));
 sg13g2_nand2_1 _0868_ (.Y(_0283_),
    .A(_0148_),
    .B(_0184_));
 sg13g2_buf_1 _0869_ (.A(_0283_),
    .X(_0284_));
 sg13g2_nor2_1 _0870_ (.A(_0239_),
    .B(net22),
    .Y(_0285_));
 sg13g2_a221oi_1 _0871_ (.B2(_0285_),
    .C1(_0198_),
    .B1(_0282_),
    .A1(_0278_),
    .Y(_0119_),
    .A2(_0279_));
 sg13g2_inv_1 _0872_ (.Y(_0286_),
    .A(\vcount[3] ));
 sg13g2_inv_1 _0873_ (.Y(_0287_),
    .A(\vcount[7] ));
 sg13g2_nor4_1 _0874_ (.A(_0286_),
    .B(_0233_),
    .C(_0287_),
    .D(\vcount[6] ),
    .Y(_0288_));
 sg13g2_a21oi_1 _0875_ (.A1(_0232_),
    .A2(_0288_),
    .Y(_0289_),
    .B1(_0238_));
 sg13g2_nor2_1 _0876_ (.A(net33),
    .B(_0289_),
    .Y(_0120_));
 sg13g2_or2_1 _0877_ (.X(_0290_),
    .B(_0138_),
    .A(_0135_));
 sg13g2_nand2b_1 _0878_ (.Y(_0291_),
    .B(\cutoff2[0] ),
    .A_N(\l2[0] ));
 sg13g2_or2_1 _0879_ (.X(_0292_),
    .B(\l2[1] ),
    .A(\l2[2] ));
 sg13g2_a21oi_1 _0880_ (.A1(_0253_),
    .A2(_0291_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_nand2b_1 _0881_ (.Y(_0294_),
    .B(\cutoff2[3] ),
    .A_N(\l2[3] ));
 sg13g2_nand3b_1 _0882_ (.B(_0254_),
    .C(\cutoff2[1] ),
    .Y(_0295_),
    .A_N(\l2[1] ));
 sg13g2_nand2b_1 _0883_ (.Y(_0296_),
    .B(_0254_),
    .A_N(\l2[2] ));
 sg13g2_nand3_1 _0884_ (.B(_0295_),
    .C(_0296_),
    .A(_0294_),
    .Y(_0297_));
 sg13g2_nand2b_1 _0885_ (.Y(_0298_),
    .B(\l2[3] ),
    .A_N(\cutoff2[3] ));
 sg13g2_o21ai_1 _0886_ (.B1(_0298_),
    .Y(_0299_),
    .A1(_0293_),
    .A2(_0297_));
 sg13g2_nor2b_1 _0887_ (.A(_0254_),
    .B_N(\l2[2] ),
    .Y(_0300_));
 sg13g2_nand2b_1 _0888_ (.Y(_0301_),
    .B(_0254_),
    .A_N(\l2[1] ));
 sg13g2_o21ai_1 _0889_ (.B1(_0301_),
    .Y(_0302_),
    .A1(_0253_),
    .A2(_0300_));
 sg13g2_nor2b_1 _0890_ (.A(_0291_),
    .B_N(_0298_),
    .Y(_0303_));
 sg13g2_inv_1 _0891_ (.Y(_0304_),
    .A(_0002_));
 sg13g2_a21oi_2 _0892_ (.B1(_0304_),
    .Y(_0305_),
    .A2(_0303_),
    .A1(_0302_));
 sg13g2_nor2b_1 _0893_ (.A(vborder2),
    .B_N(\count2[1] ),
    .Y(_0306_));
 sg13g2_a21oi_1 _0894_ (.A1(_0299_),
    .A2(_0305_),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_inv_1 _0895_ (.Y(_0308_),
    .A(net1));
 sg13g2_nand2_1 _0896_ (.Y(_0309_),
    .A(\vga_sync.yvisible ),
    .B(\vga_sync.xvisible ));
 sg13g2_nor2_1 _0897_ (.A(_0308_),
    .B(_0309_),
    .Y(_0310_));
 sg13g2_o21ai_1 _0898_ (.B1(_0310_),
    .Y(_0311_),
    .A1(_0135_),
    .A2(_0139_));
 sg13g2_a21oi_1 _0899_ (.A1(_0290_),
    .A2(_0307_),
    .Y(_0011_),
    .B1(_0311_));
 sg13g2_nor2_1 _0900_ (.A(_0135_),
    .B(_0138_),
    .Y(_0312_));
 sg13g2_nand3_1 _0901_ (.B(_0299_),
    .C(_0305_),
    .A(_0310_),
    .Y(_0313_));
 sg13g2_o21ai_1 _0902_ (.B1(_0140_),
    .Y(_0012_),
    .A1(_0312_),
    .A2(_0313_));
 sg13g2_and2_1 _0903_ (.A(_0299_),
    .B(_0305_),
    .X(_0314_));
 sg13g2_a21oi_1 _0904_ (.A1(_0290_),
    .A2(_0314_),
    .Y(_0013_),
    .B1(_0124_));
 sg13g2_buf_1 _0905_ (.A(_0308_),
    .X(_0315_));
 sg13g2_nand2_1 _0906_ (.Y(_0316_),
    .A(\color_ditherer.dither ),
    .B(\bd[0] ));
 sg13g2_xor2_1 _0907_ (.B(_0316_),
    .A(\bd[1] ),
    .X(_0317_));
 sg13g2_nor2_1 _0908_ (.A(net39),
    .B(_0317_),
    .Y(_0014_));
 sg13g2_nand3_1 _0909_ (.B(\bd[0] ),
    .C(\bd[1] ),
    .A(\color_ditherer.dither ),
    .Y(_0318_));
 sg13g2_xor2_1 _0910_ (.B(_0318_),
    .A(\bd[2] ),
    .X(_0319_));
 sg13g2_nor2_1 _0911_ (.A(_0315_),
    .B(_0319_),
    .Y(_0015_));
 sg13g2_nand2_1 _0912_ (.Y(_0320_),
    .A(\color_ditherer.gin[0] ),
    .B(\color_ditherer.dither ));
 sg13g2_xor2_1 _0913_ (.B(_0320_),
    .A(\color_ditherer.gin[1] ),
    .X(_0321_));
 sg13g2_nor2_1 _0914_ (.A(_0315_),
    .B(_0321_),
    .Y(_0016_));
 sg13g2_nand3_1 _0915_ (.B(\color_ditherer.dither ),
    .C(\color_ditherer.gin[1] ),
    .A(\color_ditherer.gin[0] ),
    .Y(_0322_));
 sg13g2_xor2_1 _0916_ (.B(_0322_),
    .A(\color_ditherer.gin[2] ),
    .X(_0323_));
 sg13g2_nor2_1 _0917_ (.A(net39),
    .B(_0323_),
    .Y(_0017_));
 sg13g2_buf_1 _0918_ (.A(_0284_),
    .X(_0324_));
 sg13g2_nor2_1 _0919_ (.A(\count1b[0] ),
    .B(net11),
    .Y(_0325_));
 sg13g2_buf_1 _0920_ (.A(net25),
    .X(_0326_));
 sg13g2_buf_1 _0921_ (.A(net24),
    .X(_0327_));
 sg13g2_inv_1 _0922_ (.Y(_0328_),
    .A(\count1[0] ));
 sg13g2_nor2_1 _0923_ (.A(_0328_),
    .B(net35),
    .Y(_0329_));
 sg13g2_a221oi_1 _0924_ (.B2(net20),
    .C1(_0329_),
    .B1(_0326_),
    .A1(_0004_),
    .Y(_0330_),
    .A2(net35));
 sg13g2_buf_1 _0925_ (.A(_0121_),
    .X(_0331_));
 sg13g2_buf_1 _0926_ (.A(net38),
    .X(_0332_));
 sg13g2_o21ai_1 _0927_ (.B1(net32),
    .Y(_0018_),
    .A1(_0325_),
    .A2(_0330_));
 sg13g2_nor2_1 _0928_ (.A(\count1b[1] ),
    .B(net11),
    .Y(_0333_));
 sg13g2_a21o_1 _0929_ (.A2(net35),
    .A1(\count1[0] ),
    .B1(\count1[1] ),
    .X(_0334_));
 sg13g2_nand3_1 _0930_ (.B(\count1[1] ),
    .C(net35),
    .A(\count1[0] ),
    .Y(_0335_));
 sg13g2_a21oi_1 _0931_ (.A1(_0334_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(_0259_));
 sg13g2_o21ai_1 _0932_ (.B1(net32),
    .Y(_0019_),
    .A1(_0333_),
    .A2(_0336_));
 sg13g2_nor2_1 _0933_ (.A(\count1b[2] ),
    .B(net11),
    .Y(_0337_));
 sg13g2_buf_1 _0934_ (.A(_0259_),
    .X(_0338_));
 sg13g2_xnor2_1 _0935_ (.Y(_0339_),
    .A(\count1[2] ),
    .B(_0335_));
 sg13g2_nor2_1 _0936_ (.A(_0338_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_o21ai_1 _0937_ (.B1(_0332_),
    .Y(_0020_),
    .A1(_0337_),
    .A2(_0340_));
 sg13g2_buf_1 _0938_ (.A(net41),
    .X(_0341_));
 sg13g2_and3_1 _0939_ (.X(_0342_),
    .A(\vcount[7] ),
    .B(\vcount[6] ),
    .C(\vcount[8] ));
 sg13g2_nor2_1 _0940_ (.A(\vcount[4] ),
    .B(\vcount[9] ),
    .Y(_0343_));
 sg13g2_nand3_1 _0941_ (.B(_0342_),
    .C(_0343_),
    .A(\vcount[5] ),
    .Y(_0344_));
 sg13g2_nor2_1 _0942_ (.A(\vcount[3] ),
    .B(_0233_),
    .Y(_0345_));
 sg13g2_nor2b_1 _0943_ (.A(net40),
    .B_N(\vcount[1] ),
    .Y(_0346_));
 sg13g2_nand4_1 _0944_ (.B(_0182_),
    .C(_0345_),
    .A(_0181_),
    .Y(_0347_),
    .D(_0346_));
 sg13g2_nor3_2 _0945_ (.A(net27),
    .B(_0344_),
    .C(_0347_),
    .Y(_0348_));
 sg13g2_nand2b_1 _0946_ (.Y(_0349_),
    .B(\count1b[0] ),
    .A_N(_0348_));
 sg13g2_nand2_1 _0947_ (.Y(_0350_),
    .A(_0008_),
    .B(_0348_));
 sg13g2_nand3_1 _0948_ (.B(_0349_),
    .C(_0350_),
    .A(net37),
    .Y(_0021_));
 sg13g2_inv_1 _0949_ (.Y(_0351_),
    .A(\count1b[0] ));
 sg13g2_nor4_2 _0950_ (.A(_0351_),
    .B(net27),
    .C(_0344_),
    .Y(_0352_),
    .D(_0347_));
 sg13g2_xnor2_1 _0951_ (.Y(_0353_),
    .A(\count1b[1] ),
    .B(_0352_));
 sg13g2_nand2_1 _0952_ (.Y(_0022_),
    .A(net32),
    .B(_0353_));
 sg13g2_nand2_1 _0953_ (.Y(_0354_),
    .A(\count1b[2] ),
    .B(net38));
 sg13g2_nand2b_1 _0954_ (.Y(_0355_),
    .B(net38),
    .A_N(\count1b[2] ));
 sg13g2_nand2_1 _0955_ (.Y(_0356_),
    .A(\count1b[1] ),
    .B(_0352_));
 sg13g2_mux2_1 _0956_ (.A0(_0354_),
    .A1(_0355_),
    .S(_0356_),
    .X(_0023_));
 sg13g2_nor2_1 _0957_ (.A(\count2b[0] ),
    .B(_0324_),
    .Y(_0357_));
 sg13g2_and2_1 _0958_ (.A(\count2[0] ),
    .B(_0309_),
    .X(_0358_));
 sg13g2_a221oi_1 _0959_ (.B2(net20),
    .C1(_0358_),
    .B1(net21),
    .A1(_0003_),
    .Y(_0359_),
    .A2(net35));
 sg13g2_o21ai_1 _0960_ (.B1(net32),
    .Y(_0024_),
    .A1(_0357_),
    .A2(_0359_));
 sg13g2_nor2_1 _0961_ (.A(\count2b[1] ),
    .B(_0324_),
    .Y(_0360_));
 sg13g2_nand2_1 _0962_ (.Y(_0361_),
    .A(\count2[0] ),
    .B(_0123_));
 sg13g2_xnor2_1 _0963_ (.Y(_0362_),
    .A(\count2[1] ),
    .B(_0361_));
 sg13g2_nor2_1 _0964_ (.A(_0338_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_o21ai_1 _0965_ (.B1(net32),
    .Y(_0025_),
    .A1(_0360_),
    .A2(_0363_));
 sg13g2_nand4_1 _0966_ (.B(_0342_),
    .C(_0343_),
    .A(\vcount[5] ),
    .Y(_0364_),
    .D(_0345_));
 sg13g2_nand2_1 _0967_ (.Y(_0365_),
    .A(count2low),
    .B(_0346_));
 sg13g2_nor4_2 _0968_ (.A(net27),
    .B(_0215_),
    .C(_0364_),
    .Y(_0366_),
    .D(_0365_));
 sg13g2_buf_8 _0969_ (.A(_0366_),
    .X(_0367_));
 sg13g2_xnor2_1 _0970_ (.Y(_0368_),
    .A(\count2b[0] ),
    .B(net18));
 sg13g2_nand2_1 _0971_ (.Y(_0026_),
    .A(net32),
    .B(_0368_));
 sg13g2_a21oi_1 _0972_ (.A1(\count2b[0] ),
    .A2(_0366_),
    .Y(_0369_),
    .B1(\count2b[1] ));
 sg13g2_and3_1 _0973_ (.X(_0370_),
    .A(\count2b[1] ),
    .B(\count2b[0] ),
    .C(_0366_));
 sg13g2_o21ai_1 _0974_ (.B1(_0332_),
    .Y(_0027_),
    .A1(_0369_),
    .A2(_0370_));
 sg13g2_nand2b_1 _0975_ (.Y(_0371_),
    .B(count2low),
    .A_N(_0348_));
 sg13g2_nand2_1 _0976_ (.Y(_0372_),
    .A(_0009_),
    .B(_0348_));
 sg13g2_nand3_1 _0977_ (.B(_0371_),
    .C(_0372_),
    .A(net37),
    .Y(_0028_));
 sg13g2_nand3_1 _0978_ (.B(_0309_),
    .C(net22),
    .A(\color_ditherer.dither ),
    .Y(_0373_));
 sg13g2_o21ai_1 _0979_ (.B1(_0005_),
    .Y(_0374_),
    .A1(net35),
    .A2(_0259_));
 sg13g2_a21oi_1 _0980_ (.A1(_0373_),
    .A2(_0374_),
    .Y(_0029_),
    .B1(net39));
 sg13g2_nand2_1 _0981_ (.Y(_0375_),
    .A(\lfsr1b[0] ),
    .B(net19));
 sg13g2_xor2_1 _0982_ (.B(\lfsr1[9] ),
    .A(\lfsr1[6] ),
    .X(_0376_));
 sg13g2_nand3_1 _0983_ (.B(_0122_),
    .C(_0136_),
    .A(_0328_),
    .Y(_0377_));
 sg13g2_buf_1 _0984_ (.A(_0377_),
    .X(_0378_));
 sg13g2_mux2_1 _0985_ (.A0(_0376_),
    .A1(\l1[0] ),
    .S(net28),
    .X(_0379_));
 sg13g2_nand2_1 _0986_ (.Y(_0380_),
    .A(net11),
    .B(_0379_));
 sg13g2_nand3_1 _0987_ (.B(_0375_),
    .C(_0380_),
    .A(net37),
    .Y(_0030_));
 sg13g2_nand2_1 _0988_ (.Y(_0381_),
    .A(\lfsr1b[1] ),
    .B(net19));
 sg13g2_xor2_1 _0989_ (.B(\lfsr1[8] ),
    .A(\lfsr1[5] ),
    .X(_0382_));
 sg13g2_mux2_1 _0990_ (.A0(_0382_),
    .A1(\l1[1] ),
    .S(net28),
    .X(_0383_));
 sg13g2_nand2_1 _0991_ (.Y(_0384_),
    .A(net11),
    .B(_0383_));
 sg13g2_nand3_1 _0992_ (.B(_0381_),
    .C(_0384_),
    .A(net37),
    .Y(_0031_));
 sg13g2_nand2_1 _0993_ (.Y(_0385_),
    .A(\lfsr1b[2] ),
    .B(net19));
 sg13g2_xor2_1 _0994_ (.B(\lfsr1[7] ),
    .A(\lfsr1[4] ),
    .X(_0386_));
 sg13g2_mux2_1 _0995_ (.A0(_0386_),
    .A1(\l1[2] ),
    .S(net28),
    .X(_0387_));
 sg13g2_nand2_1 _0996_ (.Y(_0388_),
    .A(net11),
    .B(_0387_));
 sg13g2_nand3_1 _0997_ (.B(_0385_),
    .C(_0388_),
    .A(net37),
    .Y(_0032_));
 sg13g2_nor2_1 _0998_ (.A(\lfsr1b[3] ),
    .B(net11),
    .Y(_0389_));
 sg13g2_nand4_1 _0999_ (.B(\lfsr1[6] ),
    .C(net35),
    .A(_0328_),
    .Y(_0390_),
    .D(_0136_));
 sg13g2_xnor2_1 _1000_ (.Y(_0391_),
    .A(\l1[3] ),
    .B(_0390_));
 sg13g2_nor2_1 _1001_ (.A(net19),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_o21ai_1 _1002_ (.B1(net32),
    .Y(_0033_),
    .A1(_0389_),
    .A2(_0392_));
 sg13g2_nor2_1 _1003_ (.A(\lfsr1b[4] ),
    .B(net11),
    .Y(_0393_));
 sg13g2_mux2_1 _1004_ (.A0(\l1[0] ),
    .A1(\lfsr1[4] ),
    .S(net28),
    .X(_0394_));
 sg13g2_nor2_1 _1005_ (.A(net19),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_o21ai_1 _1006_ (.B1(net32),
    .Y(_0034_),
    .A1(_0393_),
    .A2(_0395_));
 sg13g2_nor2_1 _1007_ (.A(\lfsr1b[5] ),
    .B(net22),
    .Y(_0396_));
 sg13g2_mux2_1 _1008_ (.A0(\l1[1] ),
    .A1(\lfsr1[5] ),
    .S(net28),
    .X(_0397_));
 sg13g2_nor2_1 _1009_ (.A(net19),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_buf_1 _1010_ (.A(net38),
    .X(_0399_));
 sg13g2_o21ai_1 _1011_ (.B1(net31),
    .Y(_0035_),
    .A1(_0396_),
    .A2(_0398_));
 sg13g2_nor2_1 _1012_ (.A(\lfsr1b[6] ),
    .B(net22),
    .Y(_0400_));
 sg13g2_mux2_1 _1013_ (.A0(\l1[2] ),
    .A1(\lfsr1[6] ),
    .S(net28),
    .X(_0401_));
 sg13g2_nor2_1 _1014_ (.A(net19),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_o21ai_1 _1015_ (.B1(net31),
    .Y(_0036_),
    .A1(_0400_),
    .A2(_0402_));
 sg13g2_nor2_1 _1016_ (.A(\lfsr1b[7] ),
    .B(net22),
    .Y(_0403_));
 sg13g2_mux2_1 _1017_ (.A0(\l1[3] ),
    .A1(\lfsr1[7] ),
    .S(net28),
    .X(_0404_));
 sg13g2_nor2_1 _1018_ (.A(_0259_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_o21ai_1 _1019_ (.B1(net31),
    .Y(_0037_),
    .A1(_0403_),
    .A2(_0405_));
 sg13g2_nor2_1 _1020_ (.A(\lfsr1b[8] ),
    .B(net22),
    .Y(_0406_));
 sg13g2_mux2_1 _1021_ (.A0(\lfsr1[4] ),
    .A1(\lfsr1[8] ),
    .S(net28),
    .X(_0407_));
 sg13g2_nor2_1 _1022_ (.A(_0259_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_o21ai_1 _1023_ (.B1(net31),
    .Y(_0038_),
    .A1(_0406_),
    .A2(_0408_));
 sg13g2_nor2_1 _1024_ (.A(\lfsr1b[9] ),
    .B(net22),
    .Y(_0409_));
 sg13g2_mux2_1 _1025_ (.A0(\lfsr1[5] ),
    .A1(\lfsr1[9] ),
    .S(_0378_),
    .X(_0410_));
 sg13g2_nor2_1 _1026_ (.A(_0259_),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_o21ai_1 _1027_ (.B1(net31),
    .Y(_0039_),
    .A1(_0409_),
    .A2(_0411_));
 sg13g2_or3_1 _1028_ (.A(\count1b[1] ),
    .B(\count1b[0] ),
    .C(\count1b[2] ),
    .X(_0412_));
 sg13g2_nor4_1 _1029_ (.A(net27),
    .B(_0344_),
    .C(_0347_),
    .D(_0412_),
    .Y(_0413_));
 sg13g2_buf_1 _1030_ (.A(_0413_),
    .X(_0414_));
 sg13g2_nand2b_1 _1031_ (.Y(_0415_),
    .B(\lfsr1b[0] ),
    .A_N(net17));
 sg13g2_xor2_1 _1032_ (.B(\lfsr1b[9] ),
    .A(\lfsr1b[6] ),
    .X(_0416_));
 sg13g2_buf_1 _1033_ (.A(_0413_),
    .X(_0417_));
 sg13g2_nand2_1 _1034_ (.Y(_0418_),
    .A(_0416_),
    .B(net16));
 sg13g2_nand3_1 _1035_ (.B(_0415_),
    .C(_0418_),
    .A(net37),
    .Y(_0040_));
 sg13g2_xor2_1 _1036_ (.B(\lfsr1b[8] ),
    .A(\lfsr1b[5] ),
    .X(_0419_));
 sg13g2_nand2_1 _1037_ (.Y(_0420_),
    .A(net16),
    .B(_0419_));
 sg13g2_nand2b_1 _1038_ (.Y(_0421_),
    .B(\lfsr1b[1] ),
    .A_N(net17));
 sg13g2_nand3_1 _1039_ (.B(_0420_),
    .C(_0421_),
    .A(net37),
    .Y(_0041_));
 sg13g2_xor2_1 _1040_ (.B(\lfsr1b[7] ),
    .A(\lfsr1b[4] ),
    .X(_0422_));
 sg13g2_nand2_1 _1041_ (.Y(_0423_),
    .A(net16),
    .B(_0422_));
 sg13g2_nand2b_1 _1042_ (.Y(_0424_),
    .B(\lfsr1b[2] ),
    .A_N(net17));
 sg13g2_nand3_1 _1043_ (.B(_0423_),
    .C(_0424_),
    .A(net37),
    .Y(_0042_));
 sg13g2_nand2b_1 _1044_ (.Y(_0425_),
    .B(net41),
    .A_N(\lfsr1b[3] ));
 sg13g2_a21oi_1 _1045_ (.A1(\lfsr1b[6] ),
    .A2(_0417_),
    .Y(_0426_),
    .B1(_0425_));
 sg13g2_nand4_1 _1046_ (.B(\lfsr1b[6] ),
    .C(\lfsr1b[3] ),
    .A(net41),
    .Y(_0427_),
    .D(net17));
 sg13g2_nor2b_1 _1047_ (.A(_0426_),
    .B_N(_0427_),
    .Y(_0043_));
 sg13g2_buf_1 _1048_ (.A(net41),
    .X(_0428_));
 sg13g2_nand2b_1 _1049_ (.Y(_0429_),
    .B(\lfsr1b[4] ),
    .A_N(net17));
 sg13g2_nand2_1 _1050_ (.Y(_0430_),
    .A(\lfsr1b[0] ),
    .B(net16));
 sg13g2_nand3_1 _1051_ (.B(_0429_),
    .C(_0430_),
    .A(net36),
    .Y(_0044_));
 sg13g2_nand2b_1 _1052_ (.Y(_0431_),
    .B(\lfsr1b[5] ),
    .A_N(net17));
 sg13g2_nand2_1 _1053_ (.Y(_0432_),
    .A(\lfsr1b[1] ),
    .B(net16));
 sg13g2_nand3_1 _1054_ (.B(_0431_),
    .C(_0432_),
    .A(net36),
    .Y(_0045_));
 sg13g2_nand2b_1 _1055_ (.Y(_0433_),
    .B(\lfsr1b[6] ),
    .A_N(_0414_));
 sg13g2_nand2_1 _1056_ (.Y(_0434_),
    .A(\lfsr1b[2] ),
    .B(net16));
 sg13g2_nand3_1 _1057_ (.B(_0433_),
    .C(_0434_),
    .A(net36),
    .Y(_0046_));
 sg13g2_nand2b_1 _1058_ (.Y(_0435_),
    .B(\lfsr1b[7] ),
    .A_N(_0414_));
 sg13g2_nand2_1 _1059_ (.Y(_0436_),
    .A(\lfsr1b[3] ),
    .B(_0417_));
 sg13g2_nand3_1 _1060_ (.B(_0435_),
    .C(_0436_),
    .A(net36),
    .Y(_0047_));
 sg13g2_nand2b_1 _1061_ (.Y(_0437_),
    .B(\lfsr1b[8] ),
    .A_N(net17));
 sg13g2_nand2_1 _1062_ (.Y(_0438_),
    .A(\lfsr1b[4] ),
    .B(net16));
 sg13g2_nand3_1 _1063_ (.B(_0437_),
    .C(_0438_),
    .A(net36),
    .Y(_0048_));
 sg13g2_nand2b_1 _1064_ (.Y(_0439_),
    .B(\lfsr1b[9] ),
    .A_N(net17));
 sg13g2_nand2_1 _1065_ (.Y(_0440_),
    .A(\lfsr1b[5] ),
    .B(net16));
 sg13g2_nand3_1 _1066_ (.B(_0439_),
    .C(_0440_),
    .A(net36),
    .Y(_0049_));
 sg13g2_nor2_1 _1067_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .Y(_0441_));
 sg13g2_a22oi_1 _1068_ (.Y(_0442_),
    .B1(_0441_),
    .B2(_0123_),
    .A2(_0184_),
    .A1(_0148_));
 sg13g2_buf_1 _1069_ (.A(_0442_),
    .X(_0443_));
 sg13g2_nor3_1 _1070_ (.A(\lfsr2b[0] ),
    .B(net23),
    .C(net26),
    .Y(_0444_));
 sg13g2_xor2_1 _1071_ (.B(\lfsr2[9] ),
    .A(\lfsr2[6] ),
    .X(_0445_));
 sg13g2_a21oi_1 _1072_ (.A1(net21),
    .A2(net20),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_nor3_1 _1073_ (.A(net15),
    .B(_0444_),
    .C(_0446_),
    .Y(_0447_));
 sg13g2_nand2_1 _1074_ (.Y(_0448_),
    .A(\l2[0] ),
    .B(net15));
 sg13g2_nand3b_1 _1075_ (.B(net36),
    .C(_0448_),
    .Y(_0050_),
    .A_N(_0447_));
 sg13g2_nor3_1 _1076_ (.A(\lfsr2b[1] ),
    .B(_0272_),
    .C(_0273_),
    .Y(_0449_));
 sg13g2_xor2_1 _1077_ (.B(\lfsr2[5] ),
    .A(\lfsr2[8] ),
    .X(_0450_));
 sg13g2_a21oi_1 _1078_ (.A1(_0326_),
    .A2(net20),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_nor3_1 _1079_ (.A(_0442_),
    .B(_0449_),
    .C(_0451_),
    .Y(_0452_));
 sg13g2_nand2_1 _1080_ (.Y(_0453_),
    .A(\l2[1] ),
    .B(net15));
 sg13g2_nand3b_1 _1081_ (.B(net36),
    .C(_0453_),
    .Y(_0051_),
    .A_N(_0452_));
 sg13g2_nor3_1 _1082_ (.A(\lfsr2b[2] ),
    .B(_0272_),
    .C(_0273_),
    .Y(_0454_));
 sg13g2_xor2_1 _1083_ (.B(\lfsr2[4] ),
    .A(\lfsr2[7] ),
    .X(_0455_));
 sg13g2_a21oi_1 _1084_ (.A1(net21),
    .A2(_0327_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_nor3_1 _1085_ (.A(_0442_),
    .B(_0454_),
    .C(_0456_),
    .Y(_0457_));
 sg13g2_nand2_1 _1086_ (.Y(_0458_),
    .A(\l2[2] ),
    .B(net15));
 sg13g2_nand3b_1 _1087_ (.B(_0428_),
    .C(_0458_),
    .Y(_0052_),
    .A_N(_0457_));
 sg13g2_nor2_1 _1088_ (.A(\lfsr2b[3] ),
    .B(net22),
    .Y(_0459_));
 sg13g2_inv_1 _1089_ (.Y(_0460_),
    .A(\lfsr2[6] ));
 sg13g2_nor4_1 _1090_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .C(_0460_),
    .D(_0309_),
    .Y(_0461_));
 sg13g2_xor2_1 _1091_ (.B(_0461_),
    .A(\l2[3] ),
    .X(_0462_));
 sg13g2_nor2_1 _1092_ (.A(_0259_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _1093_ (.B1(net31),
    .Y(_0053_),
    .A1(_0459_),
    .A2(_0463_));
 sg13g2_nand2b_1 _1094_ (.Y(_0464_),
    .B(net15),
    .A_N(\lfsr2[4] ));
 sg13g2_nand2_1 _1095_ (.Y(_0465_),
    .A(_0122_),
    .B(_0441_));
 sg13g2_o21ai_1 _1096_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0214_),
    .A2(_0215_));
 sg13g2_buf_1 _1097_ (.A(_0466_),
    .X(_0467_));
 sg13g2_buf_1 _1098_ (.A(net25),
    .X(_0468_));
 sg13g2_nand3_1 _1099_ (.B(net14),
    .C(net20),
    .A(\lfsr2b[4] ),
    .Y(_0469_));
 sg13g2_o21ai_1 _1100_ (.B1(\l2[0] ),
    .Y(_0470_),
    .A1(net23),
    .A2(net26));
 sg13g2_nand3_1 _1101_ (.B(_0469_),
    .C(_0470_),
    .A(_0467_),
    .Y(_0471_));
 sg13g2_and3_1 _1102_ (.X(_0054_),
    .A(_0428_),
    .B(_0464_),
    .C(_0471_));
 sg13g2_nand2b_1 _1103_ (.Y(_0472_),
    .B(_0443_),
    .A_N(\lfsr2[5] ));
 sg13g2_nand3_1 _1104_ (.B(net14),
    .C(net20),
    .A(\lfsr2b[5] ),
    .Y(_0473_));
 sg13g2_o21ai_1 _1105_ (.B1(\l2[1] ),
    .Y(_0474_),
    .A1(net23),
    .A2(net26));
 sg13g2_nand3_1 _1106_ (.B(_0473_),
    .C(_0474_),
    .A(_0467_),
    .Y(_0475_));
 sg13g2_and3_1 _1107_ (.X(_0055_),
    .A(net38),
    .B(_0472_),
    .C(_0475_));
 sg13g2_nand2_1 _1108_ (.Y(_0476_),
    .A(_0460_),
    .B(net15));
 sg13g2_nand3_1 _1109_ (.B(net14),
    .C(_0327_),
    .A(\lfsr2b[6] ),
    .Y(_0477_));
 sg13g2_o21ai_1 _1110_ (.B1(\l2[2] ),
    .Y(_0478_),
    .A1(net23),
    .A2(net26));
 sg13g2_nand3_1 _1111_ (.B(_0477_),
    .C(_0478_),
    .A(_0467_),
    .Y(_0479_));
 sg13g2_and3_1 _1112_ (.X(_0056_),
    .A(net38),
    .B(_0476_),
    .C(_0479_));
 sg13g2_nand2b_1 _1113_ (.Y(_0480_),
    .B(_0443_),
    .A_N(\lfsr2[7] ));
 sg13g2_nand3_1 _1114_ (.B(net14),
    .C(net20),
    .A(\lfsr2b[7] ),
    .Y(_0481_));
 sg13g2_o21ai_1 _1115_ (.B1(\l2[3] ),
    .Y(_0482_),
    .A1(net23),
    .A2(net26));
 sg13g2_nand3_1 _1116_ (.B(_0481_),
    .C(_0482_),
    .A(_0467_),
    .Y(_0483_));
 sg13g2_and3_1 _1117_ (.X(_0057_),
    .A(_0331_),
    .B(_0480_),
    .C(_0483_));
 sg13g2_nand2b_1 _1118_ (.Y(_0484_),
    .B(net15),
    .A_N(\lfsr2[8] ));
 sg13g2_o21ai_1 _1119_ (.B1(\lfsr2[4] ),
    .Y(_0485_),
    .A1(net23),
    .A2(net26));
 sg13g2_nand3_1 _1120_ (.B(_0468_),
    .C(_0185_),
    .A(\lfsr2b[8] ),
    .Y(_0486_));
 sg13g2_nand3_1 _1121_ (.B(_0485_),
    .C(_0486_),
    .A(_0467_),
    .Y(_0487_));
 sg13g2_a21o_1 _1122_ (.A2(_0487_),
    .A1(_0484_),
    .B1(_0308_),
    .X(_0058_));
 sg13g2_nand2b_1 _1123_ (.Y(_0488_),
    .B(net15),
    .A_N(\lfsr2[9] ));
 sg13g2_nand3_1 _1124_ (.B(_0468_),
    .C(net20),
    .A(\lfsr2b[9] ),
    .Y(_0489_));
 sg13g2_o21ai_1 _1125_ (.B1(\lfsr2[5] ),
    .Y(_0490_),
    .A1(net23),
    .A2(net26));
 sg13g2_nand3_1 _1126_ (.B(_0489_),
    .C(_0490_),
    .A(_0467_),
    .Y(_0491_));
 sg13g2_and3_1 _1127_ (.X(_0059_),
    .A(_0331_),
    .B(_0488_),
    .C(_0491_));
 sg13g2_nor2_1 _1128_ (.A(\count2b[1] ),
    .B(\count2b[0] ),
    .Y(_0492_));
 sg13g2_buf_1 _1129_ (.A(_0492_),
    .X(_0493_));
 sg13g2_a21oi_1 _1130_ (.A1(net18),
    .A2(net30),
    .Y(_0494_),
    .B1(\lfsr2b[0] ));
 sg13g2_or4_1 _1131_ (.A(net27),
    .B(_0215_),
    .C(_0364_),
    .D(_0365_),
    .X(_0495_));
 sg13g2_buf_1 _1132_ (.A(_0495_),
    .X(_0496_));
 sg13g2_or2_1 _1133_ (.X(_0497_),
    .B(\count2b[0] ),
    .A(\count2b[1] ));
 sg13g2_buf_1 _1134_ (.A(_0497_),
    .X(_0498_));
 sg13g2_xor2_1 _1135_ (.B(\lfsr2b[9] ),
    .A(\lfsr2b[6] ),
    .X(_0499_));
 sg13g2_nor3_1 _1136_ (.A(net13),
    .B(net29),
    .C(_0499_),
    .Y(_0500_));
 sg13g2_o21ai_1 _1137_ (.B1(net31),
    .Y(_0060_),
    .A1(_0494_),
    .A2(_0500_));
 sg13g2_a21oi_1 _1138_ (.A1(net18),
    .A2(net30),
    .Y(_0501_),
    .B1(\lfsr2b[1] ));
 sg13g2_xor2_1 _1139_ (.B(\lfsr2b[8] ),
    .A(\lfsr2b[5] ),
    .X(_0502_));
 sg13g2_nor3_1 _1140_ (.A(net13),
    .B(net29),
    .C(_0502_),
    .Y(_0503_));
 sg13g2_o21ai_1 _1141_ (.B1(net31),
    .Y(_0061_),
    .A1(_0501_),
    .A2(_0503_));
 sg13g2_a21oi_1 _1142_ (.A1(net18),
    .A2(_0493_),
    .Y(_0504_),
    .B1(\lfsr2b[2] ));
 sg13g2_xor2_1 _1143_ (.B(\lfsr2b[7] ),
    .A(\lfsr2b[4] ),
    .X(_0505_));
 sg13g2_nor3_1 _1144_ (.A(_0496_),
    .B(_0498_),
    .C(_0505_),
    .Y(_0506_));
 sg13g2_o21ai_1 _1145_ (.B1(_0399_),
    .Y(_0062_),
    .A1(_0504_),
    .A2(_0506_));
 sg13g2_nand2_1 _1146_ (.Y(_0507_),
    .A(net38),
    .B(\lfsr2b[3] ));
 sg13g2_nand2b_1 _1147_ (.Y(_0508_),
    .B(net38),
    .A_N(\lfsr2b[3] ));
 sg13g2_nand3_1 _1148_ (.B(_0366_),
    .C(net30),
    .A(\lfsr2b[6] ),
    .Y(_0509_));
 sg13g2_mux2_1 _1149_ (.A0(_0507_),
    .A1(_0508_),
    .S(_0509_),
    .X(_0063_));
 sg13g2_o21ai_1 _1150_ (.B1(\lfsr2b[4] ),
    .Y(_0510_),
    .A1(net13),
    .A2(net29));
 sg13g2_nand3_1 _1151_ (.B(_0367_),
    .C(net30),
    .A(\lfsr2b[0] ),
    .Y(_0511_));
 sg13g2_a21oi_1 _1152_ (.A1(_0510_),
    .A2(_0511_),
    .Y(_0064_),
    .B1(net39));
 sg13g2_o21ai_1 _1153_ (.B1(\lfsr2b[5] ),
    .Y(_0512_),
    .A1(net13),
    .A2(net29));
 sg13g2_nand3_1 _1154_ (.B(net18),
    .C(net30),
    .A(\lfsr2b[1] ),
    .Y(_0513_));
 sg13g2_a21oi_1 _1155_ (.A1(_0512_),
    .A2(_0513_),
    .Y(_0065_),
    .B1(net39));
 sg13g2_o21ai_1 _1156_ (.B1(\lfsr2b[6] ),
    .Y(_0514_),
    .A1(net13),
    .A2(net29));
 sg13g2_nand3_1 _1157_ (.B(_0367_),
    .C(net30),
    .A(\lfsr2b[2] ),
    .Y(_0515_));
 sg13g2_a21oi_1 _1158_ (.A1(_0514_),
    .A2(_0515_),
    .Y(_0066_),
    .B1(net39));
 sg13g2_o21ai_1 _1159_ (.B1(\lfsr2b[7] ),
    .Y(_0516_),
    .A1(net13),
    .A2(net29));
 sg13g2_nand3_1 _1160_ (.B(net18),
    .C(net30),
    .A(\lfsr2b[3] ),
    .Y(_0517_));
 sg13g2_a21oi_1 _1161_ (.A1(_0516_),
    .A2(_0517_),
    .Y(_0067_),
    .B1(net39));
 sg13g2_nor3_1 _1162_ (.A(\lfsr2b[4] ),
    .B(net13),
    .C(net29),
    .Y(_0518_));
 sg13g2_a21oi_1 _1163_ (.A1(net18),
    .A2(_0493_),
    .Y(_0519_),
    .B1(\lfsr2b[8] ));
 sg13g2_o21ai_1 _1164_ (.B1(_0399_),
    .Y(_0068_),
    .A1(_0518_),
    .A2(_0519_));
 sg13g2_o21ai_1 _1165_ (.B1(\lfsr2b[9] ),
    .Y(_0520_),
    .A1(net13),
    .A2(net29));
 sg13g2_nand3_1 _1166_ (.B(net18),
    .C(net30),
    .A(\lfsr2b[5] ),
    .Y(_0521_));
 sg13g2_a21oi_1 _1167_ (.A1(_0520_),
    .A2(_0521_),
    .Y(_0069_),
    .B1(net39));
 sg13g2_nand2_1 _1168_ (.Y(_0522_),
    .A(\count2[1] ),
    .B(_0278_));
 sg13g2_a21oi_1 _1169_ (.A1(_0299_),
    .A2(_0305_),
    .Y(_0523_),
    .B1(_0522_));
 sg13g2_a21oi_1 _1170_ (.A1(_0290_),
    .A2(_0523_),
    .Y(_0071_),
    .B1(_0124_));
 sg13g2_nand2_1 _1171_ (.Y(_0524_),
    .A(_0310_),
    .B(_0306_));
 sg13g2_a21oi_1 _1172_ (.A1(_0299_),
    .A2(_0305_),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_and2_1 _1173_ (.A(_0310_),
    .B(_0137_),
    .X(_0526_));
 sg13g2_mux2_1 _1174_ (.A0(_0525_),
    .A1(_0526_),
    .S(_0312_),
    .X(_0072_));
 sg13g2_nor4_1 _1175_ (.A(_0143_),
    .B(\hcount[3] ),
    .C(\hcount[2] ),
    .D(\hcount[8] ),
    .Y(_0527_));
 sg13g2_nand2_1 _1176_ (.Y(_0528_),
    .A(_0141_),
    .B(_0149_));
 sg13g2_nor4_1 _1177_ (.A(_0145_),
    .B(_0174_),
    .C(_0166_),
    .D(_0528_),
    .Y(_0529_));
 sg13g2_a21oi_1 _1178_ (.A1(_0527_),
    .A2(_0529_),
    .Y(_0530_),
    .B1(hsync));
 sg13g2_o21ai_1 _1179_ (.B1(_0341_),
    .Y(_0073_),
    .A1(net19),
    .A2(_0530_));
 sg13g2_or4_1 _1180_ (.A(net40),
    .B(_0286_),
    .C(_0233_),
    .D(_0344_),
    .X(_0531_));
 sg13g2_inv_1 _1181_ (.Y(_0532_),
    .A(\vcount[1] ));
 sg13g2_a21oi_1 _1182_ (.A1(\vga_sync.vga_vsync ),
    .A2(_0531_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nor3_1 _1183_ (.A(net40),
    .B(_0286_),
    .C(_0344_),
    .Y(_0534_));
 sg13g2_a21oi_1 _1184_ (.A1(_0233_),
    .A2(_0534_),
    .Y(_0535_),
    .B1(\vga_sync.vga_vsync ));
 sg13g2_o21ai_1 _1185_ (.B1(_0341_),
    .Y(_0074_),
    .A1(_0533_),
    .A2(_0535_));
 sg13g2_nor4_1 _1186_ (.A(\vcount[4] ),
    .B(\vcount[5] ),
    .C(\vcount[7] ),
    .D(\vcount[6] ),
    .Y(_0536_));
 sg13g2_nor4_1 _1187_ (.A(\vcount[1] ),
    .B(_0286_),
    .C(_0234_),
    .D(\vcount[8] ),
    .Y(_0537_));
 sg13g2_nand4_1 _1188_ (.B(\vcount[9] ),
    .C(_0536_),
    .A(_0227_),
    .Y(_0538_),
    .D(_0537_));
 sg13g2_o21ai_1 _1189_ (.B1(net41),
    .Y(_0539_),
    .A1(_0153_),
    .A2(_0538_));
 sg13g2_buf_1 _1190_ (.A(_0539_),
    .X(_0540_));
 sg13g2_xnor2_1 _1191_ (.Y(_0541_),
    .A(_0228_),
    .B(_0153_));
 sg13g2_nand2b_1 _1192_ (.Y(_0085_),
    .B(_0541_),
    .A_N(net10));
 sg13g2_o21ai_1 _1193_ (.B1(\vcount[1] ),
    .Y(_0542_),
    .A1(_0228_),
    .A2(_0153_));
 sg13g2_nand4_1 _1194_ (.B(_0532_),
    .C(net21),
    .A(net40),
    .Y(_0543_),
    .D(_0152_));
 sg13g2_a21oi_1 _1195_ (.A1(_0542_),
    .A2(_0543_),
    .Y(_0086_),
    .B1(_0540_));
 sg13g2_nor2_1 _1196_ (.A(_0228_),
    .B(_0532_),
    .Y(_0544_));
 sg13g2_nand3_1 _1197_ (.B(_0152_),
    .C(_0544_),
    .A(net21),
    .Y(_0545_));
 sg13g2_xnor2_1 _1198_ (.Y(_0546_),
    .A(_0234_),
    .B(_0545_));
 sg13g2_nor2_1 _1199_ (.A(net10),
    .B(_0546_),
    .Y(_0087_));
 sg13g2_nand4_1 _1200_ (.B(net14),
    .C(_0152_),
    .A(_0233_),
    .Y(_0547_),
    .D(_0544_));
 sg13g2_xnor2_1 _1201_ (.Y(_0548_),
    .A(_0286_),
    .B(_0547_));
 sg13g2_nor2_1 _1202_ (.A(net10),
    .B(_0548_),
    .Y(_0088_));
 sg13g2_nand4_1 _1203_ (.B(\vcount[1] ),
    .C(\vcount[3] ),
    .A(net40),
    .Y(_0549_),
    .D(_0233_));
 sg13g2_nor4_2 _1204_ (.A(_0149_),
    .B(_0150_),
    .C(_0151_),
    .Y(_0550_),
    .D(_0549_));
 sg13g2_nand2_1 _1205_ (.Y(_0551_),
    .A(net21),
    .B(_0550_));
 sg13g2_xor2_1 _1206_ (.B(_0551_),
    .A(\vcount[4] ),
    .X(_0552_));
 sg13g2_nor2_1 _1207_ (.A(net10),
    .B(_0552_),
    .Y(_0089_));
 sg13g2_nand3_1 _1208_ (.B(net21),
    .C(_0550_),
    .A(\vcount[4] ),
    .Y(_0553_));
 sg13g2_xor2_1 _1209_ (.B(_0553_),
    .A(\vcount[5] ),
    .X(_0554_));
 sg13g2_nor2_1 _1210_ (.A(net10),
    .B(_0554_),
    .Y(_0090_));
 sg13g2_nand3_1 _1211_ (.B(_0231_),
    .C(_0550_),
    .A(net21),
    .Y(_0555_));
 sg13g2_xnor2_1 _1212_ (.Y(_0556_),
    .A(_0235_),
    .B(_0555_));
 sg13g2_nor2_1 _1213_ (.A(net10),
    .B(_0556_),
    .Y(_0091_));
 sg13g2_nand4_1 _1214_ (.B(net14),
    .C(_0231_),
    .A(\vcount[6] ),
    .Y(_0557_),
    .D(_0550_));
 sg13g2_xnor2_1 _1215_ (.Y(_0558_),
    .A(_0287_),
    .B(_0557_));
 sg13g2_nor2_1 _1216_ (.A(_0540_),
    .B(_0558_),
    .Y(_0092_));
 sg13g2_nor2_1 _1217_ (.A(_0287_),
    .B(_0235_),
    .Y(_0559_));
 sg13g2_nand4_1 _1218_ (.B(_0231_),
    .C(_0559_),
    .A(net14),
    .Y(_0560_),
    .D(_0550_));
 sg13g2_xor2_1 _1219_ (.B(_0560_),
    .A(\vcount[8] ),
    .X(_0561_));
 sg13g2_nor2_1 _1220_ (.A(net10),
    .B(_0561_),
    .Y(_0093_));
 sg13g2_nand4_1 _1221_ (.B(_0231_),
    .C(_0342_),
    .A(net14),
    .Y(_0562_),
    .D(_0550_));
 sg13g2_xor2_1 _1222_ (.B(_0562_),
    .A(\vcount[9] ),
    .X(_0563_));
 sg13g2_nor2_1 _1223_ (.A(net10),
    .B(_0563_),
    .Y(_0094_));
 sg13g2_nor2_1 _1224_ (.A(\hcount[5] ),
    .B(\hcount[4] ),
    .Y(_0564_));
 sg13g2_nand4_1 _1225_ (.B(_0142_),
    .C(_0527_),
    .A(_0145_),
    .Y(_0565_),
    .D(_0564_));
 sg13g2_nor2_1 _1226_ (.A(\hcount[9] ),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_o21ai_1 _1227_ (.B1(_0169_),
    .Y(_0567_),
    .A1(\vga_sync.xvisible ),
    .A2(_0566_));
 sg13g2_o21ai_1 _1228_ (.B1(\vga_sync.xvisible ),
    .Y(_0568_),
    .A1(_0174_),
    .A2(_0565_));
 sg13g2_a21oi_1 _1229_ (.A1(_0567_),
    .A2(_0568_),
    .Y(_0095_),
    .B1(_0308_));
 sg13g2_nand2_1 _1230_ (.Y(_0569_),
    .A(net40),
    .B(_0532_));
 sg13g2_o21ai_1 _1231_ (.B1(\vga_sync.yvisible ),
    .Y(_0570_),
    .A1(_0364_),
    .A2(_0569_));
 sg13g2_nand4_1 _1232_ (.B(_0229_),
    .C(_0345_),
    .A(net40),
    .Y(_0571_),
    .D(_0536_));
 sg13g2_a21oi_1 _1233_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0096_),
    .B1(_0308_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \bd[0]$_SDFF_PN0__58  (.L_HI(net58));
 sg13g2_buf_1 _1236_ (.A(net42),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1237_ (.A(net43),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1238_ (.A(net44),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1239_ (.A(net45),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1240_ (.A(net46),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1241_ (.A(net47),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1242_ (.A(net48),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1243_ (.A(net49),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1244_ (.A(net50),
    .X(uio_out[0]));
 sg13g2_buf_1 _1245_ (.A(net51),
    .X(uio_out[1]));
 sg13g2_buf_1 _1246_ (.A(net52),
    .X(uio_out[2]));
 sg13g2_buf_1 _1247_ (.A(net53),
    .X(uio_out[3]));
 sg13g2_buf_1 _1248_ (.A(net54),
    .X(uio_out[4]));
 sg13g2_buf_1 _1249_ (.A(net55),
    .X(uio_out[5]));
 sg13g2_buf_1 _1250_ (.A(net56),
    .X(uio_out[6]));
 sg13g2_buf_1 _1251_ (.A(net57),
    .X(uio_out[7]));
 sg13g2_buf_1 _1252_ (.A(net3),
    .X(net2));
 sg13g2_buf_1 _1253_ (.A(\vga_sync.vga_vsync ),
    .X(net5));
 sg13g2_buf_1 _1254_ (.A(net7),
    .X(net6));
 sg13g2_buf_1 _1255_ (.A(hsync),
    .X(net9));
 sg13g2_dfrbp_1 \bd[0]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net58),
    .D(_0011_),
    .Q_N(_0670_),
    .Q(\bd[0] ));
 sg13g2_dfrbp_1 \bd[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net59),
    .D(_0012_),
    .Q_N(_0669_),
    .Q(\bd[1] ));
 sg13g2_dfrbp_1 \bd[2]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net60),
    .D(_0013_),
    .Q_N(_0668_),
    .Q(\bd[2] ));
 sg13g2_dfrbp_1 \color_ditherer.bout[0]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net61),
    .D(_0014_),
    .Q_N(_0667_),
    .Q(net8));
 sg13g2_dfrbp_1 \color_ditherer.bout[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net62),
    .D(_0015_),
    .Q_N(_0666_),
    .Q(net4));
 sg13g2_dfrbp_1 \color_ditherer.gout[0]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net63),
    .D(_0016_),
    .Q_N(_0665_),
    .Q(net7));
 sg13g2_dfrbp_1 \color_ditherer.gout[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net64),
    .D(_0017_),
    .Q_N(_0664_),
    .Q(net3));
 sg13g2_dfrbp_1 \count1[0]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net65),
    .D(_0018_),
    .Q_N(_0004_),
    .Q(\count1[0] ));
 sg13g2_dfrbp_1 \count1[1]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(_0019_),
    .Q_N(_0663_),
    .Q(\count1[1] ));
 sg13g2_dfrbp_1 \count1[2]$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net67),
    .D(_0020_),
    .Q_N(_0662_),
    .Q(\count1[2] ));
 sg13g2_dfrbp_1 \count1b[0]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net68),
    .D(_0021_),
    .Q_N(_0008_),
    .Q(\count1b[0] ));
 sg13g2_dfrbp_1 \count1b[1]$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net69),
    .D(_0022_),
    .Q_N(_0661_),
    .Q(\count1b[1] ));
 sg13g2_dfrbp_1 \count1b[2]$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net70),
    .D(_0023_),
    .Q_N(_0660_),
    .Q(\count1b[2] ));
 sg13g2_dfrbp_1 \count2[0]$_SDFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net71),
    .D(_0024_),
    .Q_N(_0003_),
    .Q(\count2[0] ));
 sg13g2_dfrbp_1 \count2[1]$_SDFFE_PN1P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net72),
    .D(_0025_),
    .Q_N(_0659_),
    .Q(\count2[1] ));
 sg13g2_dfrbp_1 \count2b[0]$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net73),
    .D(_0026_),
    .Q_N(_0658_),
    .Q(\count2b[0] ));
 sg13g2_dfrbp_1 \count2b[1]$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net74),
    .D(_0027_),
    .Q_N(_0657_),
    .Q(\count2b[1] ));
 sg13g2_dfrbp_1 \count2low$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net75),
    .D(_0028_),
    .Q_N(_0009_),
    .Q(count2low));
 sg13g2_dfrbp_1 \dither$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net76),
    .D(_0029_),
    .Q_N(_0005_),
    .Q(\color_ditherer.dither ));
 sg13g2_dfrbp_1 \lfsr1[0]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net77),
    .D(_0030_),
    .Q_N(_0656_),
    .Q(\l1[0] ));
 sg13g2_dfrbp_1 \lfsr1[1]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net78),
    .D(_0031_),
    .Q_N(_0655_),
    .Q(\l1[1] ));
 sg13g2_dfrbp_1 \lfsr1[2]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net79),
    .D(_0032_),
    .Q_N(_0654_),
    .Q(\l1[2] ));
 sg13g2_dfrbp_1 \lfsr1[3]$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net80),
    .D(_0033_),
    .Q_N(_0653_),
    .Q(\l1[3] ));
 sg13g2_dfrbp_1 \lfsr1[4]$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net81),
    .D(_0034_),
    .Q_N(_0652_),
    .Q(\lfsr1[4] ));
 sg13g2_dfrbp_1 \lfsr1[5]$_SDFFE_PN1P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net82),
    .D(_0035_),
    .Q_N(_0651_),
    .Q(\lfsr1[5] ));
 sg13g2_dfrbp_1 \lfsr1[6]$_SDFFE_PN1P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net83),
    .D(_0036_),
    .Q_N(_0650_),
    .Q(\lfsr1[6] ));
 sg13g2_dfrbp_1 \lfsr1[7]$_SDFFE_PN1P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net84),
    .D(_0037_),
    .Q_N(_0649_),
    .Q(\lfsr1[7] ));
 sg13g2_dfrbp_1 \lfsr1[8]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net85),
    .D(_0038_),
    .Q_N(_0648_),
    .Q(\lfsr1[8] ));
 sg13g2_dfrbp_1 \lfsr1[9]$_SDFFE_PN1P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net86),
    .D(_0039_),
    .Q_N(_0647_),
    .Q(\lfsr1[9] ));
 sg13g2_dfrbp_1 \lfsr1b[0]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net87),
    .D(_0040_),
    .Q_N(_0646_),
    .Q(\lfsr1b[0] ));
 sg13g2_dfrbp_1 \lfsr1b[1]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net88),
    .D(_0041_),
    .Q_N(_0645_),
    .Q(\lfsr1b[1] ));
 sg13g2_dfrbp_1 \lfsr1b[2]$_SDFFE_PN1P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net89),
    .D(_0042_),
    .Q_N(_0644_),
    .Q(\lfsr1b[2] ));
 sg13g2_dfrbp_1 \lfsr1b[3]$_SDFFE_PN1P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net90),
    .D(_0043_),
    .Q_N(_0643_),
    .Q(\lfsr1b[3] ));
 sg13g2_dfrbp_1 \lfsr1b[4]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net91),
    .D(_0044_),
    .Q_N(_0642_),
    .Q(\lfsr1b[4] ));
 sg13g2_dfrbp_1 \lfsr1b[5]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(_0045_),
    .Q_N(_0641_),
    .Q(\lfsr1b[5] ));
 sg13g2_dfrbp_1 \lfsr1b[6]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net93),
    .D(_0046_),
    .Q_N(_0640_),
    .Q(\lfsr1b[6] ));
 sg13g2_dfrbp_1 \lfsr1b[7]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net94),
    .D(_0047_),
    .Q_N(_0639_),
    .Q(\lfsr1b[7] ));
 sg13g2_dfrbp_1 \lfsr1b[8]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net95),
    .D(_0048_),
    .Q_N(_0638_),
    .Q(\lfsr1b[8] ));
 sg13g2_dfrbp_1 \lfsr1b[9]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net96),
    .D(_0049_),
    .Q_N(_0637_),
    .Q(\lfsr1b[9] ));
 sg13g2_dfrbp_1 \lfsr2[0]$_SDFFE_PN1P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net97),
    .D(_0050_),
    .Q_N(_0636_),
    .Q(\l2[0] ));
 sg13g2_dfrbp_1 \lfsr2[1]$_SDFFE_PN1P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net98),
    .D(_0051_),
    .Q_N(_0635_),
    .Q(\l2[1] ));
 sg13g2_dfrbp_1 \lfsr2[2]$_SDFFE_PN1P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net99),
    .D(_0052_),
    .Q_N(_0634_),
    .Q(\l2[2] ));
 sg13g2_dfrbp_1 \lfsr2[3]$_SDFFE_PN1P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net100),
    .D(_0053_),
    .Q_N(_0633_),
    .Q(\l2[3] ));
 sg13g2_dfrbp_1 \lfsr2[4]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net101),
    .D(_0054_),
    .Q_N(_0632_),
    .Q(\lfsr2[4] ));
 sg13g2_dfrbp_1 \lfsr2[5]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net102),
    .D(_0055_),
    .Q_N(_0631_),
    .Q(\lfsr2[5] ));
 sg13g2_dfrbp_1 \lfsr2[6]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net103),
    .D(_0056_),
    .Q_N(_0630_),
    .Q(\lfsr2[6] ));
 sg13g2_dfrbp_1 \lfsr2[7]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net104),
    .D(_0057_),
    .Q_N(_0629_),
    .Q(\lfsr2[7] ));
 sg13g2_dfrbp_1 \lfsr2[8]$_SDFFE_PN1P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net105),
    .D(_0058_),
    .Q_N(_0628_),
    .Q(\lfsr2[8] ));
 sg13g2_dfrbp_1 \lfsr2[9]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net106),
    .D(_0059_),
    .Q_N(_0627_),
    .Q(\lfsr2[9] ));
 sg13g2_dfrbp_1 \lfsr2b[0]$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net107),
    .D(_0060_),
    .Q_N(_0626_),
    .Q(\lfsr2b[0] ));
 sg13g2_dfrbp_1 \lfsr2b[1]$_SDFFE_PN1P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net108),
    .D(_0061_),
    .Q_N(_0625_),
    .Q(\lfsr2b[1] ));
 sg13g2_dfrbp_1 \lfsr2b[2]$_SDFFE_PN1P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net109),
    .D(_0062_),
    .Q_N(_0624_),
    .Q(\lfsr2b[2] ));
 sg13g2_dfrbp_1 \lfsr2b[3]$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net110),
    .D(_0063_),
    .Q_N(_0623_),
    .Q(\lfsr2b[3] ));
 sg13g2_dfrbp_1 \lfsr2b[4]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net111),
    .D(_0064_),
    .Q_N(_0622_),
    .Q(\lfsr2b[4] ));
 sg13g2_dfrbp_1 \lfsr2b[5]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net112),
    .D(_0065_),
    .Q_N(_0621_),
    .Q(\lfsr2b[5] ));
 sg13g2_dfrbp_1 \lfsr2b[6]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net113),
    .D(_0066_),
    .Q_N(_0620_),
    .Q(\lfsr2b[6] ));
 sg13g2_dfrbp_1 \lfsr2b[7]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net114),
    .D(_0067_),
    .Q_N(_0619_),
    .Q(\lfsr2b[7] ));
 sg13g2_dfrbp_1 \lfsr2b[8]$_SDFFE_PN1P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net115),
    .D(_0068_),
    .Q_N(_0618_),
    .Q(\lfsr2b[8] ));
 sg13g2_dfrbp_1 \lfsr2b[9]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net116),
    .D(_0069_),
    .Q_N(_0617_),
    .Q(\lfsr2b[9] ));
 sg13g2_dfrbp_1 \rd[0]$_SDFF_PP0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net117),
    .D(_0070_),
    .Q_N(_0616_),
    .Q(\color_ditherer.gin[0] ));
 sg13g2_dfrbp_1 \rd[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net118),
    .D(_0071_),
    .Q_N(_0615_),
    .Q(\color_ditherer.gin[1] ));
 sg13g2_dfrbp_1 \rd[2]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net119),
    .D(_0072_),
    .Q_N(_0614_),
    .Q(\color_ditherer.gin[2] ));
 sg13g2_dfrbp_1 \vga_sync.vga_hsync$_SDFFE_PN1P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net120),
    .D(_0073_),
    .Q_N(_0613_),
    .Q(hsync));
 sg13g2_dfrbp_1 \vga_sync.vga_vsync$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net121),
    .D(_0074_),
    .Q_N(_0612_),
    .Q(\vga_sync.vga_vsync ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[0]$_SDFF_PP1_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net122),
    .D(_0075_),
    .Q_N(_0010_),
    .Q(\hcount[0] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[1]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net123),
    .D(_0076_),
    .Q_N(_0611_),
    .Q(\hcount[1] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[2]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net124),
    .D(_0077_),
    .Q_N(_0610_),
    .Q(\hcount[2] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[3]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net125),
    .D(_0078_),
    .Q_N(_0609_),
    .Q(\hcount[3] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[4]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net126),
    .D(_0079_),
    .Q_N(_0608_),
    .Q(\hcount[4] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[5]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net127),
    .D(_0080_),
    .Q_N(_0607_),
    .Q(\hcount[5] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[6]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net128),
    .D(_0081_),
    .Q_N(_0606_),
    .Q(\hcount[6] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[7]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net129),
    .D(_0082_),
    .Q_N(_0605_),
    .Q(\hcount[7] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[8]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net130),
    .D(_0083_),
    .Q_N(_0604_),
    .Q(\hcount[8] ));
 sg13g2_dfrbp_1 \vga_sync.vga_xpos[9]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net131),
    .D(_0084_),
    .Q_N(_0603_),
    .Q(\hcount[9] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[0]$_SDFFE_PN1N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net132),
    .D(_0085_),
    .Q_N(_0602_),
    .Q(\vcount[0] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[1]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net133),
    .D(_0086_),
    .Q_N(_0601_),
    .Q(\vcount[1] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[2]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net134),
    .D(_0087_),
    .Q_N(_0600_),
    .Q(\vcount[2] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[3]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net135),
    .D(_0088_),
    .Q_N(_0599_),
    .Q(\vcount[3] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[4]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net136),
    .D(_0089_),
    .Q_N(_0598_),
    .Q(\vcount[4] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[5]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net137),
    .D(_0090_),
    .Q_N(_0597_),
    .Q(\vcount[5] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[6]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net138),
    .D(_0091_),
    .Q_N(_0596_),
    .Q(\vcount[6] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[7]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net139),
    .D(_0092_),
    .Q_N(_0595_),
    .Q(\vcount[7] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[8]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net140),
    .D(_0093_),
    .Q_N(_0594_),
    .Q(\vcount[8] ));
 sg13g2_dfrbp_1 \vga_sync.vga_ypos[9]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net141),
    .D(_0094_),
    .Q_N(_0593_),
    .Q(\vcount[9] ));
 sg13g2_dfrbp_1 \vga_sync.xvisible$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net142),
    .D(_0095_),
    .Q_N(_0592_),
    .Q(\vga_sync.xvisible ));
 sg13g2_dfrbp_1 \vga_sync.yvisible$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net143),
    .D(_0096_),
    .Q_N(_0591_),
    .Q(\vga_sync.yvisible ));
 sg13g2_dfrbp_1 \vscheudler1.blockline[0]$_SDFFE_PP1P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net144),
    .D(_0097_),
    .Q_N(_0590_),
    .Q(\vscheudler1.blockline[0] ));
 sg13g2_dfrbp_1 \vscheudler1.blockline[1]$_SDFFE_PP1P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net145),
    .D(_0098_),
    .Q_N(_0589_),
    .Q(\vscheudler1.blockline[1] ));
 sg13g2_dfrbp_1 \vscheudler1.blockline[2]$_SDFFE_PP1P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net146),
    .D(_0099_),
    .Q_N(_0588_),
    .Q(\vscheudler1.blockline[2] ));
 sg13g2_dfrbp_1 \vscheudler1.blockline[3]$_SDFFE_PP1P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net147),
    .D(_0100_),
    .Q_N(_0587_),
    .Q(\vscheudler1.blockline[3] ));
 sg13g2_dfrbp_1 \vscheudler1.blockline[4]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net148),
    .D(_0101_),
    .Q_N(_0000_),
    .Q(\vscheudler1.blockline[4] ));
 sg13g2_dfrbp_1 \vscheudler1.blockval[0]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net149),
    .D(_0102_),
    .Q_N(_0007_),
    .Q(\cutoff1[0] ));
 sg13g2_dfrbp_1 \vscheudler1.blockval[1]$_SDFFE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net150),
    .D(_0103_),
    .Q_N(_0586_),
    .Q(\cutoff1[1] ));
 sg13g2_dfrbp_1 \vscheudler1.blockval[2]$_SDFFE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net151),
    .D(_0104_),
    .Q_N(_0585_),
    .Q(\cutoff1[2] ));
 sg13g2_dfrbp_1 \vscheudler1.blockval[3]$_SDFFE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net152),
    .D(_0105_),
    .Q_N(_0584_),
    .Q(\cutoff1[3] ));
 sg13g2_dfrbp_1 \vscheudler1.blockval[4]$_SDFFE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net153),
    .D(_0106_),
    .Q_N(_0583_),
    .Q(\cutoff1[4] ));
 sg13g2_dfrbp_1 \vscheudler1.borderreg$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net154),
    .D(_0107_),
    .Q_N(_0582_),
    .Q(vborder1));
 sg13g2_dfrbp_1 \vscheudler1.started$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net155),
    .D(_0108_),
    .Q_N(_0581_),
    .Q(\vscheudler1.started ));
 sg13g2_dfrbp_1 \vscheudler2.blockline[0]$_SDFFE_PP1P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net156),
    .D(_0109_),
    .Q_N(_0580_),
    .Q(\vscheudler2.blockline[0] ));
 sg13g2_dfrbp_1 \vscheudler2.blockline[1]$_SDFFE_PP1P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net157),
    .D(_0110_),
    .Q_N(_0579_),
    .Q(\vscheudler2.blockline[1] ));
 sg13g2_dfrbp_1 \vscheudler2.blockline[2]$_SDFFE_PP1P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net158),
    .D(_0111_),
    .Q_N(_0578_),
    .Q(\vscheudler2.blockline[2] ));
 sg13g2_dfrbp_1 \vscheudler2.blockline[3]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net159),
    .D(_0112_),
    .Q_N(_0577_),
    .Q(\vscheudler2.blockline[3] ));
 sg13g2_dfrbp_1 \vscheudler2.blockline[4]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net160),
    .D(_0113_),
    .Q_N(_0001_),
    .Q(\vscheudler2.blockline[4] ));
 sg13g2_dfrbp_1 \vscheudler2.blockval[0]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net161),
    .D(_0114_),
    .Q_N(_0006_),
    .Q(\cutoff2[0] ));
 sg13g2_dfrbp_1 \vscheudler2.blockval[1]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net162),
    .D(_0115_),
    .Q_N(_0576_),
    .Q(\cutoff2[1] ));
 sg13g2_dfrbp_1 \vscheudler2.blockval[2]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net163),
    .D(_0116_),
    .Q_N(_0575_),
    .Q(\cutoff2[2] ));
 sg13g2_dfrbp_1 \vscheudler2.blockval[3]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net164),
    .D(_0117_),
    .Q_N(_0574_),
    .Q(\cutoff2[3] ));
 sg13g2_dfrbp_1 \vscheudler2.blockval[4]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net165),
    .D(_0118_),
    .Q_N(_0002_),
    .Q(\cutoff2[4] ));
 sg13g2_dfrbp_1 \vscheudler2.borderreg$_SDFFE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net166),
    .D(_0119_),
    .Q_N(_0573_),
    .Q(vborder2));
 sg13g2_dfrbp_1 \vscheudler2.started$_SDFFE_PP0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net167),
    .D(_0120_),
    .Q_N(_0572_),
    .Q(\vscheudler2.started ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_0540_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0324_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0155_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0496_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0468_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0443_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0417_),
    .X(net16));
 sg13g2_buf_1 fanout17 (.A(_0414_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0367_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0338_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0327_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0326_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0284_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0272_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0185_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0180_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0273_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0214_),
    .X(net27));
 sg13g2_buf_4 fanout28 (.X(net28),
    .A(_0378_));
 sg13g2_buf_2 fanout29 (.A(_0498_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0493_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0399_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0332_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0199_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0178_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0123_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0428_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0341_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0331_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0315_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0227_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0121_),
    .X(net41));
 sg13g2_tielo _1236__42 (.L_LO(net42));
 sg13g2_tielo _1237__43 (.L_LO(net43));
 sg13g2_tielo _1238__44 (.L_LO(net44));
 sg13g2_tielo _1239__45 (.L_LO(net45));
 sg13g2_tielo _1240__46 (.L_LO(net46));
 sg13g2_tielo _1241__47 (.L_LO(net47));
 sg13g2_tielo _1242__48 (.L_LO(net48));
 sg13g2_tielo _1243__49 (.L_LO(net49));
 sg13g2_tielo _1244__50 (.L_LO(net50));
 sg13g2_tielo _1245__51 (.L_LO(net51));
 sg13g2_tielo _1246__52 (.L_LO(net52));
 sg13g2_tielo _1247__53 (.L_LO(net53));
 sg13g2_tielo _1248__54 (.L_LO(net54));
 sg13g2_tielo _1249__55 (.L_LO(net55));
 sg13g2_tielo _1250__56 (.L_LO(net56));
 sg13g2_tielo _1251__57 (.L_LO(net57));
 sg13g2_tiehi \bd[1]$_SDFF_PN0__59  (.L_HI(net59));
 sg13g2_tiehi \bd[2]$_SDFF_PN0__60  (.L_HI(net60));
 sg13g2_tiehi \color_ditherer.bout[0]$_SDFF_PN0__61  (.L_HI(net61));
 sg13g2_tiehi \color_ditherer.bout[1]$_SDFF_PN0__62  (.L_HI(net62));
 sg13g2_tiehi \color_ditherer.gout[0]$_SDFF_PN0__63  (.L_HI(net63));
 sg13g2_tiehi \color_ditherer.gout[1]$_SDFF_PN0__64  (.L_HI(net64));
 sg13g2_tiehi \count1[0]$_SDFFE_PN1P__65  (.L_HI(net65));
 sg13g2_tiehi \count1[1]$_SDFFE_PN1P__66  (.L_HI(net66));
 sg13g2_tiehi \count1[2]$_SDFFE_PN1P__67  (.L_HI(net67));
 sg13g2_tiehi \count1b[0]$_SDFFE_PN1P__68  (.L_HI(net68));
 sg13g2_tiehi \count1b[1]$_SDFFE_PN1P__69  (.L_HI(net69));
 sg13g2_tiehi \count1b[2]$_SDFFE_PN1P__70  (.L_HI(net70));
 sg13g2_tiehi \count2[0]$_SDFFE_PN1P__71  (.L_HI(net71));
 sg13g2_tiehi \count2[1]$_SDFFE_PN1P__72  (.L_HI(net72));
 sg13g2_tiehi \count2b[0]$_SDFFE_PN1P__73  (.L_HI(net73));
 sg13g2_tiehi \count2b[1]$_SDFFE_PN1P__74  (.L_HI(net74));
 sg13g2_tiehi \count2low$_SDFFE_PN1P__75  (.L_HI(net75));
 sg13g2_tiehi \dither$_SDFFE_PN0P__76  (.L_HI(net76));
 sg13g2_tiehi \lfsr1[0]$_SDFFE_PN1P__77  (.L_HI(net77));
 sg13g2_tiehi \lfsr1[1]$_SDFFE_PN1P__78  (.L_HI(net78));
 sg13g2_tiehi \lfsr1[2]$_SDFFE_PN1P__79  (.L_HI(net79));
 sg13g2_tiehi \lfsr1[3]$_SDFFE_PN1P__80  (.L_HI(net80));
 sg13g2_tiehi \lfsr1[4]$_SDFFE_PN1P__81  (.L_HI(net81));
 sg13g2_tiehi \lfsr1[5]$_SDFFE_PN1P__82  (.L_HI(net82));
 sg13g2_tiehi \lfsr1[6]$_SDFFE_PN1P__83  (.L_HI(net83));
 sg13g2_tiehi \lfsr1[7]$_SDFFE_PN1P__84  (.L_HI(net84));
 sg13g2_tiehi \lfsr1[8]$_SDFFE_PN1P__85  (.L_HI(net85));
 sg13g2_tiehi \lfsr1[9]$_SDFFE_PN1P__86  (.L_HI(net86));
 sg13g2_tiehi \lfsr1b[0]$_SDFFE_PN1P__87  (.L_HI(net87));
 sg13g2_tiehi \lfsr1b[1]$_SDFFE_PN1P__88  (.L_HI(net88));
 sg13g2_tiehi \lfsr1b[2]$_SDFFE_PN1P__89  (.L_HI(net89));
 sg13g2_tiehi \lfsr1b[3]$_SDFFE_PN1P__90  (.L_HI(net90));
 sg13g2_tiehi \lfsr1b[4]$_SDFFE_PN1P__91  (.L_HI(net91));
 sg13g2_tiehi \lfsr1b[5]$_SDFFE_PN1P__92  (.L_HI(net92));
 sg13g2_tiehi \lfsr1b[6]$_SDFFE_PN1P__93  (.L_HI(net93));
 sg13g2_tiehi \lfsr1b[7]$_SDFFE_PN1P__94  (.L_HI(net94));
 sg13g2_tiehi \lfsr1b[8]$_SDFFE_PN1P__95  (.L_HI(net95));
 sg13g2_tiehi \lfsr1b[9]$_SDFFE_PN1P__96  (.L_HI(net96));
 sg13g2_tiehi \lfsr2[0]$_SDFFE_PN1P__97  (.L_HI(net97));
 sg13g2_tiehi \lfsr2[1]$_SDFFE_PN1P__98  (.L_HI(net98));
 sg13g2_tiehi \lfsr2[2]$_SDFFE_PN1P__99  (.L_HI(net99));
 sg13g2_tiehi \lfsr2[3]$_SDFFE_PN1P__100  (.L_HI(net100));
 sg13g2_tiehi \lfsr2[4]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \lfsr2[5]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \lfsr2[6]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \lfsr2[7]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \lfsr2[8]$_SDFFE_PN1P__105  (.L_HI(net105));
 sg13g2_tiehi \lfsr2[9]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \lfsr2b[0]$_SDFFE_PN1P__107  (.L_HI(net107));
 sg13g2_tiehi \lfsr2b[1]$_SDFFE_PN1P__108  (.L_HI(net108));
 sg13g2_tiehi \lfsr2b[2]$_SDFFE_PN1P__109  (.L_HI(net109));
 sg13g2_tiehi \lfsr2b[3]$_SDFFE_PN1P__110  (.L_HI(net110));
 sg13g2_tiehi \lfsr2b[4]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \lfsr2b[5]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \lfsr2b[6]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \lfsr2b[7]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \lfsr2b[8]$_SDFFE_PN1P__115  (.L_HI(net115));
 sg13g2_tiehi \lfsr2b[9]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \rd[0]$_SDFF_PP0__117  (.L_HI(net117));
 sg13g2_tiehi \rd[1]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \rd[2]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \vga_sync.vga_hsync$_SDFFE_PN1P__120  (.L_HI(net120));
 sg13g2_tiehi \vga_sync.vga_vsync$_SDFFE_PN1P__121  (.L_HI(net121));
 sg13g2_tiehi \vga_sync.vga_xpos[0]$_SDFF_PP1__122  (.L_HI(net122));
 sg13g2_tiehi \vga_sync.vga_xpos[1]$_SDFF_PP0__123  (.L_HI(net123));
 sg13g2_tiehi \vga_sync.vga_xpos[2]$_SDFF_PP0__124  (.L_HI(net124));
 sg13g2_tiehi \vga_sync.vga_xpos[3]$_SDFF_PP0__125  (.L_HI(net125));
 sg13g2_tiehi \vga_sync.vga_xpos[4]$_SDFF_PP0__126  (.L_HI(net126));
 sg13g2_tiehi \vga_sync.vga_xpos[5]$_SDFF_PP0__127  (.L_HI(net127));
 sg13g2_tiehi \vga_sync.vga_xpos[6]$_SDFF_PP0__128  (.L_HI(net128));
 sg13g2_tiehi \vga_sync.vga_xpos[7]$_SDFF_PP0__129  (.L_HI(net129));
 sg13g2_tiehi \vga_sync.vga_xpos[8]$_SDFF_PP0__130  (.L_HI(net130));
 sg13g2_tiehi \vga_sync.vga_xpos[9]$_SDFF_PP0__131  (.L_HI(net131));
 sg13g2_tiehi \vga_sync.vga_ypos[0]$_SDFFE_PN1N__132  (.L_HI(net132));
 sg13g2_tiehi \vga_sync.vga_ypos[1]$_SDFFE_PN0N__133  (.L_HI(net133));
 sg13g2_tiehi \vga_sync.vga_ypos[2]$_SDFFE_PN0N__134  (.L_HI(net134));
 sg13g2_tiehi \vga_sync.vga_ypos[3]$_SDFFE_PN0N__135  (.L_HI(net135));
 sg13g2_tiehi \vga_sync.vga_ypos[4]$_SDFFE_PN0N__136  (.L_HI(net136));
 sg13g2_tiehi \vga_sync.vga_ypos[5]$_SDFFE_PN0N__137  (.L_HI(net137));
 sg13g2_tiehi \vga_sync.vga_ypos[6]$_SDFFE_PN0N__138  (.L_HI(net138));
 sg13g2_tiehi \vga_sync.vga_ypos[7]$_SDFFE_PN0N__139  (.L_HI(net139));
 sg13g2_tiehi \vga_sync.vga_ypos[8]$_SDFFE_PN0N__140  (.L_HI(net140));
 sg13g2_tiehi \vga_sync.vga_ypos[9]$_SDFFE_PN0N__141  (.L_HI(net141));
 sg13g2_tiehi \vga_sync.xvisible$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \vga_sync.yvisible$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \vscheudler1.blockline[0]$_SDFFE_PP1P__144  (.L_HI(net144));
 sg13g2_tiehi \vscheudler1.blockline[1]$_SDFFE_PP1P__145  (.L_HI(net145));
 sg13g2_tiehi \vscheudler1.blockline[2]$_SDFFE_PP1P__146  (.L_HI(net146));
 sg13g2_tiehi \vscheudler1.blockline[3]$_SDFFE_PP1P__147  (.L_HI(net147));
 sg13g2_tiehi \vscheudler1.blockline[4]$_SDFFE_PP0P__148  (.L_HI(net148));
 sg13g2_tiehi \vscheudler1.blockval[0]$_SDFFE_PP0P__149  (.L_HI(net149));
 sg13g2_tiehi \vscheudler1.blockval[1]$_SDFFE_PP0P__150  (.L_HI(net150));
 sg13g2_tiehi \vscheudler1.blockval[2]$_SDFFE_PP0P__151  (.L_HI(net151));
 sg13g2_tiehi \vscheudler1.blockval[3]$_SDFFE_PP0P__152  (.L_HI(net152));
 sg13g2_tiehi \vscheudler1.blockval[4]$_SDFFE_PP0P__153  (.L_HI(net153));
 sg13g2_tiehi \vscheudler1.borderreg$_SDFFE_PP0P__154  (.L_HI(net154));
 sg13g2_tiehi \vscheudler1.started$_SDFFE_PP0N__155  (.L_HI(net155));
 sg13g2_tiehi \vscheudler2.blockline[0]$_SDFFE_PP1P__156  (.L_HI(net156));
 sg13g2_tiehi \vscheudler2.blockline[1]$_SDFFE_PP1P__157  (.L_HI(net157));
 sg13g2_tiehi \vscheudler2.blockline[2]$_SDFFE_PP1P__158  (.L_HI(net158));
 sg13g2_tiehi \vscheudler2.blockline[3]$_SDFFE_PP0P__159  (.L_HI(net159));
 sg13g2_tiehi \vscheudler2.blockline[4]$_SDFFE_PP0P__160  (.L_HI(net160));
 sg13g2_tiehi \vscheudler2.blockval[0]$_SDFFE_PP0P__161  (.L_HI(net161));
 sg13g2_tiehi \vscheudler2.blockval[1]$_SDFFE_PP0P__162  (.L_HI(net162));
 sg13g2_tiehi \vscheudler2.blockval[2]$_SDFFE_PP0P__163  (.L_HI(net163));
 sg13g2_tiehi \vscheudler2.blockval[3]$_SDFFE_PP0P__164  (.L_HI(net164));
 sg13g2_tiehi \vscheudler2.blockval[4]$_SDFFE_PP0P__165  (.L_HI(net165));
 sg13g2_tiehi \vscheudler2.borderreg$_SDFFE_PP0P__166  (.L_HI(net166));
 sg13g2_tiehi \vscheudler2.started$_SDFFE_PP0N__167  (.L_HI(net167));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_decap_4 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_decap_8 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_194 ();
 sg13g2_decap_8 FILLER_12_201 ();
 sg13g2_fill_2 FILLER_12_208 ();
 sg13g2_fill_1 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_decap_8 FILLER_12_229 ();
 sg13g2_decap_8 FILLER_12_236 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_164 ();
 sg13g2_decap_8 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_192 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_269 ();
 sg13g2_decap_8 FILLER_13_276 ();
 sg13g2_decap_8 FILLER_13_283 ();
 sg13g2_decap_8 FILLER_13_290 ();
 sg13g2_decap_8 FILLER_13_297 ();
 sg13g2_decap_8 FILLER_13_304 ();
 sg13g2_decap_8 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_13_409 ();
 sg13g2_decap_8 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_114 ();
 sg13g2_fill_2 FILLER_14_130 ();
 sg13g2_fill_1 FILLER_14_132 ();
 sg13g2_decap_4 FILLER_14_137 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_decap_4 FILLER_14_204 ();
 sg13g2_decap_4 FILLER_14_220 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_404 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_163 ();
 sg13g2_decap_4 FILLER_15_170 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_4 FILLER_15_223 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_276 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_fill_2 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_fill_1 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_fill_1 FILLER_16_135 ();
 sg13g2_decap_4 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_177 ();
 sg13g2_decap_4 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_fill_1 FILLER_16_245 ();
 sg13g2_fill_2 FILLER_16_254 ();
 sg13g2_fill_1 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_fill_2 FILLER_16_340 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_16_413 ();
 sg13g2_fill_2 FILLER_16_417 ();
 sg13g2_decap_4 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_4 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_99 ();
 sg13g2_decap_8 FILLER_17_106 ();
 sg13g2_decap_4 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_decap_4 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_160 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_fill_2 FILLER_17_199 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_decap_4 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_61 ();
 sg13g2_decap_4 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_decap_8 FILLER_18_82 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_125 ();
 sg13g2_decap_4 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_186 ();
 sg13g2_decap_4 FILLER_18_195 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_4 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_4 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_decap_4 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_370 ();
 sg13g2_fill_1 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_16 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_39 ();
 sg13g2_fill_1 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_100 ();
 sg13g2_decap_8 FILLER_19_107 ();
 sg13g2_fill_2 FILLER_19_124 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_222 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_4 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_4 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_4 FILLER_19_332 ();
 sg13g2_fill_2 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_fill_2 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_fill_1 FILLER_19_394 ();
 sg13g2_decap_4 FILLER_19_402 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_decap_8 FILLER_20_57 ();
 sg13g2_decap_4 FILLER_20_64 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_fill_2 FILLER_20_113 ();
 sg13g2_decap_4 FILLER_20_152 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_230 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_4 FILLER_20_366 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_43 ();
 sg13g2_decap_8 FILLER_21_103 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_decap_4 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_decap_4 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_167 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_decap_4 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_387 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_19 ();
 sg13g2_decap_8 FILLER_22_26 ();
 sg13g2_decap_8 FILLER_22_33 ();
 sg13g2_decap_8 FILLER_22_40 ();
 sg13g2_decap_4 FILLER_22_47 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_decap_4 FILLER_22_61 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_111 ();
 sg13g2_decap_4 FILLER_22_118 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_decap_4 FILLER_22_150 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_decap_4 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_229 ();
 sg13g2_decap_8 FILLER_22_234 ();
 sg13g2_decap_4 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_349 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_419 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_decap_4 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_decap_8 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_118 ();
 sg13g2_decap_4 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_fill_2 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_192 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_decap_8 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_decap_4 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_4 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_fill_2 FILLER_24_32 ();
 sg13g2_fill_1 FILLER_24_34 ();
 sg13g2_decap_4 FILLER_24_73 ();
 sg13g2_decap_4 FILLER_24_85 ();
 sg13g2_fill_2 FILLER_24_95 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_decap_4 FILLER_24_222 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_decap_4 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_fill_2 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_4 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_41 ();
 sg13g2_decap_4 FILLER_25_47 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_99 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_decap_4 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_decap_4 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_397 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_fill_1 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_20 ();
 sg13g2_decap_8 FILLER_26_27 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_69 ();
 sg13g2_fill_2 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_decap_4 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_2 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_decap_4 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_376 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_44 ();
 sg13g2_decap_8 FILLER_27_51 ();
 sg13g2_decap_4 FILLER_27_58 ();
 sg13g2_fill_2 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_97 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_decap_4 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_129 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_decap_4 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_decap_4 FILLER_27_216 ();
 sg13g2_decap_4 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_decap_4 FILLER_27_255 ();
 sg13g2_decap_4 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_8 ();
 sg13g2_fill_1 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_decap_8 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_decap_4 FILLER_28_100 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_fill_2 FILLER_28_232 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_4 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_25 ();
 sg13g2_fill_2 FILLER_29_37 ();
 sg13g2_fill_2 FILLER_29_43 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_decap_4 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_decap_4 FILLER_29_89 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_4 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_decap_4 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_124 ();
 sg13g2_decap_8 FILLER_29_131 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_decap_4 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_149 ();
 sg13g2_decap_4 FILLER_29_155 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_decap_4 FILLER_29_267 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_decap_4 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_409 ();
 sg13g2_decap_8 FILLER_29_416 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_18 ();
 sg13g2_decap_4 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_33 ();
 sg13g2_decap_4 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_fill_2 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_decap_8 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_213 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_decap_4 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_155 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_236 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_decap_4 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_4 FILLER_31_366 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_4 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_decap_4 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_decap_8 FILLER_32_72 ();
 sg13g2_decap_8 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_4 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_decap_4 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_fill_1 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_24 ();
 sg13g2_decap_8 FILLER_33_31 ();
 sg13g2_decap_8 FILLER_33_38 ();
 sg13g2_decap_8 FILLER_33_45 ();
 sg13g2_decap_8 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_92 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_decap_4 FILLER_33_177 ();
 sg13g2_decap_4 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_decap_8 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_411 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_15 ();
 sg13g2_fill_1 FILLER_34_19 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_2 FILLER_34_32 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_57 ();
 sg13g2_decap_4 FILLER_34_69 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_89 ();
 sg13g2_decap_8 FILLER_34_101 ();
 sg13g2_decap_4 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_261 ();
 sg13g2_decap_4 FILLER_34_268 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_decap_4 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_370 ();
 sg13g2_fill_1 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_75 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_decap_4 FILLER_35_89 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_4 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_decap_4 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_179 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_353 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_35_417 ();
 sg13g2_decap_4 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_decap_8 FILLER_36_45 ();
 sg13g2_decap_8 FILLER_36_52 ();
 sg13g2_decap_4 FILLER_36_59 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_97 ();
 sg13g2_decap_8 FILLER_36_108 ();
 sg13g2_decap_8 FILLER_36_115 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_decap_8 FILLER_36_129 ();
 sg13g2_decap_8 FILLER_36_136 ();
 sg13g2_decap_8 FILLER_36_143 ();
 sg13g2_decap_8 FILLER_36_150 ();
 sg13g2_decap_4 FILLER_36_157 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_decap_8 FILLER_36_257 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_367 ();
 sg13g2_fill_1 FILLER_36_369 ();
 sg13g2_fill_2 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_4 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_decap_4 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_4 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_decap_8 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_288 ();
 sg13g2_decap_4 FILLER_38_295 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_318 ();
 sg13g2_decap_8 FILLER_38_325 ();
 sg13g2_decap_8 FILLER_38_332 ();
 sg13g2_decap_8 FILLER_38_339 ();
 sg13g2_decap_8 FILLER_38_346 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_decap_8 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_8 FILLER_38_404 ();
 sg13g2_decap_8 FILLER_38_411 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
