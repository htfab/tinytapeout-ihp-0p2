module tt_um_algofoogle_vga_fun_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire clknet_0_clk;
 wire net80;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[28] ;
 wire \counter[29] ;
 wire \counter[2] ;
 wire \counter[30] ;
 wire \counter[31] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \depth[0] ;
 wire \depth[1] ;
 wire \depth[2] ;
 wire hsync;
 wire \i_project.controller_0.divider[0] ;
 wire \i_project.controller_0.divider[1] ;
 wire \i_project.controller_0.grey_pass[10] ;
 wire \i_project.controller_0.grey_pass[11] ;
 wire \i_project.controller_0.grey_pass[12] ;
 wire \i_project.controller_0.grey_pass[13] ;
 wire \i_project.controller_0.grey_pass[14] ;
 wire \i_project.controller_0.grey_pass[15] ;
 wire \i_project.controller_0.h[0] ;
 wire \i_project.controller_0.h[1] ;
 wire \i_project.controller_0.h[2] ;
 wire \i_project.controller_0.h[3] ;
 wire \i_project.controller_0.h[4] ;
 wire \i_project.controller_0.h[5] ;
 wire \i_project.controller_0.h[6] ;
 wire \i_project.controller_0.h[7] ;
 wire \i_project.controller_0.h[8] ;
 wire \i_project.controller_0.h[9] ;
 wire \i_project.controller_0.mode[0] ;
 wire \i_project.controller_0.mode[1] ;
 wire \i_project.controller_0.mode[2] ;
 wire \i_project.controller_0.mode_ramp_base[0] ;
 wire \i_project.controller_0.mode_ramp_base[1] ;
 wire \i_project.controller_0.mode_ramp_base[2] ;
 wire \i_project.controller_0.mode_ramp_base[3] ;
 wire \i_project.controller_0.mode_ramp_base[4] ;
 wire \i_project.controller_0.mode_ramp_base[5] ;
 wire \i_project.controller_0.mode_ramp_base[6] ;
 wire \i_project.controller_0.mode_ramp_base[7] ;
 wire \i_project.controller_0.rst_n ;
 wire \i_project.controller_0.t[10] ;
 wire \i_project.controller_0.t[11] ;
 wire \i_project.controller_0.t[8] ;
 wire \i_project.controller_0.t[9] ;
 wire \i_project.controller_0.v[0] ;
 wire \i_project.controller_0.v[1] ;
 wire \i_project.controller_0.v[2] ;
 wire \i_project.controller_0.v[3] ;
 wire \i_project.controller_0.v[4] ;
 wire \i_project.controller_0.v[5] ;
 wire \i_project.controller_0.v[6] ;
 wire \i_project.controller_0.v[7] ;
 wire \i_project.controller_0.v[8] ;
 wire \i_project.controller_0.v[9] ;
 wire \i_project.controller_0.vga_sync.hsync ;
 wire \i_project.controller_0.vga_sync.mode ;
 wire \i_project.controller_0.vga_sync.o_vsync ;
 wire \i_project.controller_0.vga_sync.vsync ;
 wire \i_project.controller_0.voffset[0] ;
 wire \i_project.controller_0.voffset[1] ;
 wire \i_project.controller_0.voffset[2] ;
 wire \i_project.controller_0.voffset[3] ;
 wire \i_project.controller_0.voffset[4] ;
 wire \i_project.controller_0.voffset[5] ;
 wire \i_project.controller_0.voffset[6] ;
 wire \i_project.controller_0.voffset[7] ;
 wire \lfsr[0] ;
 wire \lfsr[10] ;
 wire \lfsr[11] ;
 wire \lfsr[12] ;
 wire \lfsr[13] ;
 wire \lfsr[14] ;
 wire \lfsr[15] ;
 wire \lfsr[16] ;
 wire \lfsr[17] ;
 wire \lfsr[18] ;
 wire \lfsr[19] ;
 wire \lfsr[1] ;
 wire \lfsr[20] ;
 wire \lfsr[21] ;
 wire \lfsr[22] ;
 wire \lfsr[23] ;
 wire \lfsr[24] ;
 wire \lfsr[25] ;
 wire \lfsr[26] ;
 wire \lfsr[27] ;
 wire \lfsr[28] ;
 wire \lfsr[29] ;
 wire \lfsr[2] ;
 wire \lfsr[30] ;
 wire \lfsr[31] ;
 wire \lfsr[3] ;
 wire \lfsr[4] ;
 wire \lfsr[5] ;
 wire \lfsr[6] ;
 wire \lfsr[7] ;
 wire \lfsr[8] ;
 wire \lfsr[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_a21oi_1 _1989_ (.A1(_0637_),
    .A2(net48),
    .Y(_1110_),
    .B1(net35));
 sg13g2_nand2_1 _1990_ (.Y(_1111_),
    .A(_1109_),
    .B(_1110_));
 sg13g2_nand2_1 _1991_ (.Y(_1112_),
    .A(_1111_),
    .B(_0246_));
 sg13g2_nand2_1 _1992_ (.Y(_1113_),
    .A(_1112_),
    .B(_0248_));
 sg13g2_nand4_1 _1993_ (.B(_0259_),
    .C(_0270_),
    .A(_1113_),
    .Y(_1114_),
    .D(_0261_));
 sg13g2_nand2_1 _1994_ (.Y(_1115_),
    .A(_1114_),
    .B(_0375_));
 sg13g2_nand3_1 _1995_ (.B(_0313_),
    .C(_0319_),
    .A(_1080_),
    .Y(_1116_));
 sg13g2_xnor2_1 _1996_ (.Y(_1117_),
    .A(_0987_),
    .B(_0982_));
 sg13g2_nand2_1 _1997_ (.Y(_1118_),
    .A(_1087_),
    .B(_1117_));
 sg13g2_nand3_1 _1998_ (.B(_1015_),
    .C(_0979_),
    .A(_1086_),
    .Y(_1119_));
 sg13g2_nand3_1 _1999_ (.B(_1119_),
    .C(net49),
    .A(_1118_),
    .Y(_1120_));
 sg13g2_a21o_1 _2000_ (.A2(_1061_),
    .A1(_1059_),
    .B1(_1049_),
    .X(_1121_));
 sg13g2_xnor2_1 _2001_ (.Y(_1122_),
    .A(_1052_),
    .B(_1121_));
 sg13g2_inv_1 _2002_ (.Y(_1123_),
    .A(_1040_));
 sg13g2_a21o_1 _2003_ (.A2(_1041_),
    .A1(_1039_),
    .B1(_1029_),
    .X(_1124_));
 sg13g2_xnor2_1 _2004_ (.Y(_1125_),
    .A(_1123_),
    .B(_1124_));
 sg13g2_nor2_1 _2005_ (.A(_1122_),
    .B(_1125_),
    .Y(_1126_));
 sg13g2_a21oi_1 _2006_ (.A1(_1125_),
    .A2(_1122_),
    .Y(_1127_),
    .B1(_0293_));
 sg13g2_nand2b_1 _2007_ (.Y(_1128_),
    .B(_1127_),
    .A_N(_1126_));
 sg13g2_nand2_1 _2008_ (.Y(_1129_),
    .A(_1128_),
    .B(_0846_));
 sg13g2_nand3_1 _2009_ (.B(_1129_),
    .C(_0363_),
    .A(_1120_),
    .Y(_1130_));
 sg13g2_xor2_1 _2010_ (.B(_0200_),
    .A(_1698_),
    .X(_1131_));
 sg13g2_a21oi_1 _2011_ (.A1(_1131_),
    .A2(_0303_),
    .Y(_1132_),
    .B1(net42));
 sg13g2_nand2_1 _2012_ (.Y(_1133_),
    .A(_1130_),
    .B(_1132_));
 sg13g2_a21oi_1 _2013_ (.A1(_1863_),
    .A2(_0304_),
    .Y(_1134_),
    .B1(net29));
 sg13g2_nand2_1 _2014_ (.Y(_1135_),
    .A(_1133_),
    .B(_1134_));
 sg13g2_a21oi_1 _2015_ (.A1(_1135_),
    .A2(net22),
    .Y(_1136_),
    .B1(net52));
 sg13g2_nor2_1 _2016_ (.A(_0331_),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_nand2b_1 _2017_ (.Y(_1138_),
    .B(_1137_),
    .A_N(_0339_));
 sg13g2_nand2_1 _2018_ (.Y(_1139_),
    .A(_1116_),
    .B(_1138_));
 sg13g2_nor2_1 _2019_ (.A(_1115_),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_nor2_1 _2020_ (.A(_1083_),
    .B(_1140_),
    .Y(_1141_));
 sg13g2_inv_1 _2021_ (.Y(_1142_),
    .A(_1141_));
 sg13g2_inv_4 _2022_ (.A(_1081_),
    .Y(_1143_));
 sg13g2_nand2_1 _2023_ (.Y(_1144_),
    .A(_0266_),
    .B(_0043_));
 sg13g2_inv_1 _2024_ (.Y(_1145_),
    .A(_1144_));
 sg13g2_nand3_1 _2025_ (.B(_0259_),
    .C(_0261_),
    .A(_1113_),
    .Y(_1146_));
 sg13g2_nor2_1 _2026_ (.A(_0413_),
    .B(_1146_),
    .Y(_1147_));
 sg13g2_inv_1 _2027_ (.Y(_1148_),
    .A(_1147_));
 sg13g2_nand2b_1 _2028_ (.Y(_1149_),
    .B(_1014_),
    .A_N(_1011_));
 sg13g2_nand3_1 _2029_ (.B(net46),
    .C(_1086_),
    .A(_1149_),
    .Y(_1150_));
 sg13g2_o21ai_1 _2030_ (.B1(_1046_),
    .Y(_1151_),
    .A1(_1058_),
    .A2(_1060_));
 sg13g2_xnor2_1 _2031_ (.Y(_1152_),
    .A(_1047_),
    .B(_1151_));
 sg13g2_xor2_1 _2032_ (.B(_1039_),
    .A(_1041_),
    .X(_1153_));
 sg13g2_xor2_1 _2033_ (.B(_1153_),
    .A(_1152_),
    .X(_1154_));
 sg13g2_o21ai_1 _2034_ (.B1(_0760_),
    .Y(_1155_),
    .A1(net39),
    .A2(_1154_));
 sg13g2_nand3_1 _2035_ (.B(net33),
    .C(_1155_),
    .A(_1150_),
    .Y(_1156_));
 sg13g2_a21oi_1 _2036_ (.A1(net23),
    .A2(_1696_),
    .Y(_1157_),
    .B1(net33));
 sg13g2_o21ai_1 _2037_ (.B1(_1157_),
    .Y(_1158_),
    .A1(_1696_),
    .A2(net23));
 sg13g2_nand3_1 _2038_ (.B(net38),
    .C(_1158_),
    .A(_1156_),
    .Y(_1159_));
 sg13g2_nand2_1 _2039_ (.Y(_1160_),
    .A(net32),
    .B(_0968_));
 sg13g2_nand3_1 _2040_ (.B(_0420_),
    .C(_1160_),
    .A(_1159_),
    .Y(_1161_));
 sg13g2_a21o_1 _2041_ (.A2(_0309_),
    .A1(_1161_),
    .B1(net52),
    .X(_1162_));
 sg13g2_a21oi_1 _2042_ (.A1(_1162_),
    .A2(_0521_),
    .Y(_1163_),
    .B1(_0329_));
 sg13g2_nand2_1 _2043_ (.Y(_1164_),
    .A(_1148_),
    .B(_1163_));
 sg13g2_a21oi_1 _2044_ (.A1(_1143_),
    .A2(_1145_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_nor3_1 _2045_ (.A(net30),
    .B(_1143_),
    .C(_1165_),
    .Y(_1166_));
 sg13g2_a21o_1 _2046_ (.A2(_1165_),
    .A1(_1143_),
    .B1(_1166_),
    .X(_1167_));
 sg13g2_xnor2_1 _2047_ (.Y(_1168_),
    .A(net58),
    .B(_0974_));
 sg13g2_inv_1 _2048_ (.Y(_1169_),
    .A(_1000_));
 sg13g2_nand2_1 _2049_ (.Y(_1170_),
    .A(_1168_),
    .B(_1169_));
 sg13g2_inv_1 _2050_ (.Y(_1171_),
    .A(_1010_));
 sg13g2_a21oi_1 _2051_ (.A1(_1170_),
    .A2(_1008_),
    .Y(_1172_),
    .B1(_1171_));
 sg13g2_nor3_1 _2052_ (.A(_1172_),
    .B(_1014_),
    .C(_1015_),
    .Y(_1173_));
 sg13g2_nor2b_1 _2053_ (.A(_1173_),
    .B_N(_0990_),
    .Y(_1174_));
 sg13g2_nand2b_1 _2054_ (.Y(_1175_),
    .B(_1006_),
    .A_N(_1008_));
 sg13g2_nand2_1 _2055_ (.Y(_1176_),
    .A(_1010_),
    .B(_1170_));
 sg13g2_nor2_1 _2056_ (.A(_1175_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_nand4_1 _2057_ (.B(_1085_),
    .C(_1007_),
    .A(_1117_),
    .Y(_1178_),
    .D(_1177_));
 sg13g2_nand2_1 _2058_ (.Y(_1179_),
    .A(_1174_),
    .B(_1178_));
 sg13g2_inv_1 _2059_ (.Y(_1180_),
    .A(_0958_));
 sg13g2_nand2_1 _2060_ (.Y(_1181_),
    .A(_1179_),
    .B(_1180_));
 sg13g2_nand3_1 _2061_ (.B(_1178_),
    .C(_0958_),
    .A(_1174_),
    .Y(_1182_));
 sg13g2_nand3_1 _2062_ (.B(_1182_),
    .C(net49),
    .A(_1181_),
    .Y(_1183_));
 sg13g2_nand2_1 _2063_ (.Y(_1184_),
    .A(_1121_),
    .B(_1051_));
 sg13g2_nand2_1 _2064_ (.Y(_1185_),
    .A(_1184_),
    .B(_1054_));
 sg13g2_xnor2_1 _2065_ (.Y(_1186_),
    .A(_1050_),
    .B(_1185_));
 sg13g2_nand3_1 _2066_ (.B(_1027_),
    .C(_1031_),
    .A(_1098_),
    .Y(_1187_));
 sg13g2_nand2_1 _2067_ (.Y(_1188_),
    .A(_1100_),
    .B(_1187_));
 sg13g2_nor2_1 _2068_ (.A(_1186_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_a21oi_1 _2069_ (.A1(_1188_),
    .A2(_1186_),
    .Y(_1190_),
    .B1(_0293_));
 sg13g2_nand2b_1 _2070_ (.Y(_1191_),
    .B(_1190_),
    .A_N(_1189_));
 sg13g2_a21oi_1 _2071_ (.A1(_1191_),
    .A2(_0867_),
    .Y(_1192_),
    .B1(_0186_));
 sg13g2_nand2_1 _2072_ (.Y(_1193_),
    .A(_1183_),
    .B(_1192_));
 sg13g2_xnor2_1 _2073_ (.Y(_1194_),
    .A(_1690_),
    .B(net27));
 sg13g2_a21oi_1 _2074_ (.A1(_1194_),
    .A2(_0186_),
    .Y(_1195_),
    .B1(net48));
 sg13g2_nand2_1 _2075_ (.Y(_1196_),
    .A(_1193_),
    .B(_1195_));
 sg13g2_a21oi_1 _2076_ (.A1(_0942_),
    .A2(net48),
    .Y(_1197_),
    .B1(net35));
 sg13g2_nand2_1 _2077_ (.Y(_1198_),
    .A(_1196_),
    .B(_1197_));
 sg13g2_nand2_1 _2078_ (.Y(_1199_),
    .A(_1198_),
    .B(_0246_));
 sg13g2_nand2_1 _2079_ (.Y(_1200_),
    .A(_1199_),
    .B(_0248_));
 sg13g2_nand2_1 _2080_ (.Y(_1201_),
    .A(_1200_),
    .B(_0407_));
 sg13g2_nor2_1 _2081_ (.A(_0339_),
    .B(_1201_),
    .Y(_1202_));
 sg13g2_nor2b_1 _2082_ (.A(_1202_),
    .B_N(_0375_),
    .Y(_1203_));
 sg13g2_nand4_1 _2083_ (.B(_0259_),
    .C(_0319_),
    .A(_1200_),
    .Y(_1204_),
    .D(_0407_));
 sg13g2_nand2_1 _2084_ (.Y(_1205_),
    .A(_1203_),
    .B(_1204_));
 sg13g2_nand2_1 _2085_ (.Y(_1206_),
    .A(_1205_),
    .B(_1082_));
 sg13g2_nand2_1 _2086_ (.Y(_1207_),
    .A(_1143_),
    .B(_0270_));
 sg13g2_nand2_1 _2087_ (.Y(_1208_),
    .A(_1206_),
    .B(_1207_));
 sg13g2_buf_2 _2088_ (.A(_1208_),
    .X(_1209_));
 sg13g2_nor2_1 _2089_ (.A(_0441_),
    .B(_1201_),
    .Y(_1210_));
 sg13g2_xnor2_1 _2090_ (.Y(_1211_),
    .A(_1007_),
    .B(_1175_));
 sg13g2_nand2_1 _2091_ (.Y(_1212_),
    .A(_1211_),
    .B(net46));
 sg13g2_nand2b_1 _2092_ (.Y(_1213_),
    .B(_0432_),
    .A_N(_0427_));
 sg13g2_nand3_1 _2093_ (.B(_0363_),
    .C(_1213_),
    .A(_1212_),
    .Y(_1214_));
 sg13g2_a21oi_1 _2094_ (.A1(_0200_),
    .A2(_1701_),
    .Y(_1215_),
    .B1(_0363_));
 sg13g2_o21ai_1 _2095_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_1701_),
    .A2(net24));
 sg13g2_nand3_1 _2096_ (.B(net38),
    .C(_1216_),
    .A(_1214_),
    .Y(_1217_));
 sg13g2_nand2_1 _2097_ (.Y(_1218_),
    .A(net37),
    .B(_0996_));
 sg13g2_nand3_1 _2098_ (.B(_0420_),
    .C(_1218_),
    .A(_1217_),
    .Y(_1219_));
 sg13g2_a21oi_1 _2099_ (.A1(_0448_),
    .A2(_1219_),
    .Y(_1220_),
    .B1(_0328_));
 sg13g2_nor2b_1 _2100_ (.A(_1210_),
    .B_N(_1220_),
    .Y(_1221_));
 sg13g2_nand2_1 _2101_ (.Y(_1222_),
    .A(_1116_),
    .B(_1221_));
 sg13g2_nor2_1 _2102_ (.A(_0270_),
    .B(_0414_),
    .Y(_1223_));
 sg13g2_nand3b_1 _2103_ (.B(_1080_),
    .C(_0313_),
    .Y(_1224_),
    .A_N(_1223_));
 sg13g2_nor2_2 _2104_ (.A(_0535_),
    .B(_1146_),
    .Y(_1225_));
 sg13g2_inv_2 _2105_ (.Y(_1226_),
    .A(_1225_));
 sg13g2_nand2_1 _2106_ (.Y(_1227_),
    .A(_1224_),
    .B(_1226_));
 sg13g2_nor2_1 _2107_ (.A(_1222_),
    .B(_1227_),
    .Y(_1228_));
 sg13g2_inv_1 _2108_ (.Y(_1229_),
    .A(_1205_));
 sg13g2_nand2_1 _2109_ (.Y(_1230_),
    .A(_1229_),
    .B(_1207_));
 sg13g2_nor2_1 _2110_ (.A(_1230_),
    .B(_1228_),
    .Y(_1231_));
 sg13g2_a21oi_1 _2111_ (.A1(_1209_),
    .A2(_1228_),
    .Y(_1232_),
    .B1(_1231_));
 sg13g2_nand4_1 _2112_ (.B(_0259_),
    .C(_0410_),
    .A(_1200_),
    .Y(_1233_),
    .D(_0407_));
 sg13g2_nor2_1 _2113_ (.A(_1685_),
    .B(_0426_),
    .Y(_1234_));
 sg13g2_nor3_1 _2114_ (.A(_0168_),
    .B(_1234_),
    .C(_1007_),
    .Y(_1235_));
 sg13g2_a21oi_1 _2115_ (.A1(net24),
    .A2(_1685_),
    .Y(_1236_),
    .B1(_0363_));
 sg13g2_o21ai_1 _2116_ (.B1(_1236_),
    .Y(_1237_),
    .A1(_1685_),
    .A2(net24));
 sg13g2_o21ai_1 _2117_ (.B1(_1237_),
    .Y(_1238_),
    .A1(net34),
    .A2(_1235_));
 sg13g2_nand2_1 _2118_ (.Y(_1239_),
    .A(net37),
    .B(_1683_));
 sg13g2_nand3_1 _2119_ (.B(_0420_),
    .C(_1239_),
    .A(_1238_),
    .Y(_1240_));
 sg13g2_a22oi_1 _2120_ (.Y(_1241_),
    .B1(_0338_),
    .B2(_1137_),
    .A2(_1240_),
    .A1(_0818_));
 sg13g2_nand2_1 _2121_ (.Y(_1242_),
    .A(_1233_),
    .B(_1241_));
 sg13g2_nor2_1 _2122_ (.A(_1242_),
    .B(_1115_),
    .Y(_1243_));
 sg13g2_nor2_1 _2123_ (.A(_0415_),
    .B(_1146_),
    .Y(_1244_));
 sg13g2_nor2_1 _2124_ (.A(_0419_),
    .B(_1081_),
    .Y(_1245_));
 sg13g2_nor2_1 _2125_ (.A(_1244_),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_nand3_1 _2126_ (.B(_1148_),
    .C(_1246_),
    .A(_1243_),
    .Y(_1247_));
 sg13g2_inv_1 _2127_ (.Y(_1248_),
    .A(_1247_));
 sg13g2_nand2_1 _2128_ (.Y(_1249_),
    .A(_1248_),
    .B(_1141_));
 sg13g2_nand2_1 _2129_ (.Y(_1250_),
    .A(_1232_),
    .B(_1249_));
 sg13g2_nor2_1 _2130_ (.A(_0535_),
    .B(_1081_),
    .Y(_1251_));
 sg13g2_nand3_1 _2131_ (.B(_0338_),
    .C(_0261_),
    .A(_1113_),
    .Y(_1252_));
 sg13g2_o21ai_1 _2132_ (.B1(net46),
    .Y(_1253_),
    .A1(_1009_),
    .A2(_1176_));
 sg13g2_a21oi_1 _2133_ (.A1(_1176_),
    .A2(_1009_),
    .Y(_1254_),
    .B1(_1253_));
 sg13g2_xnor2_1 _2134_ (.Y(_1255_),
    .A(_1059_),
    .B(_1060_));
 sg13g2_xor2_1 _2135_ (.B(_1035_),
    .A(_1036_),
    .X(_1256_));
 sg13g2_xor2_1 _2136_ (.B(_1256_),
    .A(_1255_),
    .X(_1257_));
 sg13g2_o21ai_1 _2137_ (.B1(_0812_),
    .Y(_1258_),
    .A1(net39),
    .A2(_1257_));
 sg13g2_nand3b_1 _2138_ (.B(net33),
    .C(_1258_),
    .Y(_1259_),
    .A_N(_1254_));
 sg13g2_a21oi_1 _2139_ (.A1(net24),
    .A2(net70),
    .Y(_1260_),
    .B1(net33));
 sg13g2_o21ai_1 _2140_ (.B1(_1260_),
    .Y(_1261_),
    .A1(_1700_),
    .A2(net24));
 sg13g2_nand3_1 _2141_ (.B(net38),
    .C(_1261_),
    .A(_1259_),
    .Y(_1262_));
 sg13g2_nand2b_1 _2142_ (.Y(_1263_),
    .B(net37),
    .A_N(_0042_));
 sg13g2_nand3_1 _2143_ (.B(_0420_),
    .C(_1263_),
    .A(_1262_),
    .Y(_1264_));
 sg13g2_a21oi_1 _2144_ (.A1(_1264_),
    .A2(net22),
    .Y(_1265_),
    .B1(net52));
 sg13g2_nand2b_1 _2145_ (.Y(_1266_),
    .B(_0561_),
    .A_N(_1265_));
 sg13g2_nand3_1 _2146_ (.B(_1252_),
    .C(_1266_),
    .A(_1204_),
    .Y(_1267_));
 sg13g2_nor3_1 _2147_ (.A(_1115_),
    .B(_1251_),
    .C(_1267_),
    .Y(_1268_));
 sg13g2_nand2_1 _2148_ (.Y(_1269_),
    .A(_1113_),
    .B(_0261_));
 sg13g2_o21ai_1 _2149_ (.B1(net26),
    .Y(_1270_),
    .A1(_0837_),
    .A2(_1269_));
 sg13g2_nor2_2 _2150_ (.A(_1225_),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_nor2b_1 _2151_ (.A(_1268_),
    .B_N(_1271_),
    .Y(_1272_));
 sg13g2_nor2_1 _2152_ (.A(_1231_),
    .B(_1272_),
    .Y(_1273_));
 sg13g2_nand2_1 _2153_ (.Y(_1274_),
    .A(_1250_),
    .B(_1273_));
 sg13g2_nor2_2 _2154_ (.A(_1083_),
    .B(_1271_),
    .Y(_1275_));
 sg13g2_nand2_1 _2155_ (.Y(_1276_),
    .A(_1268_),
    .B(_1275_));
 sg13g2_nand2_1 _2156_ (.Y(_1277_),
    .A(_1274_),
    .B(_1276_));
 sg13g2_or2_1 _2157_ (.X(_1278_),
    .B(_1277_),
    .A(_1167_));
 sg13g2_nor2b_1 _2158_ (.A(_1166_),
    .B_N(_1278_),
    .Y(_1279_));
 sg13g2_xnor2_1 _2159_ (.Y(_1280_),
    .A(_1167_),
    .B(_1277_));
 sg13g2_nand2b_1 _2160_ (.Y(_1281_),
    .B(_1276_),
    .A_N(_1272_));
 sg13g2_nand2_1 _2161_ (.Y(_1282_),
    .A(_1209_),
    .B(_1228_));
 sg13g2_a21oi_1 _2162_ (.A1(_1249_),
    .A2(_1282_),
    .Y(_1283_),
    .B1(_1231_));
 sg13g2_xnor2_1 _2163_ (.Y(_1284_),
    .A(_1281_),
    .B(_1283_));
 sg13g2_nand2_1 _2164_ (.Y(_1285_),
    .A(_1247_),
    .B(_1140_));
 sg13g2_and3_1 _2165_ (.X(_1286_),
    .A(_1232_),
    .B(_1249_),
    .C(_1285_));
 sg13g2_nand3_1 _2166_ (.B(_1284_),
    .C(_1286_),
    .A(_1280_),
    .Y(_1287_));
 sg13g2_nor2b_1 _2167_ (.A(_1279_),
    .B_N(_1287_),
    .Y(_1288_));
 sg13g2_inv_1 _2168_ (.Y(_1289_),
    .A(_1222_));
 sg13g2_nor2_1 _2169_ (.A(_1223_),
    .B(_1081_),
    .Y(_1290_));
 sg13g2_nor2_1 _2170_ (.A(_1225_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_nand2_1 _2171_ (.Y(_1292_),
    .A(_1289_),
    .B(_1291_));
 sg13g2_nor2b_1 _2172_ (.A(_1205_),
    .B_N(_1207_),
    .Y(_1293_));
 sg13g2_nand2_1 _2173_ (.Y(_1294_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_nand3_1 _2174_ (.B(\lfsr[1] ),
    .C(_1294_),
    .A(_1282_),
    .Y(_1295_));
 sg13g2_nand2_1 _2175_ (.Y(_1296_),
    .A(_1285_),
    .B(\lfsr[0] ));
 sg13g2_nand3_1 _2176_ (.B(_1296_),
    .C(_1249_),
    .A(_1295_),
    .Y(_1297_));
 sg13g2_nand2_1 _2177_ (.Y(_1298_),
    .A(_1282_),
    .B(_1294_));
 sg13g2_nand2_1 _2178_ (.Y(_1299_),
    .A(_1298_),
    .B(\lfsr[1] ));
 sg13g2_nand2_1 _2179_ (.Y(_1300_),
    .A(_1250_),
    .B(_1299_));
 sg13g2_nand2_1 _2180_ (.Y(_1301_),
    .A(_1297_),
    .B(_1300_));
 sg13g2_nand2_1 _2181_ (.Y(_1302_),
    .A(_1301_),
    .B(_1749_));
 sg13g2_nor2_1 _2182_ (.A(_1749_),
    .B(_1301_),
    .Y(_1303_));
 sg13g2_a21oi_1 _2183_ (.A1(_1302_),
    .A2(_1284_),
    .Y(_1304_),
    .B1(_1303_));
 sg13g2_nand2_1 _2184_ (.Y(_1305_),
    .A(_1280_),
    .B(\lfsr[3] ));
 sg13g2_nand2_1 _2185_ (.Y(_1306_),
    .A(_1304_),
    .B(_1305_));
 sg13g2_nand2_1 _2186_ (.Y(_1307_),
    .A(_1277_),
    .B(_1167_));
 sg13g2_nand3_1 _2187_ (.B(_1750_),
    .C(_1307_),
    .A(_1278_),
    .Y(_1308_));
 sg13g2_nand2_1 _2188_ (.Y(_1309_),
    .A(_1306_),
    .B(_1308_));
 sg13g2_nand2_1 _2189_ (.Y(_1310_),
    .A(_1288_),
    .B(_1309_));
 sg13g2_nand3_1 _2190_ (.B(_1279_),
    .C(_1308_),
    .A(_1306_),
    .Y(_1311_));
 sg13g2_buf_1 _2191_ (.A(_1311_),
    .X(_1312_));
 sg13g2_nand2_1 _2192_ (.Y(_1313_),
    .A(_1310_),
    .B(_1312_));
 sg13g2_xnor2_1 _2193_ (.Y(net18),
    .A(_1142_),
    .B(_1313_));
 sg13g2_xnor2_1 _2194_ (.Y(_1314_),
    .A(_1209_),
    .B(_1312_));
 sg13g2_nand2_1 _2195_ (.Y(_1315_),
    .A(_1313_),
    .B(_1141_));
 sg13g2_xnor2_1 _2196_ (.Y(net19),
    .A(_1314_),
    .B(_1315_));
 sg13g2_xnor2_1 _2197_ (.Y(_1316_),
    .A(_1275_),
    .B(_1209_));
 sg13g2_inv_1 _2198_ (.Y(_1317_),
    .A(_1316_));
 sg13g2_a21oi_1 _2199_ (.A1(_1310_),
    .A2(_1312_),
    .Y(_1318_),
    .B1(_1142_));
 sg13g2_nand2_1 _2200_ (.Y(_1319_),
    .A(_1318_),
    .B(_1314_));
 sg13g2_nand2b_1 _2201_ (.Y(_1320_),
    .B(_1312_),
    .A_N(_1209_));
 sg13g2_nand2_1 _2202_ (.Y(_1321_),
    .A(_1319_),
    .B(_1320_));
 sg13g2_xnor2_1 _2203_ (.Y(net20),
    .A(_1317_),
    .B(_1321_));
 sg13g2_nand2_1 _2204_ (.Y(_1322_),
    .A(_1209_),
    .B(_1271_));
 sg13g2_o21ai_1 _2205_ (.B1(_1322_),
    .Y(_1323_),
    .A1(_1317_),
    .A2(_1320_));
 sg13g2_xnor2_1 _2206_ (.Y(_1324_),
    .A(_1143_),
    .B(_1275_));
 sg13g2_nand4_1 _2207_ (.B(_1209_),
    .C(_1279_),
    .A(_1306_),
    .Y(_1325_),
    .D(_1308_));
 sg13g2_nand3_1 _2208_ (.B(_1325_),
    .C(_1316_),
    .A(_1320_),
    .Y(_1326_));
 sg13g2_nor2_1 _2209_ (.A(_1315_),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_nor3_1 _2210_ (.A(_1323_),
    .B(_1324_),
    .C(_1327_),
    .Y(_1328_));
 sg13g2_o21ai_1 _2211_ (.B1(_1081_),
    .Y(_1329_),
    .A1(net30),
    .A2(_1271_));
 sg13g2_nor2b_1 _2212_ (.A(_1328_),
    .B_N(_1329_),
    .Y(net21));
 sg13g2_buf_1 _2213_ (.A(\counter[21] ),
    .X(_1330_));
 sg13g2_buf_1 _2214_ (.A(\counter[20] ),
    .X(_1331_));
 sg13g2_buf_1 _2215_ (.A(\counter[23] ),
    .X(_1332_));
 sg13g2_buf_1 _2216_ (.A(\counter[22] ),
    .X(_1333_));
 sg13g2_nor4_1 _2217_ (.A(_1330_),
    .B(_1331_),
    .C(_1332_),
    .D(_1333_),
    .Y(_1334_));
 sg13g2_nor4_1 _2218_ (.A(\counter[17] ),
    .B(\counter[16] ),
    .C(\counter[19] ),
    .D(\counter[18] ),
    .Y(_1335_));
 sg13g2_buf_1 _2219_ (.A(\counter[25] ),
    .X(_1336_));
 sg13g2_buf_1 _2220_ (.A(\counter[24] ),
    .X(_1337_));
 sg13g2_buf_1 _2221_ (.A(\counter[26] ),
    .X(_1338_));
 sg13g2_nor3_1 _2222_ (.A(_1336_),
    .B(_1337_),
    .C(_1338_),
    .Y(_1339_));
 sg13g2_and3_1 _2223_ (.X(_1340_),
    .A(_1334_),
    .B(_1335_),
    .C(_1339_));
 sg13g2_nor4_1 _2224_ (.A(\counter[5] ),
    .B(\counter[4] ),
    .C(\counter[7] ),
    .D(\counter[6] ),
    .Y(_1341_));
 sg13g2_nor4_1 _2225_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .C(\counter[3] ),
    .D(\counter[2] ),
    .Y(_1342_));
 sg13g2_inv_1 _2226_ (.Y(_1343_),
    .A(\counter[9] ));
 sg13g2_inv_1 _2227_ (.Y(_1344_),
    .A(\counter[8] ));
 sg13g2_inv_1 _2228_ (.Y(_1345_),
    .A(\counter[11] ));
 sg13g2_inv_1 _2229_ (.Y(_1346_),
    .A(\counter[10] ));
 sg13g2_nand4_1 _2230_ (.B(_1344_),
    .C(_1345_),
    .A(_1343_),
    .Y(_1347_),
    .D(_1346_));
 sg13g2_nor4_1 _2231_ (.A(\counter[13] ),
    .B(\counter[12] ),
    .C(\counter[15] ),
    .D(\counter[14] ),
    .Y(_1348_));
 sg13g2_nor2b_1 _2232_ (.A(_1347_),
    .B_N(_1348_),
    .Y(_1349_));
 sg13g2_nand4_1 _2233_ (.B(_1341_),
    .C(_1342_),
    .A(_1340_),
    .Y(_0008_),
    .D(_1349_));
 sg13g2_buf_2 _2234_ (.A(\i_project.controller_0.rst_n ),
    .X(_1350_));
 sg13g2_buf_2 _2235_ (.A(\i_project.controller_0.divider[0] ),
    .X(_1351_));
 sg13g2_inv_1 _2236_ (.Y(_1352_),
    .A(_1351_));
 sg13g2_nor2_1 _2237_ (.A(_1350_),
    .B(\i_project.controller_0.grey_pass[10] ),
    .Y(_1353_));
 sg13g2_a21oi_1 _2238_ (.A1(_1350_),
    .A2(_1352_),
    .Y(_0003_),
    .B1(_1353_));
 sg13g2_buf_1 _2239_ (.A(_1350_),
    .X(_1354_));
 sg13g2_buf_1 _2240_ (.A(\i_project.controller_0.divider[1] ),
    .X(_1355_));
 sg13g2_inv_1 _2241_ (.Y(_1356_),
    .A(net76));
 sg13g2_nor2_1 _2242_ (.A(_1350_),
    .B(\i_project.controller_0.grey_pass[11] ),
    .Y(_1357_));
 sg13g2_a21oi_1 _2243_ (.A1(net66),
    .A2(net65),
    .Y(_0004_),
    .B1(_1357_));
 sg13g2_buf_1 _2244_ (.A(rst_n),
    .X(_1358_));
 sg13g2_inv_1 _2245_ (.Y(_1359_),
    .A(net77));
 sg13g2_buf_1 _2246_ (.A(_1359_),
    .X(_1360_));
 sg13g2_inv_1 _2247_ (.Y(_1361_),
    .A(_1336_));
 sg13g2_inv_1 _2248_ (.Y(_1362_),
    .A(\counter[7] ));
 sg13g2_inv_1 _2249_ (.Y(_1363_),
    .A(\counter[6] ));
 sg13g2_nand2_1 _2250_ (.Y(_1364_),
    .A(\counter[5] ),
    .B(\counter[4] ));
 sg13g2_nand2_1 _2251_ (.Y(_1365_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_nor2b_1 _2252_ (.A(_1365_),
    .B_N(\counter[2] ),
    .Y(_1366_));
 sg13g2_nand2_1 _2253_ (.Y(_1367_),
    .A(_1366_),
    .B(\counter[3] ));
 sg13g2_nor2_1 _2254_ (.A(_1364_),
    .B(_1367_),
    .Y(_1368_));
 sg13g2_inv_1 _2255_ (.Y(_1369_),
    .A(_1368_));
 sg13g2_nor3_1 _2256_ (.A(_1362_),
    .B(_1363_),
    .C(_1369_),
    .Y(_1370_));
 sg13g2_nand2_1 _2257_ (.Y(_1371_),
    .A(_1370_),
    .B(\counter[8] ));
 sg13g2_nor2_1 _2258_ (.A(_1343_),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_nand2_1 _2259_ (.Y(_1373_),
    .A(_1372_),
    .B(\counter[10] ));
 sg13g2_nor2_1 _2260_ (.A(_1345_),
    .B(_1373_),
    .Y(_1374_));
 sg13g2_nand2_1 _2261_ (.Y(_1375_),
    .A(_1374_),
    .B(\counter[12] ));
 sg13g2_nor2b_1 _2262_ (.A(_1375_),
    .B_N(\counter[13] ),
    .Y(_1376_));
 sg13g2_nand2_1 _2263_ (.Y(_1377_),
    .A(_1376_),
    .B(\counter[14] ));
 sg13g2_nor2b_1 _2264_ (.A(_1377_),
    .B_N(\counter[15] ),
    .Y(_1378_));
 sg13g2_nand2_1 _2265_ (.Y(_1379_),
    .A(_1378_),
    .B(\counter[16] ));
 sg13g2_nor2b_1 _2266_ (.A(_1379_),
    .B_N(\counter[17] ),
    .Y(_1380_));
 sg13g2_nand2_1 _2267_ (.Y(_1381_),
    .A(_1380_),
    .B(\counter[18] ));
 sg13g2_nor2b_1 _2268_ (.A(_1381_),
    .B_N(\counter[19] ),
    .Y(_1382_));
 sg13g2_buf_2 _2269_ (.A(_1382_),
    .X(_1383_));
 sg13g2_nand2_1 _2270_ (.Y(_1384_),
    .A(_1383_),
    .B(_1331_));
 sg13g2_nor2b_1 _2271_ (.A(_1384_),
    .B_N(_1330_),
    .Y(_1385_));
 sg13g2_nand2_1 _2272_ (.Y(_1386_),
    .A(_1385_),
    .B(_1333_));
 sg13g2_nor2b_1 _2273_ (.A(_1386_),
    .B_N(_1332_),
    .Y(_1387_));
 sg13g2_nand2_1 _2274_ (.Y(_1388_),
    .A(_1387_),
    .B(_1337_));
 sg13g2_nor2_1 _2275_ (.A(_1361_),
    .B(_1388_),
    .Y(_1389_));
 sg13g2_nand2_1 _2276_ (.Y(_1390_),
    .A(_1389_),
    .B(_1338_));
 sg13g2_nor2b_1 _2277_ (.A(_1390_),
    .B_N(\counter[27] ),
    .Y(_1391_));
 sg13g2_a21oi_1 _2278_ (.A1(_1391_),
    .A2(\counter[28] ),
    .Y(_1392_),
    .B1(\counter[29] ));
 sg13g2_nand3_1 _2279_ (.B(\counter[28] ),
    .C(\counter[29] ),
    .A(_1391_),
    .Y(_1393_));
 sg13g2_inv_1 _2280_ (.Y(_1394_),
    .A(_1393_));
 sg13g2_nor3_2 _2281_ (.A(net64),
    .B(_1392_),
    .C(_1394_),
    .Y(_0074_));
 sg13g2_inv_1 _2282_ (.Y(_1395_),
    .A(_1390_));
 sg13g2_nor2_1 _2283_ (.A(\counter[27] ),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_nor3_1 _2284_ (.A(_1359_),
    .B(_1391_),
    .C(_1396_),
    .Y(_0072_));
 sg13g2_inv_1 _2285_ (.Y(_1397_),
    .A(_0072_));
 sg13g2_inv_1 _2286_ (.Y(_1398_),
    .A(\counter[28] ));
 sg13g2_nand2_1 _2287_ (.Y(_1399_),
    .A(_1330_),
    .B(_1331_));
 sg13g2_nand4_1 _2288_ (.B(_1333_),
    .C(_1336_),
    .A(_1332_),
    .Y(_1400_),
    .D(_1337_));
 sg13g2_nand3b_1 _2289_ (.B(_1338_),
    .C(\counter[27] ),
    .Y(_1401_),
    .A_N(_1400_));
 sg13g2_nor2_1 _2290_ (.A(_1399_),
    .B(_1401_),
    .Y(_1402_));
 sg13g2_nand2_1 _2291_ (.Y(_1403_),
    .A(_1383_),
    .B(_1402_));
 sg13g2_nand4_1 _2292_ (.B(_1337_),
    .C(_1338_),
    .A(_1336_),
    .Y(_1404_),
    .D(\counter[27] ));
 sg13g2_nand4_1 _2293_ (.B(_1331_),
    .C(_1332_),
    .A(_1330_),
    .Y(_1405_),
    .D(_1333_));
 sg13g2_inv_1 _2294_ (.Y(_1406_),
    .A(_1383_));
 sg13g2_nor4_1 _2295_ (.A(_1398_),
    .B(_1404_),
    .C(_1405_),
    .D(_1406_),
    .Y(_1407_));
 sg13g2_nand2b_1 _2296_ (.Y(_1408_),
    .B(net77),
    .A_N(_1407_));
 sg13g2_a21oi_1 _2297_ (.A1(_1398_),
    .A2(_1403_),
    .Y(_0073_),
    .B1(_1408_));
 sg13g2_nand2_1 _2298_ (.Y(_1409_),
    .A(_1397_),
    .B(_0073_));
 sg13g2_nor2_1 _2299_ (.A(_0073_),
    .B(_1397_),
    .Y(_1410_));
 sg13g2_a21oi_1 _2300_ (.A1(_0074_),
    .A2(_1409_),
    .Y(_0000_),
    .B1(_1410_));
 sg13g2_inv_1 _2301_ (.Y(_1411_),
    .A(_0074_));
 sg13g2_o21ai_1 _2302_ (.B1(_1409_),
    .Y(_0001_),
    .A1(_1410_),
    .A2(_1411_));
 sg13g2_a21o_1 _2303_ (.A2(_0073_),
    .A1(_0074_),
    .B1(_0072_),
    .X(_0002_));
 sg13g2_buf_2 _2304_ (.A(ui_in[7]),
    .X(_1412_));
 sg13g2_mux2_1 _2305_ (.A0(_0012_),
    .A1(net1),
    .S(_1412_),
    .X(_0009_));
 sg13g2_mux2_1 _2306_ (.A0(_0013_),
    .A1(net2),
    .S(_1412_),
    .X(_0010_));
 sg13g2_mux2_1 _2307_ (.A0(_0014_),
    .A1(net3),
    .S(_1412_),
    .X(_0011_));
 sg13g2_mux2_1 _2308_ (.A0(_1337_),
    .A1(net5),
    .S(_1412_),
    .X(_0005_));
 sg13g2_nand2_1 _2309_ (.Y(_1413_),
    .A(_1412_),
    .B(net6));
 sg13g2_o21ai_1 _2310_ (.B1(_1413_),
    .Y(_0006_),
    .A1(_1412_),
    .A2(_1361_));
 sg13g2_mux2_1 _2311_ (.A0(_1338_),
    .A1(net7),
    .S(_1412_),
    .X(_0007_));
 sg13g2_buf_1 _2312_ (.A(\i_project.controller_0.h[1] ),
    .X(_1414_));
 sg13g2_buf_1 _2313_ (.A(_1414_),
    .X(_1415_));
 sg13g2_buf_1 _2314_ (.A(\i_project.controller_0.h[0] ),
    .X(_1416_));
 sg13g2_buf_1 _2315_ (.A(_1416_),
    .X(_1417_));
 sg13g2_nor2_1 _2316_ (.A(net63),
    .B(_1417_),
    .Y(_1418_));
 sg13g2_buf_1 _2317_ (.A(\i_project.controller_0.h[2] ),
    .X(_1419_));
 sg13g2_inv_1 _2318_ (.Y(_1420_),
    .A(_1419_));
 sg13g2_buf_1 _2319_ (.A(\i_project.controller_0.h[3] ),
    .X(_1421_));
 sg13g2_inv_2 _2320_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_nand3_1 _2321_ (.B(net61),
    .C(_1422_),
    .A(_1418_),
    .Y(_1423_));
 sg13g2_buf_1 _2322_ (.A(\i_project.controller_0.h[6] ),
    .X(_1424_));
 sg13g2_inv_2 _2323_ (.Y(_1425_),
    .A(net75));
 sg13g2_buf_1 _2324_ (.A(\i_project.controller_0.h[7] ),
    .X(_1426_));
 sg13g2_inv_1 _2325_ (.Y(_1427_),
    .A(net74));
 sg13g2_buf_2 _2326_ (.A(\i_project.controller_0.h[5] ),
    .X(_1428_));
 sg13g2_buf_1 _2327_ (.A(_1428_),
    .X(_1429_));
 sg13g2_buf_1 _2328_ (.A(\i_project.controller_0.h[4] ),
    .X(_1430_));
 sg13g2_buf_1 _2329_ (.A(_1430_),
    .X(_1431_));
 sg13g2_nand2_1 _2330_ (.Y(_1432_),
    .A(net60),
    .B(net59));
 sg13g2_nor3_1 _2331_ (.A(_1425_),
    .B(_1427_),
    .C(_1432_),
    .Y(_1433_));
 sg13g2_buf_2 _2332_ (.A(\i_project.controller_0.h[8] ),
    .X(_1434_));
 sg13g2_buf_1 _2333_ (.A(\i_project.controller_0.h[9] ),
    .X(_1435_));
 sg13g2_inv_1 _2334_ (.Y(_1436_),
    .A(_1435_));
 sg13g2_nor2_1 _2335_ (.A(_1434_),
    .B(_1436_),
    .Y(_1437_));
 sg13g2_nand3b_1 _2336_ (.B(_1433_),
    .C(_1437_),
    .Y(_1438_),
    .A_N(_1423_));
 sg13g2_nor2_1 _2337_ (.A(_1350_),
    .B(net77),
    .Y(_1439_));
 sg13g2_buf_2 _2338_ (.A(_1439_),
    .X(_1440_));
 sg13g2_inv_1 _2339_ (.Y(_1441_),
    .A(_1440_));
 sg13g2_nand3_1 _2340_ (.B(_0027_),
    .C(_1441_),
    .A(_1438_),
    .Y(_1442_));
 sg13g2_nand2_1 _2341_ (.Y(_1443_),
    .A(_1425_),
    .B(net74));
 sg13g2_inv_1 _2342_ (.Y(_1444_),
    .A(_1437_));
 sg13g2_inv_2 _2343_ (.Y(_1445_),
    .A(net59));
 sg13g2_nor2_1 _2344_ (.A(net60),
    .B(_1445_),
    .Y(_1446_));
 sg13g2_inv_1 _2345_ (.Y(_1447_),
    .A(_1446_));
 sg13g2_nor4_1 _2346_ (.A(_1443_),
    .B(_1444_),
    .C(_1447_),
    .D(_1423_),
    .Y(_1448_));
 sg13g2_nor3_1 _2347_ (.A(_1425_),
    .B(net74),
    .C(_1432_),
    .Y(_1449_));
 sg13g2_inv_1 _2348_ (.Y(_1450_),
    .A(_1449_));
 sg13g2_inv_1 _2349_ (.Y(_1451_),
    .A(_1434_));
 sg13g2_nor2_1 _2350_ (.A(_1435_),
    .B(_1451_),
    .Y(_1452_));
 sg13g2_buf_1 _2351_ (.A(_1419_),
    .X(_1453_));
 sg13g2_buf_1 _2352_ (.A(_1421_),
    .X(_1454_));
 sg13g2_nand4_1 _2353_ (.B(_1418_),
    .C(net58),
    .A(_1452_),
    .Y(_1455_),
    .D(_1454_));
 sg13g2_buf_2 _2354_ (.A(\i_project.controller_0.vga_sync.mode ),
    .X(_1456_));
 sg13g2_inv_2 _2355_ (.Y(_1457_),
    .A(_1456_));
 sg13g2_nand2_1 _2356_ (.Y(_1458_),
    .A(_1445_),
    .B(net60));
 sg13g2_inv_1 _2357_ (.Y(_1459_),
    .A(_1452_));
 sg13g2_inv_1 _2358_ (.Y(_1460_),
    .A(_1414_));
 sg13g2_nor2_1 _2359_ (.A(net62),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_nand3_1 _2360_ (.B(net61),
    .C(_1422_),
    .A(_1461_),
    .Y(_1462_));
 sg13g2_nor4_1 _2361_ (.A(_1458_),
    .B(_1459_),
    .C(_1443_),
    .D(_1462_),
    .Y(_1463_));
 sg13g2_nor3_1 _2362_ (.A(_1457_),
    .B(_1440_),
    .C(_1463_),
    .Y(_1464_));
 sg13g2_o21ai_1 _2363_ (.B1(_1464_),
    .Y(_1465_),
    .A1(_1450_),
    .A2(_1455_));
 sg13g2_o21ai_1 _2364_ (.B1(_1465_),
    .Y(_1466_),
    .A1(_1442_),
    .A2(_1448_));
 sg13g2_inv_1 _2365_ (.Y(_1467_),
    .A(\i_project.controller_0.vga_sync.hsync ));
 sg13g2_nor2b_1 _2366_ (.A(_1464_),
    .B_N(_1442_),
    .Y(_1468_));
 sg13g2_a21oi_1 _2367_ (.A1(_1466_),
    .A2(_1467_),
    .Y(_0111_),
    .B1(_1468_));
 sg13g2_buf_8 _2368_ (.A(\i_project.controller_0.v[4] ),
    .X(_1469_));
 sg13g2_buf_8 _2369_ (.A(\i_project.controller_0.v[5] ),
    .X(_1470_));
 sg13g2_inv_1 _2370_ (.Y(_1471_),
    .A(_1470_));
 sg13g2_buf_2 _2371_ (.A(\i_project.controller_0.v[7] ),
    .X(_1472_));
 sg13g2_inv_1 _2372_ (.Y(_1473_),
    .A(_1472_));
 sg13g2_buf_1 _2373_ (.A(\i_project.controller_0.v[6] ),
    .X(_1474_));
 sg13g2_inv_1 _2374_ (.Y(_1475_),
    .A(_1474_));
 sg13g2_nor4_1 _2375_ (.A(_1469_),
    .B(_1471_),
    .C(_1473_),
    .D(_1475_),
    .Y(_1476_));
 sg13g2_buf_2 _2376_ (.A(\i_project.controller_0.v[9] ),
    .X(_1477_));
 sg13g2_buf_2 _2377_ (.A(\i_project.controller_0.v[8] ),
    .X(_1478_));
 sg13g2_inv_1 _2378_ (.Y(_1479_),
    .A(_1478_));
 sg13g2_nor2_1 _2379_ (.A(_1477_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_and3_1 _2380_ (.X(_1481_),
    .A(_1476_),
    .B(_1457_),
    .C(_1480_));
 sg13g2_buf_8 _2381_ (.A(\i_project.controller_0.v[2] ),
    .X(_1482_));
 sg13g2_inv_1 _2382_ (.Y(_1483_),
    .A(_1482_));
 sg13g2_buf_8 _2383_ (.A(\i_project.controller_0.v[3] ),
    .X(_1484_));
 sg13g2_inv_4 _2384_ (.A(_1484_),
    .Y(_1485_));
 sg13g2_buf_1 _2385_ (.A(\i_project.controller_0.v[1] ),
    .X(_1486_));
 sg13g2_buf_8 _2386_ (.A(\i_project.controller_0.v[0] ),
    .X(_1487_));
 sg13g2_nor2_1 _2387_ (.A(net73),
    .B(_1487_),
    .Y(_1488_));
 sg13g2_inv_1 _2388_ (.Y(_1489_),
    .A(_1488_));
 sg13g2_nor3_1 _2389_ (.A(_1483_),
    .B(_1485_),
    .C(_1489_),
    .Y(_1490_));
 sg13g2_nand2_1 _2390_ (.Y(_1491_),
    .A(_1481_),
    .B(_1490_));
 sg13g2_nor3_1 _2391_ (.A(_1482_),
    .B(_1485_),
    .C(_1489_),
    .Y(_1492_));
 sg13g2_nor3_1 _2392_ (.A(_1469_),
    .B(_1470_),
    .C(_1474_),
    .Y(_1493_));
 sg13g2_inv_1 _2393_ (.Y(_1494_),
    .A(_1477_));
 sg13g2_nor3_1 _2394_ (.A(_1457_),
    .B(_1479_),
    .C(_1494_),
    .Y(_1495_));
 sg13g2_nand4_1 _2395_ (.B(_1472_),
    .C(_1493_),
    .A(_1492_),
    .Y(_1496_),
    .D(_1495_));
 sg13g2_nand3_1 _2396_ (.B(_1496_),
    .C(_1441_),
    .A(_1491_),
    .Y(_1497_));
 sg13g2_inv_1 _2397_ (.Y(_1498_),
    .A(_1493_));
 sg13g2_nor4_1 _2398_ (.A(_1483_),
    .B(_1484_),
    .C(_1473_),
    .D(_1498_),
    .Y(_1499_));
 sg13g2_inv_1 _2399_ (.Y(_1500_),
    .A(net73));
 sg13g2_and3_1 _2400_ (.X(_1501_),
    .A(_1495_),
    .B(_1500_),
    .C(_1487_));
 sg13g2_nor4_1 _2401_ (.A(_1487_),
    .B(_1482_),
    .C(_1500_),
    .D(_1485_),
    .Y(_1502_));
 sg13g2_a221oi_1 _2402_ (.B2(_1502_),
    .C1(\i_project.controller_0.vga_sync.vsync ),
    .B1(_1481_),
    .A1(_1499_),
    .Y(_1503_),
    .A2(_1501_));
 sg13g2_nor2_1 _2403_ (.A(_1497_),
    .B(_1503_),
    .Y(_0122_));
 sg13g2_inv_1 _2404_ (.Y(_1504_),
    .A(\i_project.controller_0.voffset[0] ));
 sg13g2_nor3_1 _2405_ (.A(_1425_),
    .B(net74),
    .C(_1459_),
    .Y(_1505_));
 sg13g2_inv_1 _2406_ (.Y(_1506_),
    .A(_1418_));
 sg13g2_nor4_1 _2407_ (.A(net58),
    .B(_1422_),
    .C(_1458_),
    .D(_1506_),
    .Y(_1507_));
 sg13g2_o21ai_1 _2408_ (.B1(_1434_),
    .Y(_1508_),
    .A1(net75),
    .A2(net74));
 sg13g2_buf_1 _2409_ (.A(_0025_),
    .X(_1509_));
 sg13g2_inv_1 _2410_ (.Y(_1510_),
    .A(_1509_));
 sg13g2_o21ai_1 _2411_ (.B1(net60),
    .Y(_1511_),
    .A1(_1431_),
    .A2(_1510_));
 sg13g2_a22oi_1 _2412_ (.Y(_1512_),
    .B1(_1511_),
    .B2(_1505_),
    .A2(_1508_),
    .A1(_1436_));
 sg13g2_a21o_1 _2413_ (.A2(_1507_),
    .A1(_1505_),
    .B1(_1512_),
    .X(_1513_));
 sg13g2_inv_1 _2414_ (.Y(_1514_),
    .A(_0028_));
 sg13g2_nor4_1 _2415_ (.A(net60),
    .B(_1431_),
    .C(_1443_),
    .D(_1423_),
    .Y(_1515_));
 sg13g2_nor3_1 _2416_ (.A(_1434_),
    .B(_1514_),
    .C(_1515_),
    .Y(_1516_));
 sg13g2_nor3_1 _2417_ (.A(_1456_),
    .B(_1436_),
    .C(_1516_),
    .Y(_1517_));
 sg13g2_a21oi_1 _2418_ (.A1(_1456_),
    .A2(_1513_),
    .Y(_1518_),
    .B1(_1517_));
 sg13g2_xor2_1 _2419_ (.B(\i_project.controller_0.grey_pass[14] ),
    .A(\i_project.controller_0.mode[2] ),
    .X(_1519_));
 sg13g2_buf_2 _2420_ (.A(\i_project.controller_0.mode[1] ),
    .X(_1520_));
 sg13g2_xor2_1 _2421_ (.B(\i_project.controller_0.grey_pass[13] ),
    .A(_1520_),
    .X(_1521_));
 sg13g2_nor2_1 _2422_ (.A(_1519_),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_buf_2 _2423_ (.A(\i_project.controller_0.mode[0] ),
    .X(_1523_));
 sg13g2_xnor2_1 _2424_ (.Y(_1524_),
    .A(_1523_),
    .B(\i_project.controller_0.grey_pass[12] ));
 sg13g2_inv_1 _2425_ (.Y(_1525_),
    .A(_0029_));
 sg13g2_nor3_2 _2426_ (.A(_1520_),
    .B(_1523_),
    .C(_1525_),
    .Y(_1526_));
 sg13g2_buf_1 _2427_ (.A(_1526_),
    .X(_1527_));
 sg13g2_a21oi_1 _2428_ (.A1(_1522_),
    .A2(_1524_),
    .Y(_1528_),
    .B1(_1527_));
 sg13g2_nand2b_1 _2429_ (.Y(_1529_),
    .B(_1528_),
    .A_N(_1518_));
 sg13g2_nand2_1 _2430_ (.Y(_1530_),
    .A(_1529_),
    .B(_1350_));
 sg13g2_buf_2 _2431_ (.A(_1530_),
    .X(_1531_));
 sg13g2_inv_1 _2432_ (.Y(_1532_),
    .A(_1531_));
 sg13g2_nand2b_1 _2433_ (.Y(_1533_),
    .B(net66),
    .A_N(_1524_));
 sg13g2_inv_1 _2434_ (.Y(_1534_),
    .A(\i_project.controller_0.mode[2] ));
 sg13g2_nor3_1 _2435_ (.A(_1520_),
    .B(_1350_),
    .C(_1534_),
    .Y(_1535_));
 sg13g2_nand2_1 _2436_ (.Y(_1536_),
    .A(_1535_),
    .B(_0016_));
 sg13g2_nor2b_2 _2437_ (.A(_1532_),
    .B_N(_1536_),
    .Y(_1537_));
 sg13g2_a22oi_1 _2438_ (.Y(_0123_),
    .B1(_1533_),
    .B2(_1537_),
    .A2(_1532_),
    .A1(_1504_));
 sg13g2_a22oi_1 _2439_ (.Y(_1538_),
    .B1(net66),
    .B2(_1521_),
    .A2(_0015_),
    .A1(_1535_));
 sg13g2_buf_2 _2440_ (.A(\i_project.controller_0.voffset[1] ),
    .X(_1539_));
 sg13g2_nor2_1 _2441_ (.A(_1539_),
    .B(_1531_),
    .Y(_1540_));
 sg13g2_a21oi_1 _2442_ (.A1(_1531_),
    .A2(_1538_),
    .Y(_0124_),
    .B1(_1540_));
 sg13g2_inv_1 _2443_ (.Y(_1541_),
    .A(\i_project.controller_0.voffset[2] ));
 sg13g2_nand2_1 _2444_ (.Y(_1542_),
    .A(_1519_),
    .B(net66));
 sg13g2_a22oi_1 _2445_ (.Y(_0125_),
    .B1(_1542_),
    .B2(_1537_),
    .A2(_1532_),
    .A1(_1541_));
 sg13g2_inv_1 _2446_ (.Y(_1543_),
    .A(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_1 _2447_ (.Y(_1544_),
    .A(_1535_),
    .B(_0164_));
 sg13g2_o21ai_1 _2448_ (.B1(_1544_),
    .Y(_0126_),
    .A1(_1543_),
    .A2(_1531_));
 sg13g2_inv_1 _2449_ (.Y(_1545_),
    .A(\i_project.controller_0.voffset[4] ));
 sg13g2_o21ai_1 _2450_ (.B1(_1536_),
    .Y(_0127_),
    .A1(_1545_),
    .A2(_1531_));
 sg13g2_inv_1 _2451_ (.Y(_1546_),
    .A(\i_project.controller_0.voffset[5] ));
 sg13g2_buf_1 _2452_ (.A(_1350_),
    .X(_1547_));
 sg13g2_nand2_1 _2453_ (.Y(_1548_),
    .A(net56),
    .B(\i_project.controller_0.grey_pass[10] ));
 sg13g2_a22oi_1 _2454_ (.Y(_0128_),
    .B1(_1548_),
    .B2(_1537_),
    .A2(_1532_),
    .A1(_1546_));
 sg13g2_inv_1 _2455_ (.Y(_1549_),
    .A(\i_project.controller_0.voffset[6] ));
 sg13g2_nand2_1 _2456_ (.Y(_1550_),
    .A(net56),
    .B(\i_project.controller_0.grey_pass[11] ));
 sg13g2_a22oi_1 _2457_ (.Y(_0129_),
    .B1(_1550_),
    .B2(_1537_),
    .A2(_1532_),
    .A1(_1549_));
 sg13g2_inv_1 _2458_ (.Y(_1551_),
    .A(\i_project.controller_0.voffset[7] ));
 sg13g2_nand3_1 _2459_ (.B(_1354_),
    .C(\i_project.controller_0.grey_pass[15] ),
    .A(_1531_),
    .Y(_1552_));
 sg13g2_o21ai_1 _2460_ (.B1(_1552_),
    .Y(_0130_),
    .A1(_1551_),
    .A2(_1531_));
 sg13g2_inv_1 _2461_ (.Y(_1553_),
    .A(_1523_));
 sg13g2_nor2_1 _2462_ (.A(net56),
    .B(\i_project.controller_0.grey_pass[12] ),
    .Y(_1554_));
 sg13g2_a21oi_1 _2463_ (.A1(_1553_),
    .A2(net56),
    .Y(_0085_),
    .B1(_1554_));
 sg13g2_inv_1 _2464_ (.Y(_1555_),
    .A(_1520_));
 sg13g2_nor2_1 _2465_ (.A(net56),
    .B(\i_project.controller_0.grey_pass[13] ),
    .Y(_1556_));
 sg13g2_a21oi_1 _2466_ (.A1(_1555_),
    .A2(net56),
    .Y(_0086_),
    .B1(_1556_));
 sg13g2_nor2_1 _2467_ (.A(_1547_),
    .B(\i_project.controller_0.grey_pass[14] ),
    .Y(_1557_));
 sg13g2_a21oi_1 _2468_ (.A1(_1534_),
    .A2(_1547_),
    .Y(_0087_),
    .B1(_1557_));
 sg13g2_nor2_1 _2469_ (.A(net66),
    .B(\i_project.controller_0.grey_pass[15] ),
    .Y(_1558_));
 sg13g2_a21oi_1 _2470_ (.A1(_1457_),
    .A2(net56),
    .Y(_0088_),
    .B1(_1558_));
 sg13g2_inv_1 _2471_ (.Y(_1559_),
    .A(_0049_));
 sg13g2_nor4_1 _2472_ (.A(_1435_),
    .B(_1457_),
    .C(_1425_),
    .D(_1427_),
    .Y(_1560_));
 sg13g2_nor2_1 _2473_ (.A(_1453_),
    .B(_1560_),
    .Y(_1561_));
 sg13g2_nand2_2 _2474_ (.Y(_1562_),
    .A(net63),
    .B(net62));
 sg13g2_nand4_1 _2475_ (.B(_1425_),
    .C(_1427_),
    .A(_1457_),
    .Y(_1563_),
    .D(_1435_));
 sg13g2_nand2_1 _2476_ (.Y(_1564_),
    .A(_1563_),
    .B(net58));
 sg13g2_inv_1 _2477_ (.Y(_1565_),
    .A(_0026_));
 sg13g2_nand3_1 _2478_ (.B(_1565_),
    .C(_1446_),
    .A(_1564_),
    .Y(_1566_));
 sg13g2_nor4_2 _2479_ (.A(_1509_),
    .B(_1561_),
    .C(_1562_),
    .Y(_1567_),
    .D(_1566_));
 sg13g2_nor2_1 _2480_ (.A(_1440_),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_inv_1 _2481_ (.Y(_1569_),
    .A(_1568_));
 sg13g2_nor2_1 _2482_ (.A(_1559_),
    .B(net31),
    .Y(_0101_));
 sg13g2_inv_1 _2483_ (.Y(_1570_),
    .A(_1562_));
 sg13g2_nor3_1 _2484_ (.A(_1418_),
    .B(_1570_),
    .C(net31),
    .Y(_0102_));
 sg13g2_nor2_1 _2485_ (.A(_1453_),
    .B(_1570_),
    .Y(_1571_));
 sg13g2_nor2_1 _2486_ (.A(net61),
    .B(_1562_),
    .Y(_1572_));
 sg13g2_nor3_1 _2487_ (.A(_1571_),
    .B(_1572_),
    .C(_1569_),
    .Y(_0103_));
 sg13g2_nor2_1 _2488_ (.A(_1454_),
    .B(_1572_),
    .Y(_1573_));
 sg13g2_nor3_1 _2489_ (.A(net61),
    .B(_1422_),
    .C(_1562_),
    .Y(_1574_));
 sg13g2_nor3_1 _2490_ (.A(_1573_),
    .B(_1574_),
    .C(net31),
    .Y(_0104_));
 sg13g2_nor2_1 _2491_ (.A(net59),
    .B(_1574_),
    .Y(_1575_));
 sg13g2_nand2_1 _2492_ (.Y(_1576_),
    .A(_1574_),
    .B(net59));
 sg13g2_inv_1 _2493_ (.Y(_1577_),
    .A(_1576_));
 sg13g2_nor3_1 _2494_ (.A(_1575_),
    .B(_1577_),
    .C(_1569_),
    .Y(_0105_));
 sg13g2_nor2_1 _2495_ (.A(_1429_),
    .B(_1577_),
    .Y(_1578_));
 sg13g2_inv_1 _2496_ (.Y(_1579_),
    .A(_1428_));
 sg13g2_nor2_1 _2497_ (.A(_1579_),
    .B(_1576_),
    .Y(_1580_));
 sg13g2_nor3_1 _2498_ (.A(_1578_),
    .B(_1580_),
    .C(net31),
    .Y(_0106_));
 sg13g2_nor2_1 _2499_ (.A(_1424_),
    .B(_1580_),
    .Y(_1581_));
 sg13g2_nand2_1 _2500_ (.Y(_1582_),
    .A(_1580_),
    .B(_1424_));
 sg13g2_inv_1 _2501_ (.Y(_1583_),
    .A(_1582_));
 sg13g2_nor3_1 _2502_ (.A(_1581_),
    .B(_1583_),
    .C(net31),
    .Y(_0107_));
 sg13g2_nand2_1 _2503_ (.Y(_1584_),
    .A(_1583_),
    .B(_1427_));
 sg13g2_nand2_1 _2504_ (.Y(_1585_),
    .A(_1582_),
    .B(net74));
 sg13g2_a21oi_1 _2505_ (.A1(_1584_),
    .A2(_1585_),
    .Y(_0108_),
    .B1(net31));
 sg13g2_a21oi_1 _2506_ (.A1(_1583_),
    .A2(_1426_),
    .Y(_1586_),
    .B1(_1434_));
 sg13g2_nor3_1 _2507_ (.A(_1427_),
    .B(_1451_),
    .C(_1582_),
    .Y(_1587_));
 sg13g2_nor3_1 _2508_ (.A(_1586_),
    .B(_1587_),
    .C(net31),
    .Y(_0109_));
 sg13g2_xnor2_1 _2509_ (.Y(_1588_),
    .A(_1435_),
    .B(_1587_));
 sg13g2_nor2_1 _2510_ (.A(_1588_),
    .B(net31),
    .Y(_0110_));
 sg13g2_inv_1 _2511_ (.Y(_1589_),
    .A(_1487_));
 sg13g2_nor4_1 _2512_ (.A(_1509_),
    .B(_0026_),
    .C(_1562_),
    .D(_1447_),
    .Y(_1590_));
 sg13g2_nand3b_1 _2513_ (.B(_1564_),
    .C(_1590_),
    .Y(_1591_),
    .A_N(_1561_));
 sg13g2_buf_1 _2514_ (.A(_1591_),
    .X(_1592_));
 sg13g2_nor2_1 _2515_ (.A(_1589_),
    .B(_1592_),
    .Y(_1593_));
 sg13g2_nor4_1 _2516_ (.A(_1456_),
    .B(_1472_),
    .C(_1478_),
    .D(_1498_),
    .Y(_1594_));
 sg13g2_nand2_1 _2517_ (.Y(_1595_),
    .A(net73),
    .B(_1487_));
 sg13g2_nand2_1 _2518_ (.Y(_1596_),
    .A(_1472_),
    .B(_1478_));
 sg13g2_inv_1 _2519_ (.Y(_1597_),
    .A(_1596_));
 sg13g2_nor2_1 _2520_ (.A(_1482_),
    .B(_1484_),
    .Y(_1598_));
 sg13g2_nand4_1 _2521_ (.B(_1598_),
    .C(_1456_),
    .A(_1597_),
    .Y(_1599_),
    .D(_1475_));
 sg13g2_nor4_1 _2522_ (.A(_1469_),
    .B(_1471_),
    .C(_1595_),
    .D(_1599_),
    .Y(_1600_));
 sg13g2_a21o_1 _2523_ (.A2(_1594_),
    .A1(_1490_),
    .B1(_1600_),
    .X(_1601_));
 sg13g2_inv_1 _2524_ (.Y(_1602_),
    .A(_0030_));
 sg13g2_nand2_2 _2525_ (.Y(_1603_),
    .A(_1601_),
    .B(_1602_));
 sg13g2_a21oi_1 _2526_ (.A1(_1603_),
    .A2(_1567_),
    .Y(_1604_),
    .B1(_1487_));
 sg13g2_nor3_1 _2527_ (.A(_1440_),
    .B(_1593_),
    .C(_1604_),
    .Y(_0112_));
 sg13g2_nor2_1 _2528_ (.A(net73),
    .B(_1593_),
    .Y(_1605_));
 sg13g2_nand2_1 _2529_ (.Y(_1606_),
    .A(_1593_),
    .B(net73));
 sg13g2_inv_1 _2530_ (.Y(_1607_),
    .A(_1606_));
 sg13g2_nor3_1 _2531_ (.A(_1440_),
    .B(_1605_),
    .C(_1607_),
    .Y(_0113_));
 sg13g2_nor2_1 _2532_ (.A(_1483_),
    .B(_1606_),
    .Y(_1608_));
 sg13g2_nor2_1 _2533_ (.A(_1482_),
    .B(_1607_),
    .Y(_1609_));
 sg13g2_inv_1 _2534_ (.Y(_1610_),
    .A(_1603_));
 sg13g2_nand2_1 _2535_ (.Y(_1611_),
    .A(_1610_),
    .B(_1567_));
 sg13g2_nand2_1 _2536_ (.Y(_1612_),
    .A(_1611_),
    .B(_1441_));
 sg13g2_nor3_1 _2537_ (.A(_1608_),
    .B(_1609_),
    .C(_1612_),
    .Y(_0114_));
 sg13g2_nor2_1 _2538_ (.A(_1484_),
    .B(_1608_),
    .Y(_1613_));
 sg13g2_nor2_1 _2539_ (.A(_1483_),
    .B(_1595_),
    .Y(_1614_));
 sg13g2_nand2_1 _2540_ (.Y(_1615_),
    .A(_1614_),
    .B(_1484_));
 sg13g2_inv_1 _2541_ (.Y(_1616_),
    .A(_1615_));
 sg13g2_nand2_1 _2542_ (.Y(_1617_),
    .A(_1567_),
    .B(_1616_));
 sg13g2_inv_1 _2543_ (.Y(_1618_),
    .A(_1617_));
 sg13g2_nor3_1 _2544_ (.A(_1613_),
    .B(_1618_),
    .C(_1612_),
    .Y(_0115_));
 sg13g2_inv_1 _2545_ (.Y(_1619_),
    .A(_1469_));
 sg13g2_xnor2_1 _2546_ (.Y(_1620_),
    .A(_1619_),
    .B(_1617_));
 sg13g2_nor2_1 _2547_ (.A(_1440_),
    .B(_1620_),
    .Y(_0116_));
 sg13g2_nor2_1 _2548_ (.A(_1619_),
    .B(_1615_),
    .Y(_1621_));
 sg13g2_xor2_1 _2549_ (.B(_1621_),
    .A(_0031_),
    .X(_1622_));
 sg13g2_nand3b_1 _2550_ (.B(_1603_),
    .C(_1441_),
    .Y(_1623_),
    .A_N(_1592_));
 sg13g2_nand2_1 _2551_ (.Y(_1624_),
    .A(_1568_),
    .B(_1470_));
 sg13g2_o21ai_1 _2552_ (.B1(_1624_),
    .Y(_0117_),
    .A1(_1622_),
    .A2(_1623_));
 sg13g2_nor3_1 _2553_ (.A(_1619_),
    .B(_1471_),
    .C(_1617_),
    .Y(_1625_));
 sg13g2_xnor2_1 _2554_ (.Y(_1626_),
    .A(_1474_),
    .B(_1625_));
 sg13g2_nor2_1 _2555_ (.A(_1440_),
    .B(_1626_),
    .Y(_0118_));
 sg13g2_nor4_2 _2556_ (.A(_1619_),
    .B(_1471_),
    .C(_1475_),
    .Y(_1627_),
    .D(_1615_));
 sg13g2_a21oi_1 _2557_ (.A1(_1567_),
    .A2(_1627_),
    .Y(_1628_),
    .B1(_1472_));
 sg13g2_nand2_1 _2558_ (.Y(_1629_),
    .A(_1627_),
    .B(_1472_));
 sg13g2_nor2_1 _2559_ (.A(_1629_),
    .B(_1592_),
    .Y(_1630_));
 sg13g2_nor3_1 _2560_ (.A(_1628_),
    .B(_1630_),
    .C(_1612_),
    .Y(_0119_));
 sg13g2_xnor2_1 _2561_ (.Y(_1631_),
    .A(_0032_),
    .B(_1629_));
 sg13g2_nand2_1 _2562_ (.Y(_1632_),
    .A(_1568_),
    .B(_1478_));
 sg13g2_o21ai_1 _2563_ (.B1(_1632_),
    .Y(_0120_),
    .A1(_1631_),
    .A2(_1623_));
 sg13g2_nand2_1 _2564_ (.Y(_1633_),
    .A(_1627_),
    .B(_1597_));
 sg13g2_xnor2_1 _2565_ (.Y(_1634_),
    .A(_0030_),
    .B(_1633_));
 sg13g2_nand2_1 _2566_ (.Y(_1635_),
    .A(_1568_),
    .B(_1477_));
 sg13g2_o21ai_1 _2567_ (.B1(_1635_),
    .Y(_0121_),
    .A1(_1634_),
    .A2(_1623_));
 sg13g2_and2_1 _2568_ (.A(_0004_),
    .B(_0003_),
    .X(_0052_));
 sg13g2_nand2_1 _2569_ (.Y(_1636_),
    .A(_1358_),
    .B(_0050_));
 sg13g2_inv_1 _2570_ (.Y(_0053_),
    .A(_1636_));
 sg13g2_buf_1 _2571_ (.A(net64),
    .X(_1637_));
 sg13g2_nor2_1 _2572_ (.A(\counter[10] ),
    .B(_1372_),
    .Y(_1638_));
 sg13g2_inv_1 _2573_ (.Y(_1639_),
    .A(_1373_));
 sg13g2_nor3_1 _2574_ (.A(net51),
    .B(_1638_),
    .C(_1639_),
    .Y(_0054_));
 sg13g2_nor2_1 _2575_ (.A(\counter[11] ),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_nor3_1 _2576_ (.A(net51),
    .B(_1374_),
    .C(_1640_),
    .Y(_0055_));
 sg13g2_nor2_1 _2577_ (.A(\counter[12] ),
    .B(_1374_),
    .Y(_1641_));
 sg13g2_inv_1 _2578_ (.Y(_1642_),
    .A(_1375_));
 sg13g2_nor3_1 _2579_ (.A(net51),
    .B(_1641_),
    .C(_1642_),
    .Y(_0056_));
 sg13g2_nor2_1 _2580_ (.A(\counter[13] ),
    .B(_1642_),
    .Y(_1643_));
 sg13g2_nor3_1 _2581_ (.A(net51),
    .B(_1376_),
    .C(_1643_),
    .Y(_0057_));
 sg13g2_nor2_1 _2582_ (.A(\counter[14] ),
    .B(_1376_),
    .Y(_1644_));
 sg13g2_inv_1 _2583_ (.Y(_1645_),
    .A(_1377_));
 sg13g2_nor3_1 _2584_ (.A(_1637_),
    .B(_1644_),
    .C(_1645_),
    .Y(_0058_));
 sg13g2_nor2_1 _2585_ (.A(\counter[15] ),
    .B(_1645_),
    .Y(_1646_));
 sg13g2_nor3_1 _2586_ (.A(net51),
    .B(_1378_),
    .C(_1646_),
    .Y(_0059_));
 sg13g2_nor2_1 _2587_ (.A(\counter[16] ),
    .B(_1378_),
    .Y(_1647_));
 sg13g2_inv_1 _2588_ (.Y(_1648_),
    .A(_1379_));
 sg13g2_nor3_1 _2589_ (.A(net51),
    .B(_1647_),
    .C(_1648_),
    .Y(_0060_));
 sg13g2_nor2_1 _2590_ (.A(\counter[17] ),
    .B(_1648_),
    .Y(_1649_));
 sg13g2_nor3_1 _2591_ (.A(net51),
    .B(_1380_),
    .C(_1649_),
    .Y(_0061_));
 sg13g2_nor2_1 _2592_ (.A(\counter[18] ),
    .B(_1380_),
    .Y(_1650_));
 sg13g2_inv_1 _2593_ (.Y(_1651_),
    .A(_1381_));
 sg13g2_nor3_1 _2594_ (.A(net51),
    .B(_1650_),
    .C(_1651_),
    .Y(_0062_));
 sg13g2_nor2_1 _2595_ (.A(\counter[19] ),
    .B(_1651_),
    .Y(_1652_));
 sg13g2_nor3_1 _2596_ (.A(_1637_),
    .B(_1383_),
    .C(_1652_),
    .Y(_0063_));
 sg13g2_buf_1 _2597_ (.A(net64),
    .X(_1653_));
 sg13g2_nor2_1 _2598_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_1654_));
 sg13g2_inv_1 _2599_ (.Y(_1655_),
    .A(_1365_));
 sg13g2_nor3_1 _2600_ (.A(net50),
    .B(_1654_),
    .C(_1655_),
    .Y(_0064_));
 sg13g2_nor2_1 _2601_ (.A(_1331_),
    .B(_1383_),
    .Y(_1656_));
 sg13g2_inv_1 _2602_ (.Y(_1657_),
    .A(_1384_));
 sg13g2_nor3_1 _2603_ (.A(net50),
    .B(_1656_),
    .C(_1657_),
    .Y(_0065_));
 sg13g2_nor2_1 _2604_ (.A(_1330_),
    .B(_1657_),
    .Y(_1658_));
 sg13g2_nor3_1 _2605_ (.A(net50),
    .B(_1385_),
    .C(_1658_),
    .Y(_0066_));
 sg13g2_nor2_1 _2606_ (.A(_1333_),
    .B(_1385_),
    .Y(_1659_));
 sg13g2_inv_1 _2607_ (.Y(_1660_),
    .A(_1386_));
 sg13g2_nor3_1 _2608_ (.A(_1653_),
    .B(_1659_),
    .C(_1660_),
    .Y(_0067_));
 sg13g2_nor2_1 _2609_ (.A(_1332_),
    .B(_1660_),
    .Y(_1661_));
 sg13g2_nor3_1 _2610_ (.A(_1653_),
    .B(_1387_),
    .C(_1661_),
    .Y(_0068_));
 sg13g2_nor2_1 _2611_ (.A(_1337_),
    .B(_1387_),
    .Y(_1662_));
 sg13g2_inv_1 _2612_ (.Y(_1663_),
    .A(_1388_));
 sg13g2_nor3_1 _2613_ (.A(net50),
    .B(_1662_),
    .C(_1663_),
    .Y(_0069_));
 sg13g2_nor2_1 _2614_ (.A(_1336_),
    .B(_1663_),
    .Y(_1664_));
 sg13g2_nor3_1 _2615_ (.A(net50),
    .B(_1389_),
    .C(_1664_),
    .Y(_0070_));
 sg13g2_nor2_1 _2616_ (.A(_1338_),
    .B(_1389_),
    .Y(_1665_));
 sg13g2_nor3_1 _2617_ (.A(net50),
    .B(_1665_),
    .C(_1395_),
    .Y(_0071_));
 sg13g2_nor2_1 _2618_ (.A(\counter[2] ),
    .B(_1655_),
    .Y(_1666_));
 sg13g2_nor3_1 _2619_ (.A(net50),
    .B(_1366_),
    .C(_1666_),
    .Y(_0075_));
 sg13g2_inv_1 _2620_ (.Y(_1667_),
    .A(\counter[30] ));
 sg13g2_nand2_1 _2621_ (.Y(_1668_),
    .A(_1394_),
    .B(\counter[30] ));
 sg13g2_nand2_1 _2622_ (.Y(_1669_),
    .A(_1668_),
    .B(_1358_));
 sg13g2_a21oi_1 _2623_ (.A1(_1667_),
    .A2(_1393_),
    .Y(_0076_),
    .B1(_1669_));
 sg13g2_inv_1 _2624_ (.Y(_1670_),
    .A(\counter[31] ));
 sg13g2_o21ai_1 _2625_ (.B1(net77),
    .Y(_1671_),
    .A1(_1670_),
    .A2(_1668_));
 sg13g2_a21oi_1 _2626_ (.A1(_1670_),
    .A2(_1668_),
    .Y(_0077_),
    .B1(_1671_));
 sg13g2_nor2_1 _2627_ (.A(\counter[3] ),
    .B(_1366_),
    .Y(_1672_));
 sg13g2_inv_1 _2628_ (.Y(_1673_),
    .A(_1367_));
 sg13g2_nor3_1 _2629_ (.A(net50),
    .B(_1672_),
    .C(_1673_),
    .Y(_0078_));
 sg13g2_nor2b_1 _2630_ (.A(_1367_),
    .B_N(\counter[4] ),
    .Y(_1674_));
 sg13g2_nor2_1 _2631_ (.A(\counter[4] ),
    .B(_1673_),
    .Y(_1675_));
 sg13g2_nor3_1 _2632_ (.A(net64),
    .B(_1674_),
    .C(_1675_),
    .Y(_0079_));
 sg13g2_nor2_1 _2633_ (.A(\counter[5] ),
    .B(_1674_),
    .Y(_1676_));
 sg13g2_nor3_1 _2634_ (.A(net64),
    .B(_1368_),
    .C(_1676_),
    .Y(_0080_));
 sg13g2_nor2_1 _2635_ (.A(\counter[6] ),
    .B(_1368_),
    .Y(_1677_));
 sg13g2_nor2_1 _2636_ (.A(_1363_),
    .B(_1369_),
    .Y(_1678_));
 sg13g2_nor3_1 _2637_ (.A(net64),
    .B(_1677_),
    .C(_1678_),
    .Y(_0081_));
 sg13g2_nor2_1 _2638_ (.A(\counter[7] ),
    .B(_1678_),
    .Y(_1679_));
 sg13g2_nor3_1 _2639_ (.A(net64),
    .B(_1370_),
    .C(_1679_),
    .Y(_0082_));
 sg13g2_nor2_1 _2640_ (.A(\counter[8] ),
    .B(_1370_),
    .Y(_1680_));
 sg13g2_inv_1 _2641_ (.Y(_1681_),
    .A(_1371_));
 sg13g2_nor3_1 _2642_ (.A(net64),
    .B(_1680_),
    .C(_1681_),
    .Y(_0083_));
 sg13g2_nor2_1 _2643_ (.A(\counter[9] ),
    .B(_1681_),
    .Y(_1682_));
 sg13g2_nor3_1 _2644_ (.A(_1360_),
    .B(_1372_),
    .C(_1682_),
    .Y(_0084_));
 sg13g2_inv_1 _2645_ (.Y(_1683_),
    .A(_0051_));
 sg13g2_nor2_2 _2646_ (.A(_1592_),
    .B(_1603_),
    .Y(_1684_));
 sg13g2_buf_2 _2647_ (.A(\i_project.controller_0.mode_ramp_base[0] ),
    .X(_1685_));
 sg13g2_o21ai_1 _2648_ (.B1(net66),
    .Y(_1686_),
    .A1(_1685_),
    .A2(_1684_));
 sg13g2_a21oi_1 _2649_ (.A1(_1683_),
    .A2(_1684_),
    .Y(_0089_),
    .B1(_1686_));
 sg13g2_buf_1 _2650_ (.A(\i_project.controller_0.t[9] ),
    .X(_1687_));
 sg13g2_inv_1 _2651_ (.Y(_1688_),
    .A(_1687_));
 sg13g2_buf_1 _2652_ (.A(\i_project.controller_0.mode_ramp_base[5] ),
    .X(_1689_));
 sg13g2_inv_1 _2653_ (.Y(_1690_),
    .A(net72));
 sg13g2_buf_1 _2654_ (.A(\i_project.controller_0.mode_ramp_base[6] ),
    .X(_1691_));
 sg13g2_inv_2 _2655_ (.Y(_1692_),
    .A(net71));
 sg13g2_buf_2 _2656_ (.A(\i_project.controller_0.mode_ramp_base[7] ),
    .X(_1693_));
 sg13g2_inv_1 _2657_ (.Y(_1694_),
    .A(_1693_));
 sg13g2_buf_1 _2658_ (.A(\i_project.controller_0.mode_ramp_base[3] ),
    .X(_1695_));
 sg13g2_buf_1 _2659_ (.A(_1695_),
    .X(_1696_));
 sg13g2_buf_1 _2660_ (.A(\i_project.controller_0.mode_ramp_base[4] ),
    .X(_1697_));
 sg13g2_buf_1 _2661_ (.A(_1697_),
    .X(_1698_));
 sg13g2_nand2_1 _2662_ (.Y(_1699_),
    .A(net55),
    .B(net54));
 sg13g2_buf_1 _2663_ (.A(\i_project.controller_0.mode_ramp_base[2] ),
    .X(_1700_));
 sg13g2_buf_2 _2664_ (.A(\i_project.controller_0.mode_ramp_base[1] ),
    .X(_1701_));
 sg13g2_nand2_1 _2665_ (.Y(_1702_),
    .A(_1701_),
    .B(_1685_));
 sg13g2_inv_1 _2666_ (.Y(_1703_),
    .A(_1702_));
 sg13g2_nand3_1 _2667_ (.B(net70),
    .C(_1703_),
    .A(_1684_),
    .Y(_1704_));
 sg13g2_buf_1 _2668_ (.A(_1704_),
    .X(_1705_));
 sg13g2_nor2_1 _2669_ (.A(_1699_),
    .B(_1705_),
    .Y(_1706_));
 sg13g2_inv_1 _2670_ (.Y(_1707_),
    .A(_1706_));
 sg13g2_nor4_1 _2671_ (.A(_1690_),
    .B(_1692_),
    .C(_1694_),
    .D(_1707_),
    .Y(_1708_));
 sg13g2_buf_8 _2672_ (.A(\i_project.controller_0.t[8] ),
    .X(_1709_));
 sg13g2_nand2_1 _2673_ (.Y(_1710_),
    .A(_1708_),
    .B(_1709_));
 sg13g2_nor2_1 _2674_ (.A(_1688_),
    .B(_1710_),
    .Y(_1711_));
 sg13g2_nor2_1 _2675_ (.A(\i_project.controller_0.t[10] ),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_nand2_1 _2676_ (.Y(_1713_),
    .A(_1711_),
    .B(\i_project.controller_0.t[10] ));
 sg13g2_nand2_1 _2677_ (.Y(_1714_),
    .A(_1713_),
    .B(net56));
 sg13g2_nor2_1 _2678_ (.A(_1712_),
    .B(_1714_),
    .Y(_0090_));
 sg13g2_inv_1 _2679_ (.Y(_1715_),
    .A(\i_project.controller_0.t[11] ));
 sg13g2_o21ai_1 _2680_ (.B1(_1354_),
    .Y(_1716_),
    .A1(_1715_),
    .A2(_1713_));
 sg13g2_a21oi_1 _2681_ (.A1(_1715_),
    .A2(_1713_),
    .Y(_0091_),
    .B1(_1716_));
 sg13g2_inv_2 _2682_ (.Y(_1717_),
    .A(net66));
 sg13g2_a21oi_1 _2683_ (.A1(_1684_),
    .A2(_1685_),
    .Y(_1718_),
    .B1(_1701_));
 sg13g2_inv_1 _2684_ (.Y(_1719_),
    .A(_1701_));
 sg13g2_inv_1 _2685_ (.Y(_1720_),
    .A(_1685_));
 sg13g2_nor3_1 _2686_ (.A(_1719_),
    .B(_1720_),
    .C(_1611_),
    .Y(_1721_));
 sg13g2_nor3_1 _2687_ (.A(_1717_),
    .B(_1718_),
    .C(_1721_),
    .Y(_0092_));
 sg13g2_inv_1 _2688_ (.Y(_1722_),
    .A(_1705_));
 sg13g2_nor2_1 _2689_ (.A(net70),
    .B(_1721_),
    .Y(_1723_));
 sg13g2_nor3_1 _2690_ (.A(_1717_),
    .B(_1722_),
    .C(_1723_),
    .Y(_0093_));
 sg13g2_inv_1 _2691_ (.Y(_1724_),
    .A(_1695_));
 sg13g2_o21ai_1 _2692_ (.B1(net66),
    .Y(_1725_),
    .A1(_1724_),
    .A2(_1705_));
 sg13g2_a21oi_1 _2693_ (.A1(_1724_),
    .A2(_1705_),
    .Y(_0094_),
    .B1(_1725_));
 sg13g2_a21oi_1 _2694_ (.A1(_1722_),
    .A2(net55),
    .Y(_1726_),
    .B1(net54));
 sg13g2_nor3_1 _2695_ (.A(_1717_),
    .B(_1706_),
    .C(_1726_),
    .Y(_0095_));
 sg13g2_nor2_1 _2696_ (.A(net72),
    .B(_1706_),
    .Y(_1727_));
 sg13g2_nor2_1 _2697_ (.A(_1690_),
    .B(_1707_),
    .Y(_1728_));
 sg13g2_nor3_1 _2698_ (.A(_1717_),
    .B(_1727_),
    .C(_1728_),
    .Y(_0096_));
 sg13g2_inv_1 _2699_ (.Y(_1729_),
    .A(_1611_));
 sg13g2_inv_1 _2700_ (.Y(_1730_),
    .A(net70));
 sg13g2_nor4_1 _2701_ (.A(_1730_),
    .B(_1690_),
    .C(_1699_),
    .D(_1702_),
    .Y(_1731_));
 sg13g2_nand3_1 _2702_ (.B(net71),
    .C(_1731_),
    .A(_1729_),
    .Y(_1732_));
 sg13g2_inv_1 _2703_ (.Y(_1733_),
    .A(_1732_));
 sg13g2_nor2_1 _2704_ (.A(net71),
    .B(_1728_),
    .Y(_1734_));
 sg13g2_nor3_1 _2705_ (.A(_1717_),
    .B(_1733_),
    .C(_1734_),
    .Y(_0097_));
 sg13g2_nor2_1 _2706_ (.A(_1694_),
    .B(_1732_),
    .Y(_1735_));
 sg13g2_nor2_1 _2707_ (.A(_1693_),
    .B(_1733_),
    .Y(_1736_));
 sg13g2_nor3_1 _2708_ (.A(_1717_),
    .B(_1735_),
    .C(_1736_),
    .Y(_0098_));
 sg13g2_nor2_1 _2709_ (.A(_1709_),
    .B(_1735_),
    .Y(_1737_));
 sg13g2_inv_1 _2710_ (.Y(_1738_),
    .A(_1710_));
 sg13g2_nor3_1 _2711_ (.A(_1717_),
    .B(_1737_),
    .C(_1738_),
    .Y(_0099_));
 sg13g2_nor2_1 _2712_ (.A(_1687_),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_nor3_1 _2713_ (.A(_1717_),
    .B(_1711_),
    .C(_1739_),
    .Y(_0100_));
 sg13g2_xnor2_1 _2714_ (.Y(_1740_),
    .A(\lfsr[29] ),
    .B(\lfsr[31] ));
 sg13g2_xor2_1 _2715_ (.B(\lfsr[24] ),
    .A(\lfsr[25] ),
    .X(_1741_));
 sg13g2_a21oi_1 _2716_ (.A1(_1741_),
    .A2(_1740_),
    .Y(_1742_),
    .B1(_1360_));
 sg13g2_o21ai_1 _2717_ (.B1(_1742_),
    .Y(_0131_),
    .A1(_1740_),
    .A2(_1741_));
 sg13g2_buf_1 _2718_ (.A(net77),
    .X(_1743_));
 sg13g2_nand2b_1 _2719_ (.Y(_0132_),
    .B(net69),
    .A_N(\lfsr[9] ));
 sg13g2_inv_1 _2720_ (.Y(_1744_),
    .A(\lfsr[10] ));
 sg13g2_nand2_1 _2721_ (.Y(_0133_),
    .A(_1744_),
    .B(net69));
 sg13g2_nand2b_1 _2722_ (.Y(_0134_),
    .B(net69),
    .A_N(\lfsr[11] ));
 sg13g2_nand2b_1 _2723_ (.Y(_0135_),
    .B(net69),
    .A_N(\lfsr[12] ));
 sg13g2_nand2b_1 _2724_ (.Y(_0136_),
    .B(net69),
    .A_N(\lfsr[13] ));
 sg13g2_nand2b_1 _2725_ (.Y(_0137_),
    .B(net69),
    .A_N(\lfsr[14] ));
 sg13g2_buf_1 _2726_ (.A(net77),
    .X(_1745_));
 sg13g2_nand2b_1 _2727_ (.Y(_0138_),
    .B(net68),
    .A_N(\lfsr[15] ));
 sg13g2_nand2b_1 _2728_ (.Y(_0139_),
    .B(net68),
    .A_N(\lfsr[16] ));
 sg13g2_nand2b_1 _2729_ (.Y(_0140_),
    .B(_1745_),
    .A_N(\lfsr[17] ));
 sg13g2_inv_1 _2730_ (.Y(_1746_),
    .A(\lfsr[18] ));
 sg13g2_nand2_1 _2731_ (.Y(_0141_),
    .A(_1746_),
    .B(net69));
 sg13g2_nand2b_1 _2732_ (.Y(_0142_),
    .B(_1745_),
    .A_N(\lfsr[0] ));
 sg13g2_inv_1 _2733_ (.Y(_1747_),
    .A(\lfsr[19] ));
 sg13g2_nand2_1 _2734_ (.Y(_0143_),
    .A(_1747_),
    .B(_1743_));
 sg13g2_nand2b_1 _2735_ (.Y(_0144_),
    .B(net68),
    .A_N(\lfsr[20] ));
 sg13g2_nand2b_1 _2736_ (.Y(_0145_),
    .B(net68),
    .A_N(\lfsr[21] ));
 sg13g2_nand2b_1 _2737_ (.Y(_0146_),
    .B(net68),
    .A_N(\lfsr[22] ));
 sg13g2_nand2b_1 _2738_ (.Y(_0147_),
    .B(net68),
    .A_N(\lfsr[23] ));
 sg13g2_nand2b_1 _2739_ (.Y(_0148_),
    .B(net68),
    .A_N(\lfsr[24] ));
 sg13g2_nand2b_1 _2740_ (.Y(_0149_),
    .B(net68),
    .A_N(\lfsr[25] ));
 sg13g2_buf_1 _2741_ (.A(net77),
    .X(_1748_));
 sg13g2_nand2b_1 _2742_ (.Y(_0150_),
    .B(net67),
    .A_N(\lfsr[26] ));
 sg13g2_nand2b_1 _2743_ (.Y(_0151_),
    .B(net67),
    .A_N(\lfsr[27] ));
 sg13g2_nand2b_1 _2744_ (.Y(_0152_),
    .B(net67),
    .A_N(\lfsr[28] ));
 sg13g2_nand2b_1 _2745_ (.Y(_0153_),
    .B(_1748_),
    .A_N(\lfsr[1] ));
 sg13g2_nand2b_1 _2746_ (.Y(_0154_),
    .B(net67),
    .A_N(\lfsr[29] ));
 sg13g2_nand2b_1 _2747_ (.Y(_0155_),
    .B(net67),
    .A_N(\lfsr[30] ));
 sg13g2_inv_1 _2748_ (.Y(_1749_),
    .A(\lfsr[2] ));
 sg13g2_nand2_1 _2749_ (.Y(_0156_),
    .A(_1749_),
    .B(net69));
 sg13g2_inv_1 _2750_ (.Y(_1750_),
    .A(\lfsr[3] ));
 sg13g2_nand2_1 _2751_ (.Y(_0157_),
    .A(_1750_),
    .B(_1743_));
 sg13g2_nand2b_1 _2752_ (.Y(_0158_),
    .B(_1748_),
    .A_N(\lfsr[4] ));
 sg13g2_nand2b_1 _2753_ (.Y(_0159_),
    .B(net67),
    .A_N(\lfsr[5] ));
 sg13g2_nand2b_1 _2754_ (.Y(_0160_),
    .B(net67),
    .A_N(\lfsr[6] ));
 sg13g2_nand2b_1 _2755_ (.Y(_0161_),
    .B(net67),
    .A_N(\lfsr[7] ));
 sg13g2_nand2b_1 _2756_ (.Y(_0162_),
    .B(net77),
    .A_N(\lfsr[8] ));
 sg13g2_nand2_1 _2757_ (.Y(_1751_),
    .A(_1412_),
    .B(net4));
 sg13g2_inv_1 _2758_ (.Y(_0163_),
    .A(_1751_));
 sg13g2_xnor2_1 _2759_ (.Y(\i_project.controller_0.vga_sync.o_vsync ),
    .A(_1456_),
    .B(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_buf_1 _2760_ (.A(_0037_),
    .X(_1752_));
 sg13g2_inv_2 _2761_ (.Y(_1753_),
    .A(_1752_));
 sg13g2_nand2_2 _2762_ (.Y(_1754_),
    .A(_1487_),
    .B(\i_project.controller_0.voffset[0] ));
 sg13g2_nor2_1 _2763_ (.A(net73),
    .B(_1539_),
    .Y(_1755_));
 sg13g2_nand2_1 _2764_ (.Y(_1756_),
    .A(_1486_),
    .B(_1539_));
 sg13g2_o21ai_1 _2765_ (.B1(_1756_),
    .Y(_1757_),
    .A1(_1754_),
    .A2(_1755_));
 sg13g2_xnor2_1 _2766_ (.Y(_1758_),
    .A(_1470_),
    .B(\i_project.controller_0.voffset[5] ));
 sg13g2_xnor2_1 _2767_ (.Y(_1759_),
    .A(_1469_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nor2_1 _2768_ (.A(_1758_),
    .B(_1759_),
    .Y(_1760_));
 sg13g2_xnor2_1 _2769_ (.Y(_1761_),
    .A(_1482_),
    .B(\i_project.controller_0.voffset[2] ));
 sg13g2_nand2_1 _2770_ (.Y(_1762_),
    .A(_1485_),
    .B(_1543_));
 sg13g2_nand2_1 _2771_ (.Y(_1763_),
    .A(_1484_),
    .B(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_2 _2772_ (.Y(_1764_),
    .A(_1762_),
    .B(_1763_));
 sg13g2_nor2_1 _2773_ (.A(_1761_),
    .B(_1764_),
    .Y(_1765_));
 sg13g2_nand3_1 _2774_ (.B(_1760_),
    .C(_1765_),
    .A(_1757_),
    .Y(_1766_));
 sg13g2_nand2_1 _2775_ (.Y(_1767_),
    .A(_1482_),
    .B(\i_project.controller_0.voffset[2] ));
 sg13g2_nor2_1 _2776_ (.A(_1484_),
    .B(\i_project.controller_0.voffset[3] ),
    .Y(_1768_));
 sg13g2_a21oi_1 _2777_ (.A1(_1763_),
    .A2(_1767_),
    .Y(_1769_),
    .B1(_1768_));
 sg13g2_nand2_1 _2778_ (.Y(_1770_),
    .A(_1469_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nor2_1 _2779_ (.A(_1470_),
    .B(\i_project.controller_0.voffset[5] ),
    .Y(_1771_));
 sg13g2_nand2_1 _2780_ (.Y(_1772_),
    .A(_1470_),
    .B(\i_project.controller_0.voffset[5] ));
 sg13g2_o21ai_1 _2781_ (.B1(_1772_),
    .Y(_1773_),
    .A1(_1770_),
    .A2(_1771_));
 sg13g2_a21oi_1 _2782_ (.A1(_1760_),
    .A2(_1769_),
    .Y(_1774_),
    .B1(_1773_));
 sg13g2_nand2_1 _2783_ (.Y(_1775_),
    .A(_1766_),
    .B(_1774_));
 sg13g2_nor2_1 _2784_ (.A(_1474_),
    .B(\i_project.controller_0.voffset[6] ),
    .Y(_1776_));
 sg13g2_nand2_1 _2785_ (.Y(_1777_),
    .A(_1474_),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_nor2b_1 _2786_ (.A(_1776_),
    .B_N(_1777_),
    .Y(_1778_));
 sg13g2_nand2_1 _2787_ (.Y(_1779_),
    .A(_1775_),
    .B(_1778_));
 sg13g2_inv_1 _2788_ (.Y(_1780_),
    .A(_1778_));
 sg13g2_nand3_1 _2789_ (.B(_1774_),
    .C(_1780_),
    .A(_1766_),
    .Y(_1781_));
 sg13g2_nand2_1 _2790_ (.Y(_1782_),
    .A(_1779_),
    .B(_1781_));
 sg13g2_buf_8 _2791_ (.A(_1782_),
    .X(_1783_));
 sg13g2_xnor2_1 _2792_ (.Y(_1784_),
    .A(_1753_),
    .B(_1783_));
 sg13g2_xor2_1 _2793_ (.B(_1709_),
    .A(net75),
    .X(_1785_));
 sg13g2_nand2_1 _2794_ (.Y(_1786_),
    .A(net58),
    .B(net54));
 sg13g2_xnor2_1 _2795_ (.Y(_1787_),
    .A(net57),
    .B(net72));
 sg13g2_nand2_1 _2796_ (.Y(_1788_),
    .A(net57),
    .B(net72));
 sg13g2_o21ai_1 _2797_ (.B1(_1788_),
    .Y(_1789_),
    .A1(_1786_),
    .A2(_1787_));
 sg13g2_xor2_1 _2798_ (.B(_1693_),
    .A(_1428_),
    .X(_1790_));
 sg13g2_inv_1 _2799_ (.Y(_1791_),
    .A(_1790_));
 sg13g2_xor2_1 _2800_ (.B(net71),
    .A(_1430_),
    .X(_1792_));
 sg13g2_inv_1 _2801_ (.Y(_1793_),
    .A(_1792_));
 sg13g2_nor2_1 _2802_ (.A(_1791_),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_nand2_1 _2803_ (.Y(_1795_),
    .A(net59),
    .B(net71));
 sg13g2_nor2_1 _2804_ (.A(_1795_),
    .B(_1791_),
    .Y(_1796_));
 sg13g2_a221oi_1 _2805_ (.B2(_1794_),
    .C1(_1796_),
    .B1(_1789_),
    .A1(net60),
    .Y(_1797_),
    .A2(_1693_));
 sg13g2_nand2_1 _2806_ (.Y(_1798_),
    .A(net62),
    .B(net70));
 sg13g2_xnor2_1 _2807_ (.Y(_1799_),
    .A(net63),
    .B(net55));
 sg13g2_nand2_1 _2808_ (.Y(_1800_),
    .A(net63),
    .B(net55));
 sg13g2_o21ai_1 _2809_ (.B1(_1800_),
    .Y(_1801_),
    .A1(_1798_),
    .A2(_1799_));
 sg13g2_buf_1 _2810_ (.A(_1801_),
    .X(_1802_));
 sg13g2_xor2_1 _2811_ (.B(net54),
    .A(net58),
    .X(_1803_));
 sg13g2_inv_1 _2812_ (.Y(_1804_),
    .A(_1803_));
 sg13g2_nor2_1 _2813_ (.A(_1787_),
    .B(_1804_),
    .Y(_1805_));
 sg13g2_nand3_1 _2814_ (.B(_1805_),
    .C(_1794_),
    .A(_1802_),
    .Y(_1806_));
 sg13g2_nand2_1 _2815_ (.Y(_1807_),
    .A(_1797_),
    .B(_1806_));
 sg13g2_xnor2_1 _2816_ (.Y(_1808_),
    .A(_1785_),
    .B(_1807_));
 sg13g2_xor2_1 _2817_ (.B(_1808_),
    .A(_1784_),
    .X(_1809_));
 sg13g2_buf_1 _2818_ (.A(_0038_),
    .X(_1810_));
 sg13g2_nor2_1 _2819_ (.A(_1482_),
    .B(\i_project.controller_0.voffset[2] ),
    .Y(_1811_));
 sg13g2_o21ai_1 _2820_ (.B1(_1767_),
    .Y(_1812_),
    .A1(_1756_),
    .A2(_1811_));
 sg13g2_nor2_1 _2821_ (.A(_1759_),
    .B(_1764_),
    .Y(_1813_));
 sg13g2_nor2_1 _2822_ (.A(_1469_),
    .B(\i_project.controller_0.voffset[4] ),
    .Y(_1814_));
 sg13g2_o21ai_1 _2823_ (.B1(_1770_),
    .Y(_1815_),
    .A1(_1763_),
    .A2(_1814_));
 sg13g2_a21oi_1 _2824_ (.A1(_1812_),
    .A2(_1813_),
    .Y(_1816_),
    .B1(_1815_));
 sg13g2_xnor2_1 _2825_ (.Y(_1817_),
    .A(net73),
    .B(_1539_));
 sg13g2_nor2_1 _2826_ (.A(_1817_),
    .B(_1761_),
    .Y(_1818_));
 sg13g2_inv_2 _2827_ (.Y(_1819_),
    .A(_1754_));
 sg13g2_nand3_1 _2828_ (.B(_1813_),
    .C(_1819_),
    .A(_1818_),
    .Y(_1820_));
 sg13g2_nand2_1 _2829_ (.Y(_1821_),
    .A(_1816_),
    .B(_1820_));
 sg13g2_inv_1 _2830_ (.Y(_1822_),
    .A(_1758_));
 sg13g2_nand2_1 _2831_ (.Y(_1823_),
    .A(_1821_),
    .B(_1822_));
 sg13g2_nand3_1 _2832_ (.B(_1820_),
    .C(_1758_),
    .A(_1816_),
    .Y(_1824_));
 sg13g2_nand2_1 _2833_ (.Y(_1825_),
    .A(_1823_),
    .B(_1824_));
 sg13g2_buf_8 _2834_ (.A(_1825_),
    .X(_1826_));
 sg13g2_nor2_1 _2835_ (.A(_1810_),
    .B(_1826_),
    .Y(_1827_));
 sg13g2_buf_2 _2836_ (.A(_0039_),
    .X(_1828_));
 sg13g2_nand2_1 _2837_ (.Y(_1829_),
    .A(_1757_),
    .B(_1765_));
 sg13g2_inv_1 _2838_ (.Y(_1830_),
    .A(_1769_));
 sg13g2_nand2_1 _2839_ (.Y(_1831_),
    .A(_1829_),
    .B(_1830_));
 sg13g2_inv_1 _2840_ (.Y(_1832_),
    .A(_1759_));
 sg13g2_nand2_1 _2841_ (.Y(_1833_),
    .A(_1831_),
    .B(_1832_));
 sg13g2_nand3_1 _2842_ (.B(_1759_),
    .C(_1830_),
    .A(_1829_),
    .Y(_1834_));
 sg13g2_nand2_2 _2843_ (.Y(_1835_),
    .A(_1833_),
    .B(_1834_));
 sg13g2_buf_8 _2844_ (.A(_1835_),
    .X(_1836_));
 sg13g2_nor2_1 _2845_ (.A(_1828_),
    .B(net25),
    .Y(_1837_));
 sg13g2_inv_1 _2846_ (.Y(_1838_),
    .A(_1539_));
 sg13g2_nand2_1 _2847_ (.Y(_1839_),
    .A(_1500_),
    .B(_1838_));
 sg13g2_inv_1 _2848_ (.Y(_1840_),
    .A(_1756_));
 sg13g2_a21oi_1 _2849_ (.A1(_1819_),
    .A2(_1839_),
    .Y(_1841_),
    .B1(_1840_));
 sg13g2_nand2_1 _2850_ (.Y(_1842_),
    .A(_1841_),
    .B(_1761_));
 sg13g2_inv_1 _2851_ (.Y(_1843_),
    .A(_1761_));
 sg13g2_nand2_1 _2852_ (.Y(_1844_),
    .A(_1757_),
    .B(_1843_));
 sg13g2_nand2_1 _2853_ (.Y(_1845_),
    .A(_1842_),
    .B(_1844_));
 sg13g2_buf_8 _2854_ (.A(_1845_),
    .X(_1846_));
 sg13g2_xor2_1 _2855_ (.B(_1539_),
    .A(net73),
    .X(_1847_));
 sg13g2_nand2_1 _2856_ (.Y(_1848_),
    .A(_1847_),
    .B(_1819_));
 sg13g2_nand2_1 _2857_ (.Y(_1849_),
    .A(_1817_),
    .B(_1754_));
 sg13g2_nand2_1 _2858_ (.Y(_1850_),
    .A(_1848_),
    .B(_1849_));
 sg13g2_buf_8 _2859_ (.A(_1850_),
    .X(_1851_));
 sg13g2_xnor2_1 _2860_ (.Y(_1852_),
    .A(\i_project.controller_0.mode_ramp_base[2] ),
    .B(net41));
 sg13g2_nand2_1 _2861_ (.Y(_1853_),
    .A(_1589_),
    .B(_1504_));
 sg13g2_nand2_1 _2862_ (.Y(_1854_),
    .A(_1853_),
    .B(_1754_));
 sg13g2_buf_1 _2863_ (.A(_1854_),
    .X(_1855_));
 sg13g2_nor2_1 _2864_ (.A(_1719_),
    .B(net45),
    .Y(_1856_));
 sg13g2_nand2_1 _2865_ (.Y(_1857_),
    .A(_1852_),
    .B(_1856_));
 sg13g2_o21ai_1 _2866_ (.B1(_1857_),
    .Y(_1858_),
    .A1(_0042_),
    .A2(net41));
 sg13g2_xnor2_1 _2867_ (.Y(_1859_),
    .A(net55),
    .B(net36));
 sg13g2_nand2_1 _2868_ (.Y(_1860_),
    .A(_1858_),
    .B(_1859_));
 sg13g2_o21ai_1 _2869_ (.B1(_1860_),
    .Y(_1861_),
    .A1(_0041_),
    .A2(net36));
 sg13g2_buf_1 _2870_ (.A(_0040_),
    .X(_1862_));
 sg13g2_inv_1 _2871_ (.Y(_1863_),
    .A(_1862_));
 sg13g2_nand2_1 _2872_ (.Y(_1864_),
    .A(_1767_),
    .B(_1756_));
 sg13g2_inv_1 _2873_ (.Y(_1865_),
    .A(_1864_));
 sg13g2_nand2_1 _2874_ (.Y(_1866_),
    .A(_1848_),
    .B(_1865_));
 sg13g2_inv_1 _2875_ (.Y(_1867_),
    .A(_1811_));
 sg13g2_nand2_1 _2876_ (.Y(_1868_),
    .A(_1866_),
    .B(_1867_));
 sg13g2_nand2_1 _2877_ (.Y(_1869_),
    .A(_1868_),
    .B(_1764_));
 sg13g2_inv_1 _2878_ (.Y(_1870_),
    .A(_1764_));
 sg13g2_nand3_1 _2879_ (.B(_1867_),
    .C(_1870_),
    .A(_1866_),
    .Y(_1871_));
 sg13g2_nand2_1 _2880_ (.Y(_1872_),
    .A(_1869_),
    .B(_1871_));
 sg13g2_buf_1 _2881_ (.A(_1872_),
    .X(_1873_));
 sg13g2_xnor2_1 _2882_ (.Y(_1874_),
    .A(_1863_),
    .B(net28));
 sg13g2_nand2_1 _2883_ (.Y(_1875_),
    .A(_1861_),
    .B(_1874_));
 sg13g2_nand2_1 _2884_ (.Y(_1876_),
    .A(_1868_),
    .B(_1870_));
 sg13g2_nand3_1 _2885_ (.B(_1867_),
    .C(_1764_),
    .A(_1866_),
    .Y(_1877_));
 sg13g2_nand2_2 _2886_ (.Y(_1878_),
    .A(_1876_),
    .B(_1877_));
 sg13g2_nand2_1 _2887_ (.Y(_1879_),
    .A(_1878_),
    .B(_1863_));
 sg13g2_nand2_1 _2888_ (.Y(_1880_),
    .A(_1875_),
    .B(_1879_));
 sg13g2_xnor2_1 _2889_ (.Y(_1881_),
    .A(_1689_),
    .B(net25));
 sg13g2_nand2_1 _2890_ (.Y(_1882_),
    .A(_1880_),
    .B(_1881_));
 sg13g2_nand2b_1 _2891_ (.Y(_1883_),
    .B(_1882_),
    .A_N(_1837_));
 sg13g2_xnor2_1 _2892_ (.Y(_1884_),
    .A(_1691_),
    .B(_1826_));
 sg13g2_nand2_1 _2893_ (.Y(_1885_),
    .A(_1883_),
    .B(_1884_));
 sg13g2_nand2b_1 _2894_ (.Y(_1886_),
    .B(_1885_),
    .A_N(_1827_));
 sg13g2_nor2_1 _2895_ (.A(_1809_),
    .B(_1886_),
    .Y(_1887_));
 sg13g2_nand2_1 _2896_ (.Y(_1888_),
    .A(_1886_),
    .B(_1809_));
 sg13g2_nor3_1 _2897_ (.A(_1520_),
    .B(_1553_),
    .C(_1534_),
    .Y(_1889_));
 sg13g2_buf_2 _2898_ (.A(_1889_),
    .X(_1890_));
 sg13g2_buf_1 _2899_ (.A(_1890_),
    .X(_1891_));
 sg13g2_nand2_1 _2900_ (.Y(_1892_),
    .A(_1888_),
    .B(net44));
 sg13g2_nor3_1 _2901_ (.A(_1523_),
    .B(_0029_),
    .C(_1555_),
    .Y(_1893_));
 sg13g2_buf_2 _2902_ (.A(_1893_),
    .X(_1894_));
 sg13g2_inv_2 _2903_ (.Y(_0165_),
    .A(_1894_));
 sg13g2_nor3_1 _2904_ (.A(_1520_),
    .B(_1523_),
    .C(_1534_),
    .Y(_0166_));
 sg13g2_buf_8 _2905_ (.A(_0166_),
    .X(_0167_));
 sg13g2_inv_2 _2906_ (.Y(_0168_),
    .A(_0167_));
 sg13g2_nand2_1 _2907_ (.Y(_0169_),
    .A(_0165_),
    .B(_0168_));
 sg13g2_buf_2 _2908_ (.A(_0169_),
    .X(_0170_));
 sg13g2_a21oi_1 _2909_ (.A1(_1565_),
    .A2(_1352_),
    .Y(_0171_),
    .B1(_1356_));
 sg13g2_buf_1 _2910_ (.A(_1351_),
    .X(_0172_));
 sg13g2_nand2b_1 _2911_ (.Y(_0173_),
    .B(net53),
    .A_N(_0017_));
 sg13g2_nand2_1 _2912_ (.Y(_0174_),
    .A(_1514_),
    .B(_1351_));
 sg13g2_o21ai_1 _2913_ (.B1(_0174_),
    .Y(_0175_),
    .A1(_0172_),
    .A2(_0047_));
 sg13g2_inv_1 _2914_ (.Y(_0176_),
    .A(_0175_));
 sg13g2_a22oi_1 _2915_ (.Y(_0177_),
    .B1(net65),
    .B2(_0176_),
    .A2(_0173_),
    .A1(_0171_));
 sg13g2_inv_1 _2916_ (.Y(_0178_),
    .A(_0177_));
 sg13g2_xnor2_1 _2917_ (.Y(_0179_),
    .A(net75),
    .B(_1783_));
 sg13g2_a21oi_1 _2918_ (.A1(_0179_),
    .A2(_1894_),
    .Y(_0180_),
    .B1(_1890_));
 sg13g2_o21ai_1 _2919_ (.B1(_0180_),
    .Y(_0181_),
    .A1(_0170_),
    .A2(_0178_));
 sg13g2_o21ai_1 _2920_ (.B1(_0181_),
    .Y(_0182_),
    .A1(_1887_),
    .A2(_1892_));
 sg13g2_inv_1 _2921_ (.Y(_0183_),
    .A(_1783_));
 sg13g2_nor2_1 _2922_ (.A(_0047_),
    .B(_0168_),
    .Y(_0184_));
 sg13g2_nor3_1 _2923_ (.A(_1523_),
    .B(_1555_),
    .C(_1525_),
    .Y(_0185_));
 sg13g2_buf_2 _2924_ (.A(_0185_),
    .X(_0186_));
 sg13g2_buf_8 _2925_ (.A(_0186_),
    .X(_0187_));
 sg13g2_a21oi_1 _2926_ (.A1(_0183_),
    .A2(_0184_),
    .Y(_0188_),
    .B1(net43));
 sg13g2_nand2_1 _2927_ (.Y(_0189_),
    .A(_0182_),
    .B(_0188_));
 sg13g2_nand2_1 _2928_ (.Y(_0190_),
    .A(_1352_),
    .B(_0049_));
 sg13g2_a21oi_1 _2929_ (.A1(_1351_),
    .A2(_0035_),
    .Y(_0191_),
    .B1(_1355_));
 sg13g2_nand2_1 _2930_ (.Y(_0192_),
    .A(_1510_),
    .B(_1351_));
 sg13g2_o21ai_1 _2931_ (.B1(_0192_),
    .Y(_0193_),
    .A1(_1351_),
    .A2(_0034_));
 sg13g2_a22oi_1 _2932_ (.Y(_0194_),
    .B1(net76),
    .B2(_0193_),
    .A2(_0191_),
    .A1(_0190_));
 sg13g2_buf_1 _2933_ (.A(_0194_),
    .X(_0195_));
 sg13g2_nor2_1 _2934_ (.A(_1478_),
    .B(_1477_),
    .Y(_0196_));
 sg13g2_nand2_1 _2935_ (.Y(_0197_),
    .A(_0195_),
    .B(_0196_));
 sg13g2_o21ai_1 _2936_ (.B1(_0049_),
    .Y(_0198_),
    .A1(_1478_),
    .A2(_1477_));
 sg13g2_nand2_1 _2937_ (.Y(_0199_),
    .A(_0197_),
    .B(_0198_));
 sg13g2_buf_1 _2938_ (.A(_0199_),
    .X(_0200_));
 sg13g2_xnor2_1 _2939_ (.Y(_0201_),
    .A(net27),
    .B(_1783_));
 sg13g2_nor3_2 _2940_ (.A(_1520_),
    .B(_1553_),
    .C(_1525_),
    .Y(_0202_));
 sg13g2_buf_8 _2941_ (.A(_0202_),
    .X(_0203_));
 sg13g2_a21oi_1 _2942_ (.A1(_0201_),
    .A2(net43),
    .Y(_0204_),
    .B1(net48));
 sg13g2_nand2_1 _2943_ (.Y(_0205_),
    .A(_0189_),
    .B(_0204_));
 sg13g2_nor2_1 _2944_ (.A(_1444_),
    .B(_1450_),
    .Y(_0206_));
 sg13g2_buf_8 _2945_ (.A(_0206_),
    .X(_0207_));
 sg13g2_a21oi_1 _2946_ (.A1(_0183_),
    .A2(net48),
    .Y(_0208_),
    .B1(net35));
 sg13g2_nand2_1 _2947_ (.Y(_0209_),
    .A(_0205_),
    .B(_0208_));
 sg13g2_nor2_1 _2948_ (.A(_1758_),
    .B(_1780_),
    .Y(_0210_));
 sg13g2_o21ai_1 _2949_ (.B1(_1777_),
    .Y(_0211_),
    .A1(_1772_),
    .A2(_1776_));
 sg13g2_a21oi_1 _2950_ (.A1(_1821_),
    .A2(_0210_),
    .Y(_0212_),
    .B1(_0211_));
 sg13g2_nor2_1 _2951_ (.A(_1472_),
    .B(\i_project.controller_0.voffset[7] ),
    .Y(_0213_));
 sg13g2_nand2_1 _2952_ (.Y(_0214_),
    .A(_1472_),
    .B(\i_project.controller_0.voffset[7] ));
 sg13g2_inv_1 _2953_ (.Y(_0215_),
    .A(_0214_));
 sg13g2_nor2_1 _2954_ (.A(_0213_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_nand2b_1 _2955_ (.Y(_0217_),
    .B(_0216_),
    .A_N(_0212_));
 sg13g2_nand2b_1 _2956_ (.Y(_0218_),
    .B(_0212_),
    .A_N(_0216_));
 sg13g2_nand2_1 _2957_ (.Y(_0219_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_buf_8 _2958_ (.A(_0219_),
    .X(_0220_));
 sg13g2_a21oi_1 _2959_ (.A1(_0183_),
    .A2(net62),
    .Y(_0221_),
    .B1(_1415_));
 sg13g2_o21ai_1 _2960_ (.B1(_0221_),
    .Y(_0222_),
    .A1(_1417_),
    .A2(_0220_));
 sg13g2_a22oi_1 _2961_ (.Y(_0223_),
    .B1(_1461_),
    .B2(_1826_),
    .A2(net25),
    .A1(_1570_));
 sg13g2_nand2_1 _2962_ (.Y(_0224_),
    .A(_0222_),
    .B(_0223_));
 sg13g2_inv_1 _2963_ (.Y(_0225_),
    .A(_1846_));
 sg13g2_a21oi_1 _2964_ (.A1(_0225_),
    .A2(net62),
    .Y(_0226_),
    .B1(_1415_));
 sg13g2_o21ai_1 _2965_ (.B1(_0226_),
    .Y(_0227_),
    .A1(net62),
    .A2(net28));
 sg13g2_a22oi_1 _2966_ (.Y(_0228_),
    .B1(_1461_),
    .B2(net41),
    .A2(_1855_),
    .A1(_1570_));
 sg13g2_a21oi_1 _2967_ (.A1(_0227_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(net61));
 sg13g2_a21oi_1 _2968_ (.A1(_0224_),
    .A2(_1420_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_nand2b_1 _2969_ (.Y(_0231_),
    .B(_0215_),
    .A_N(_0032_));
 sg13g2_o21ai_1 _2970_ (.B1(_0231_),
    .Y(_0232_),
    .A1(_1479_),
    .A2(_0217_));
 sg13g2_nand2b_1 _2971_ (.Y(_0233_),
    .B(_1477_),
    .A_N(_0232_));
 sg13g2_inv_1 _2972_ (.Y(_0234_),
    .A(net62));
 sg13g2_nand2_1 _2973_ (.Y(_0235_),
    .A(_0232_),
    .B(_1494_));
 sg13g2_nand3_1 _2974_ (.B(_0234_),
    .C(_0235_),
    .A(_0233_),
    .Y(_0236_));
 sg13g2_nand2_1 _2975_ (.Y(_0237_),
    .A(_0214_),
    .B(_1777_));
 sg13g2_inv_1 _2976_ (.Y(_0238_),
    .A(_0237_));
 sg13g2_a21oi_1 _2977_ (.A1(_1779_),
    .A2(_0238_),
    .Y(_0239_),
    .B1(_0213_));
 sg13g2_xnor2_1 _2978_ (.Y(_0240_),
    .A(_1478_),
    .B(_0239_));
 sg13g2_nor2b_1 _2979_ (.A(_0234_),
    .B_N(_0240_),
    .Y(_0241_));
 sg13g2_nor3_1 _2980_ (.A(_0035_),
    .B(_0034_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_a21o_1 _2981_ (.A2(_0242_),
    .A1(_0236_),
    .B1(net57),
    .X(_0243_));
 sg13g2_o21ai_1 _2982_ (.B1(_0243_),
    .Y(_0244_),
    .A1(_1422_),
    .A2(_0230_));
 sg13g2_nand2_1 _2983_ (.Y(_0245_),
    .A(_0244_),
    .B(net35));
 sg13g2_buf_8 _2984_ (.A(_0245_),
    .X(_0246_));
 sg13g2_nand2_1 _2985_ (.Y(_0247_),
    .A(_0209_),
    .B(_0246_));
 sg13g2_inv_4 _2986_ (.A(_1526_),
    .Y(_0248_));
 sg13g2_buf_8 _2987_ (.A(_0248_),
    .X(_0249_));
 sg13g2_nand2_1 _2988_ (.Y(_0250_),
    .A(_0247_),
    .B(net47));
 sg13g2_a21oi_1 _2989_ (.A1(_1493_),
    .A2(_1598_),
    .Y(_0251_),
    .B1(_1473_));
 sg13g2_nand4_1 _2990_ (.B(_1488_),
    .C(_1480_),
    .A(_1476_),
    .Y(_0252_),
    .D(_1598_));
 sg13g2_nor2_1 _2991_ (.A(_0031_),
    .B(_1475_),
    .Y(_0253_));
 sg13g2_a21oi_1 _2992_ (.A1(_1597_),
    .A2(_0253_),
    .Y(_0254_),
    .B1(_1477_));
 sg13g2_nand2_1 _2993_ (.Y(_0255_),
    .A(_0252_),
    .B(_0254_));
 sg13g2_a22oi_1 _2994_ (.Y(_0256_),
    .B1(_1457_),
    .B2(_0255_),
    .A2(_0251_),
    .A1(_1495_));
 sg13g2_nand2_1 _2995_ (.Y(_0257_),
    .A(_1518_),
    .B(_0256_));
 sg13g2_nand2_1 _2996_ (.Y(_0258_),
    .A(_0257_),
    .B(_0248_));
 sg13g2_buf_8 _2997_ (.A(_0258_),
    .X(_0259_));
 sg13g2_nand2_1 _2998_ (.Y(_0260_),
    .A(_1526_),
    .B(_0048_));
 sg13g2_buf_8 _2999_ (.A(_0260_),
    .X(_0261_));
 sg13g2_nand3_1 _3000_ (.B(_0259_),
    .C(_0261_),
    .A(_0250_),
    .Y(_0262_));
 sg13g2_buf_2 _3001_ (.A(_0262_),
    .X(_0263_));
 sg13g2_inv_4 _3002_ (.A(_0263_),
    .Y(_0264_));
 sg13g2_buf_1 _3003_ (.A(\depth[1] ),
    .X(_0265_));
 sg13g2_buf_8 _3004_ (.A(\depth[0] ),
    .X(_0266_));
 sg13g2_inv_1 _3005_ (.Y(_0267_),
    .A(_0266_));
 sg13g2_inv_1 _3006_ (.Y(_0268_),
    .A(_0043_));
 sg13g2_nor3_1 _3007_ (.A(_0265_),
    .B(_0267_),
    .C(_0268_),
    .Y(_0269_));
 sg13g2_buf_2 _3008_ (.A(_0269_),
    .X(_0270_));
 sg13g2_nand2_1 _3009_ (.Y(_0271_),
    .A(_0264_),
    .B(_0270_));
 sg13g2_nand2_1 _3010_ (.Y(_0272_),
    .A(_1884_),
    .B(_1784_));
 sg13g2_nand2b_1 _3011_ (.Y(_0273_),
    .B(_1883_),
    .A_N(_0272_));
 sg13g2_nor2_1 _3012_ (.A(_1752_),
    .B(_1783_),
    .Y(_0274_));
 sg13g2_a21oi_1 _3013_ (.A1(_1784_),
    .A2(_1827_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_xnor2_1 _3014_ (.Y(_0276_),
    .A(_1426_),
    .B(_0220_));
 sg13g2_inv_2 _3015_ (.Y(_0277_),
    .A(_0276_));
 sg13g2_xor2_1 _3016_ (.B(_0036_),
    .A(_1687_),
    .X(_0278_));
 sg13g2_inv_1 _3017_ (.Y(_0279_),
    .A(_1709_));
 sg13g2_nand2_1 _3018_ (.Y(_0280_),
    .A(_1807_),
    .B(_1785_));
 sg13g2_o21ai_1 _3019_ (.B1(_0280_),
    .Y(_0281_),
    .A1(_1425_),
    .A2(_0279_));
 sg13g2_xnor2_1 _3020_ (.Y(_0282_),
    .A(_0278_),
    .B(_0281_));
 sg13g2_xnor2_1 _3021_ (.Y(_0283_),
    .A(_0277_),
    .B(_0282_));
 sg13g2_a21oi_1 _3022_ (.A1(_0273_),
    .A2(_0275_),
    .Y(_0284_),
    .B1(_0283_));
 sg13g2_nand3_1 _3023_ (.B(_0273_),
    .C(_0275_),
    .A(_0283_),
    .Y(_0285_));
 sg13g2_nand3b_1 _3024_ (.B(net44),
    .C(_0285_),
    .Y(_0286_),
    .A_N(_0284_));
 sg13g2_nand2_1 _3025_ (.Y(_0287_),
    .A(_0026_),
    .B(_1351_));
 sg13g2_o21ai_1 _3026_ (.B1(_0287_),
    .Y(_0288_),
    .A1(_0172_),
    .A2(_1514_));
 sg13g2_inv_1 _3027_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_o21ai_1 _3028_ (.B1(net76),
    .Y(_0290_),
    .A1(net53),
    .A2(_1436_));
 sg13g2_o21ai_1 _3029_ (.B1(_0290_),
    .Y(_0291_),
    .A1(net76),
    .A2(_0289_));
 sg13g2_inv_1 _3030_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_inv_2 _3031_ (.Y(_0293_),
    .A(_1890_));
 sg13g2_o21ai_1 _3032_ (.B1(_0293_),
    .Y(_0294_),
    .A1(_0165_),
    .A2(_0277_));
 sg13g2_a21oi_1 _3033_ (.A1(_0165_),
    .A2(_0292_),
    .Y(_0295_),
    .B1(_0294_));
 sg13g2_nor2_1 _3034_ (.A(net49),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_nand2_1 _3035_ (.Y(_0297_),
    .A(_0286_),
    .B(_0296_));
 sg13g2_inv_1 _3036_ (.Y(_0298_),
    .A(_0220_));
 sg13g2_nor2_1 _3037_ (.A(_0028_),
    .B(_0168_),
    .Y(_0299_));
 sg13g2_a21oi_1 _3038_ (.A1(_0298_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(net43));
 sg13g2_nand2_1 _3039_ (.Y(_0301_),
    .A(_0297_),
    .B(_0300_));
 sg13g2_xnor2_1 _3040_ (.Y(_0302_),
    .A(net27),
    .B(_0220_));
 sg13g2_buf_1 _3041_ (.A(_0187_),
    .X(_0303_));
 sg13g2_buf_8 _3042_ (.A(_0203_),
    .X(_0304_));
 sg13g2_a21oi_1 _3043_ (.A1(_0302_),
    .A2(net40),
    .Y(_0305_),
    .B1(net42));
 sg13g2_nand2_1 _3044_ (.Y(_0306_),
    .A(_0301_),
    .B(_0305_));
 sg13g2_a21oi_1 _3045_ (.A1(_0298_),
    .A2(net42),
    .Y(_0307_),
    .B1(net35));
 sg13g2_nand2_1 _3046_ (.Y(_0308_),
    .A(_0306_),
    .B(_0307_));
 sg13g2_buf_8 _3047_ (.A(_0246_),
    .X(_0309_));
 sg13g2_nand2_1 _3048_ (.Y(_0310_),
    .A(_0308_),
    .B(net22));
 sg13g2_nand3_1 _3049_ (.B(_0248_),
    .C(_0256_),
    .A(_1518_),
    .Y(_0311_));
 sg13g2_o21ai_1 _3050_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_0033_),
    .A2(_0248_));
 sg13g2_buf_2 _3051_ (.A(_0312_),
    .X(_0313_));
 sg13g2_inv_1 _3052_ (.Y(_0314_),
    .A(_0313_));
 sg13g2_a21oi_1 _3053_ (.A1(_0310_),
    .A2(net47),
    .Y(_0315_),
    .B1(_0314_));
 sg13g2_buf_2 _3054_ (.A(_0315_),
    .X(_0316_));
 sg13g2_inv_1 _3055_ (.Y(_0317_),
    .A(_0265_));
 sg13g2_nor3_1 _3056_ (.A(_0266_),
    .B(_0317_),
    .C(_0268_),
    .Y(_0318_));
 sg13g2_buf_2 _3057_ (.A(_0318_),
    .X(_0319_));
 sg13g2_nand2_1 _3058_ (.Y(_0320_),
    .A(_0316_),
    .B(_0319_));
 sg13g2_a21oi_1 _3059_ (.A1(_0317_),
    .A2(_0267_),
    .Y(_0321_),
    .B1(_0268_));
 sg13g2_inv_1 _3060_ (.Y(_0322_),
    .A(\depth[2] ));
 sg13g2_nor3_1 _3061_ (.A(_0043_),
    .B(_0317_),
    .C(_0267_),
    .Y(_0323_));
 sg13g2_nor3_1 _3062_ (.A(_0266_),
    .B(_0317_),
    .C(_0322_),
    .Y(_0324_));
 sg13g2_nor2_1 _3063_ (.A(_0323_),
    .B(_0324_),
    .Y(_0325_));
 sg13g2_o21ai_1 _3064_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0265_),
    .A2(_0322_));
 sg13g2_nor2_1 _3065_ (.A(_0321_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_buf_2 _3066_ (.A(_0327_),
    .X(_0328_));
 sg13g2_buf_8 _3067_ (.A(_0328_),
    .X(_0329_));
 sg13g2_nand2_1 _3068_ (.Y(_0330_),
    .A(net52),
    .B(_0044_));
 sg13g2_inv_1 _3069_ (.Y(_0331_),
    .A(_0330_));
 sg13g2_inv_1 _3070_ (.Y(_0332_),
    .A(_0326_));
 sg13g2_inv_4 _3071_ (.A(_0259_),
    .Y(_0333_));
 sg13g2_nor2_1 _3072_ (.A(_0332_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_nor3_1 _3073_ (.A(_0317_),
    .B(_0267_),
    .C(_0268_),
    .Y(_0335_));
 sg13g2_inv_1 _3074_ (.Y(_0336_),
    .A(_0335_));
 sg13g2_nor2_1 _3075_ (.A(_0336_),
    .B(_0333_),
    .Y(_0337_));
 sg13g2_buf_2 _3076_ (.A(_0337_),
    .X(_0338_));
 sg13g2_nor2_1 _3077_ (.A(_0334_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_buf_1 _3078_ (.A(_0293_),
    .X(_0340_));
 sg13g2_a21o_1 _3079_ (.A2(_1805_),
    .A1(_1802_),
    .B1(_1789_),
    .X(_0341_));
 sg13g2_xnor2_1 _3080_ (.Y(_0342_),
    .A(_1793_),
    .B(_0341_));
 sg13g2_xnor2_1 _3081_ (.Y(_0343_),
    .A(_1881_),
    .B(_1880_));
 sg13g2_xnor2_1 _3082_ (.Y(_0344_),
    .A(_0342_),
    .B(_0343_));
 sg13g2_nand2_1 _3083_ (.Y(_0345_),
    .A(net53),
    .B(_0046_));
 sg13g2_inv_1 _3084_ (.Y(_0346_),
    .A(_0345_));
 sg13g2_a21oi_1 _3085_ (.A1(_1352_),
    .A2(_0045_),
    .Y(_0347_),
    .B1(_0346_));
 sg13g2_nand2_1 _3086_ (.Y(_0348_),
    .A(_0347_),
    .B(net65));
 sg13g2_o21ai_1 _3087_ (.B1(_0348_),
    .Y(_0349_),
    .A1(net65),
    .A2(_0176_));
 sg13g2_inv_1 _3088_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_xnor2_1 _3089_ (.Y(_0351_),
    .A(_1445_),
    .B(net25));
 sg13g2_inv_1 _3090_ (.Y(_0352_),
    .A(_0351_));
 sg13g2_a21oi_1 _3091_ (.A1(_0352_),
    .A2(_1894_),
    .Y(_0353_),
    .B1(_1890_));
 sg13g2_o21ai_1 _3092_ (.B1(_0353_),
    .Y(_0354_),
    .A1(_0170_),
    .A2(_0350_));
 sg13g2_o21ai_1 _3093_ (.B1(_0354_),
    .Y(_0355_),
    .A1(net39),
    .A2(_0344_));
 sg13g2_inv_1 _3094_ (.Y(_0356_),
    .A(_1836_));
 sg13g2_nor2_1 _3095_ (.A(_0045_),
    .B(_0168_),
    .Y(_0357_));
 sg13g2_a21oi_1 _3096_ (.A1(_0356_),
    .A2(_0357_),
    .Y(_0358_),
    .B1(net40));
 sg13g2_nand2_1 _3097_ (.Y(_0359_),
    .A(_0355_),
    .B(_0358_));
 sg13g2_inv_1 _3098_ (.Y(_0360_),
    .A(net42));
 sg13g2_buf_1 _3099_ (.A(net27),
    .X(_0361_));
 sg13g2_inv_2 _3100_ (.Y(_0362_),
    .A(net24));
 sg13g2_inv_2 _3101_ (.Y(_0363_),
    .A(net43));
 sg13g2_a21oi_1 _3102_ (.A1(_0362_),
    .A2(_1836_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_o21ai_1 _3103_ (.B1(_0364_),
    .Y(_0365_),
    .A1(net25),
    .A2(_0362_));
 sg13g2_nand3_1 _3104_ (.B(net38),
    .C(_0365_),
    .A(_0359_),
    .Y(_0366_));
 sg13g2_buf_1 _3105_ (.A(net42),
    .X(_0367_));
 sg13g2_buf_1 _3106_ (.A(net35),
    .X(_0368_));
 sg13g2_a21oi_1 _3107_ (.A1(_0356_),
    .A2(net37),
    .Y(_0369_),
    .B1(net29));
 sg13g2_nand2_1 _3108_ (.Y(_0370_),
    .A(_0366_),
    .B(_0369_));
 sg13g2_a21oi_1 _3109_ (.A1(_0370_),
    .A2(net22),
    .Y(_0371_),
    .B1(net52));
 sg13g2_nor3_1 _3110_ (.A(_0331_),
    .B(_0339_),
    .C(_0371_),
    .Y(_0372_));
 sg13g2_nor2_1 _3111_ (.A(net30),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nand3_1 _3112_ (.B(_0320_),
    .C(_0373_),
    .A(_0271_),
    .Y(_0374_));
 sg13g2_inv_2 _3113_ (.Y(_0375_),
    .A(_0328_));
 sg13g2_buf_8 _3114_ (.A(_0375_),
    .X(_0376_));
 sg13g2_nor2_2 _3115_ (.A(net26),
    .B(_0316_),
    .Y(_0377_));
 sg13g2_inv_2 _3116_ (.Y(_0378_),
    .A(_0377_));
 sg13g2_nand2_1 _3117_ (.Y(_0379_),
    .A(_0374_),
    .B(_0378_));
 sg13g2_inv_1 _3118_ (.Y(_0380_),
    .A(_1795_));
 sg13g2_a21oi_1 _3119_ (.A1(_0341_),
    .A2(_1792_),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_xnor2_1 _3120_ (.Y(_0382_),
    .A(_1790_),
    .B(_0381_));
 sg13g2_xnor2_1 _3121_ (.Y(_0383_),
    .A(_1884_),
    .B(_0382_));
 sg13g2_a21oi_1 _3122_ (.A1(_1883_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(_0293_));
 sg13g2_o21ai_1 _3123_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_1883_),
    .A2(_0383_));
 sg13g2_nor2b_1 _3124_ (.A(net53),
    .B_N(_0046_),
    .Y(_0386_));
 sg13g2_a21oi_1 _3125_ (.A1(net53),
    .A2(_0047_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_nor2_1 _3126_ (.A(net65),
    .B(_0288_),
    .Y(_0388_));
 sg13g2_a21o_1 _3127_ (.A2(_0387_),
    .A1(net65),
    .B1(_0388_),
    .X(_0389_));
 sg13g2_inv_1 _3128_ (.Y(_0390_),
    .A(_0389_));
 sg13g2_xnor2_1 _3129_ (.Y(_0391_),
    .A(_1429_),
    .B(_1826_));
 sg13g2_a21oi_1 _3130_ (.A1(_0391_),
    .A2(_1894_),
    .Y(_0392_),
    .B1(_1890_));
 sg13g2_o21ai_1 _3131_ (.B1(_0392_),
    .Y(_0393_),
    .A1(_0170_),
    .A2(_0390_));
 sg13g2_nand2_1 _3132_ (.Y(_0394_),
    .A(_0385_),
    .B(_0393_));
 sg13g2_nand2_1 _3133_ (.Y(_0395_),
    .A(_1821_),
    .B(_1758_));
 sg13g2_nand3_1 _3134_ (.B(_1820_),
    .C(_1822_),
    .A(_1816_),
    .Y(_0396_));
 sg13g2_nand2_2 _3135_ (.Y(_0397_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_nand3b_1 _3136_ (.B(_0397_),
    .C(_0167_),
    .Y(_0398_),
    .A_N(_0046_));
 sg13g2_nand3_1 _3137_ (.B(_0363_),
    .C(_0398_),
    .A(_0394_),
    .Y(_0399_));
 sg13g2_xnor2_1 _3138_ (.Y(_0400_),
    .A(net27),
    .B(_1826_));
 sg13g2_a21oi_1 _3139_ (.A1(_0400_),
    .A2(net40),
    .Y(_0401_),
    .B1(net42));
 sg13g2_nand2_1 _3140_ (.Y(_0402_),
    .A(_0399_),
    .B(_0401_));
 sg13g2_a21oi_1 _3141_ (.A1(_0397_),
    .A2(_0304_),
    .Y(_0403_),
    .B1(_0207_));
 sg13g2_nand2_1 _3142_ (.Y(_0404_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_nand2_1 _3143_ (.Y(_0405_),
    .A(_0404_),
    .B(net22));
 sg13g2_nand2_1 _3144_ (.Y(_0406_),
    .A(_0405_),
    .B(_0249_));
 sg13g2_nand2_2 _3145_ (.Y(_0407_),
    .A(_1526_),
    .B(_0020_));
 sg13g2_nand2_1 _3146_ (.Y(_0408_),
    .A(_0406_),
    .B(_0407_));
 sg13g2_nor2_1 _3147_ (.A(_0333_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nor3_2 _3148_ (.A(_0265_),
    .B(_0266_),
    .C(_0322_),
    .Y(_0410_));
 sg13g2_nand2_1 _3149_ (.Y(_0411_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_nand2_1 _3150_ (.Y(_0412_),
    .A(_0271_),
    .B(_0411_));
 sg13g2_inv_1 _3151_ (.Y(_0413_),
    .A(_0319_));
 sg13g2_nor3_1 _3152_ (.A(_0265_),
    .B(_0267_),
    .C(_0322_),
    .Y(_0414_));
 sg13g2_inv_1 _3153_ (.Y(_0415_),
    .A(_0414_));
 sg13g2_a21oi_1 _3154_ (.A1(_0413_),
    .A2(_0415_),
    .Y(_0416_),
    .B1(_0263_));
 sg13g2_nand2_1 _3155_ (.Y(_0417_),
    .A(_0310_),
    .B(net47));
 sg13g2_nand2_2 _3156_ (.Y(_0418_),
    .A(_0417_),
    .B(_0313_));
 sg13g2_inv_1 _3157_ (.Y(_0419_),
    .A(_0324_));
 sg13g2_inv_2 _3158_ (.Y(_0420_),
    .A(net29));
 sg13g2_o21ai_1 _3159_ (.B1(_0420_),
    .Y(_0421_),
    .A1(net45),
    .A2(_0360_));
 sg13g2_o21ai_1 _3160_ (.B1(net40),
    .Y(_0422_),
    .A1(net45),
    .A2(_0362_));
 sg13g2_a21oi_1 _3161_ (.A1(net45),
    .A2(_0362_),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_buf_1 _3162_ (.A(net49),
    .X(_0424_));
 sg13g2_nor2_1 _3163_ (.A(_0049_),
    .B(net45),
    .Y(_0425_));
 sg13g2_xnor2_1 _3164_ (.Y(_0426_),
    .A(_1416_),
    .B(_1854_));
 sg13g2_a21oi_1 _3165_ (.A1(_0426_),
    .A2(_1894_),
    .Y(_0427_),
    .B1(net44));
 sg13g2_o21ai_1 _3166_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0170_),
    .A2(_0195_));
 sg13g2_xnor2_1 _3167_ (.Y(_0429_),
    .A(_1700_),
    .B(net45));
 sg13g2_xnor2_1 _3168_ (.Y(_0430_),
    .A(net62),
    .B(_1701_));
 sg13g2_a21oi_1 _3169_ (.A1(_0429_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(_0293_));
 sg13g2_o21ai_1 _3170_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0429_),
    .A2(_0430_));
 sg13g2_buf_1 _3171_ (.A(_0303_),
    .X(_0433_));
 sg13g2_a221oi_1 _3172_ (.B2(_0432_),
    .C1(net34),
    .B1(_0428_),
    .A1(net46),
    .Y(_0434_),
    .A2(_0425_));
 sg13g2_nor3_1 _3173_ (.A(net37),
    .B(_0423_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_nor2_1 _3174_ (.A(_0421_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_inv_1 _3175_ (.Y(_0437_),
    .A(_0246_));
 sg13g2_nor2_1 _3176_ (.A(_0311_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_nand2_1 _3177_ (.Y(_0439_),
    .A(_0438_),
    .B(_0323_));
 sg13g2_o21ai_1 _3178_ (.B1(_0375_),
    .Y(_0440_),
    .A1(_0436_),
    .A2(_0439_));
 sg13g2_inv_1 _3179_ (.Y(_0441_),
    .A(_0338_));
 sg13g2_nor3_1 _3180_ (.A(_0331_),
    .B(_0441_),
    .C(_0371_),
    .Y(_0442_));
 sg13g2_nor2_1 _3181_ (.A(_0440_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_o21ai_1 _3182_ (.B1(_0443_),
    .Y(_0444_),
    .A1(_0418_),
    .A2(_0419_));
 sg13g2_nor2_1 _3183_ (.A(_0416_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_nand2b_1 _3184_ (.Y(_0446_),
    .B(_0445_),
    .A_N(_0412_));
 sg13g2_nor2_1 _3185_ (.A(_0379_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_nor3_1 _3186_ (.A(_0311_),
    .B(_0325_),
    .C(_0437_),
    .Y(_0448_));
 sg13g2_xor2_1 _3187_ (.B(_1799_),
    .A(_1798_),
    .X(_0449_));
 sg13g2_xor2_1 _3188_ (.B(_1852_),
    .A(_1856_),
    .X(_0450_));
 sg13g2_xor2_1 _3189_ (.B(_0450_),
    .A(_0449_),
    .X(_0451_));
 sg13g2_nand2_1 _3190_ (.Y(_0452_),
    .A(_1352_),
    .B(_0035_));
 sg13g2_a21oi_1 _3191_ (.A1(net53),
    .A2(_0034_),
    .Y(_0453_),
    .B1(net76));
 sg13g2_nand2_1 _3192_ (.Y(_0454_),
    .A(net53),
    .B(_0045_));
 sg13g2_o21ai_1 _3193_ (.B1(_0454_),
    .Y(_0455_),
    .A1(net53),
    .A2(_1510_));
 sg13g2_inv_1 _3194_ (.Y(_0456_),
    .A(_0455_));
 sg13g2_a22oi_1 _3195_ (.Y(_0457_),
    .B1(net76),
    .B2(_0456_),
    .A2(_0453_),
    .A1(_0452_));
 sg13g2_buf_1 _3196_ (.A(_0457_),
    .X(_0458_));
 sg13g2_xnor2_1 _3197_ (.Y(_0459_),
    .A(_1460_),
    .B(net41));
 sg13g2_inv_1 _3198_ (.Y(_0460_),
    .A(_0459_));
 sg13g2_a21oi_1 _3199_ (.A1(_0460_),
    .A2(_1894_),
    .Y(_0461_),
    .B1(net44));
 sg13g2_o21ai_1 _3200_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0170_),
    .A2(_0458_));
 sg13g2_o21ai_1 _3201_ (.B1(_0462_),
    .Y(_0463_),
    .A1(net39),
    .A2(_0451_));
 sg13g2_inv_1 _3202_ (.Y(_0464_),
    .A(_1851_));
 sg13g2_nor2_1 _3203_ (.A(_0035_),
    .B(_0168_),
    .Y(_0465_));
 sg13g2_a21oi_1 _3204_ (.A1(_0464_),
    .A2(_0465_),
    .Y(_0466_),
    .B1(net34));
 sg13g2_nand2_1 _3205_ (.Y(_0467_),
    .A(_0463_),
    .B(_0466_));
 sg13g2_buf_1 _3206_ (.A(_0361_),
    .X(_0468_));
 sg13g2_buf_1 _3207_ (.A(_0363_),
    .X(_0469_));
 sg13g2_a21oi_1 _3208_ (.A1(net23),
    .A2(_0464_),
    .Y(_0470_),
    .B1(net33));
 sg13g2_o21ai_1 _3209_ (.B1(_0470_),
    .Y(_0471_),
    .A1(_0464_),
    .A2(net23));
 sg13g2_nand3_1 _3210_ (.B(net38),
    .C(_0471_),
    .A(_0467_),
    .Y(_0472_));
 sg13g2_buf_1 _3211_ (.A(net37),
    .X(_0473_));
 sg13g2_a21oi_1 _3212_ (.A1(_0464_),
    .A2(net32),
    .Y(_0474_),
    .B1(net29));
 sg13g2_nand2_1 _3213_ (.Y(_0475_),
    .A(_0472_),
    .B(_0474_));
 sg13g2_a21oi_1 _3214_ (.A1(_0448_),
    .A2(_0475_),
    .Y(_0476_),
    .B1(_0328_));
 sg13g2_o21ai_1 _3215_ (.B1(_0476_),
    .Y(_0477_),
    .A1(_0441_),
    .A2(_0408_));
 sg13g2_nand2_1 _3216_ (.Y(_0478_),
    .A(_0264_),
    .B(_0410_));
 sg13g2_nand2_1 _3217_ (.Y(_0479_),
    .A(_0413_),
    .B(_0415_));
 sg13g2_o21ai_1 _3218_ (.B1(_0316_),
    .Y(_0480_),
    .A1(_0270_),
    .A2(_0479_));
 sg13g2_nand3b_1 _3219_ (.B(_0478_),
    .C(_0480_),
    .Y(_0481_),
    .A_N(_0477_));
 sg13g2_nand2_1 _3220_ (.Y(_0482_),
    .A(_0409_),
    .B(_0319_));
 sg13g2_nand2_1 _3221_ (.Y(_0483_),
    .A(_0482_),
    .B(net26));
 sg13g2_nand2_1 _3222_ (.Y(_0484_),
    .A(_0316_),
    .B(_0270_));
 sg13g2_nor2_1 _3223_ (.A(_0415_),
    .B(_0333_),
    .Y(_0485_));
 sg13g2_nor2_1 _3224_ (.A(_0325_),
    .B(_0333_),
    .Y(_0486_));
 sg13g2_nor2_1 _3225_ (.A(_0485_),
    .B(_0486_),
    .Y(_0487_));
 sg13g2_nand2_1 _3226_ (.Y(_0488_),
    .A(_0487_),
    .B(_0441_));
 sg13g2_nand3_1 _3227_ (.B(_0407_),
    .C(_0488_),
    .A(_0406_),
    .Y(_0489_));
 sg13g2_nand3_1 _3228_ (.B(_0484_),
    .C(_0489_),
    .A(_0411_),
    .Y(_0490_));
 sg13g2_nor2_1 _3229_ (.A(_0483_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_nor3_1 _3230_ (.A(_0377_),
    .B(_0481_),
    .C(_0491_),
    .Y(_0492_));
 sg13g2_inv_1 _3231_ (.Y(_0493_),
    .A(_0491_));
 sg13g2_nand2_1 _3232_ (.Y(_0494_),
    .A(_0481_),
    .B(_0378_));
 sg13g2_nor2_1 _3233_ (.A(_0493_),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_inv_1 _3234_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_o21ai_1 _3235_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0447_),
    .A2(_0492_));
 sg13g2_nand2_1 _3236_ (.Y(_0498_),
    .A(_1802_),
    .B(_1803_));
 sg13g2_nand2_1 _3237_ (.Y(_0499_),
    .A(_0498_),
    .B(_1786_));
 sg13g2_xnor2_1 _3238_ (.Y(_0500_),
    .A(_1787_),
    .B(_0499_));
 sg13g2_xnor2_1 _3239_ (.Y(_0501_),
    .A(_1874_),
    .B(_1861_));
 sg13g2_xnor2_1 _3240_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_nor2_1 _3241_ (.A(net76),
    .B(_0455_),
    .Y(_0503_));
 sg13g2_a21o_1 _3242_ (.A2(_0387_),
    .A1(net76),
    .B1(_0503_),
    .X(_0504_));
 sg13g2_buf_1 _3243_ (.A(_0504_),
    .X(_0505_));
 sg13g2_inv_1 _3244_ (.Y(_0506_),
    .A(_0505_));
 sg13g2_xnor2_1 _3245_ (.Y(_0507_),
    .A(_1422_),
    .B(net28));
 sg13g2_inv_1 _3246_ (.Y(_0508_),
    .A(_0507_));
 sg13g2_a21oi_1 _3247_ (.A1(_0508_),
    .A2(_1894_),
    .Y(_0509_),
    .B1(_1891_));
 sg13g2_o21ai_1 _3248_ (.B1(_0509_),
    .Y(_0510_),
    .A1(_0170_),
    .A2(_0506_));
 sg13g2_o21ai_1 _3249_ (.B1(_0510_),
    .Y(_0511_),
    .A1(net39),
    .A2(_0502_));
 sg13g2_nor2_1 _3250_ (.A(_1509_),
    .B(_0168_),
    .Y(_0512_));
 sg13g2_a21oi_1 _3251_ (.A1(_1878_),
    .A2(_0512_),
    .Y(_0513_),
    .B1(net34));
 sg13g2_nand2_1 _3252_ (.Y(_0514_),
    .A(_0511_),
    .B(_0513_));
 sg13g2_a21oi_1 _3253_ (.A1(_0362_),
    .A2(net28),
    .Y(_0515_),
    .B1(_0469_));
 sg13g2_o21ai_1 _3254_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_1873_),
    .A2(_0362_));
 sg13g2_nand3_1 _3255_ (.B(net38),
    .C(_0516_),
    .A(_0514_),
    .Y(_0517_));
 sg13g2_a21oi_1 _3256_ (.A1(_1878_),
    .A2(net32),
    .Y(_0518_),
    .B1(net29));
 sg13g2_a21oi_1 _3257_ (.A1(_0517_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(_0437_));
 sg13g2_inv_1 _3258_ (.Y(_0520_),
    .A(_0334_));
 sg13g2_a21oi_1 _3259_ (.A1(_0018_),
    .A2(_1527_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_o21ai_1 _3260_ (.B1(_0521_),
    .Y(_0522_),
    .A1(net52),
    .A2(_0519_));
 sg13g2_nand2_1 _3261_ (.Y(_0523_),
    .A(_0522_),
    .B(net26));
 sg13g2_nor2_1 _3262_ (.A(_0336_),
    .B(_0418_),
    .Y(_0524_));
 sg13g2_inv_1 _3263_ (.Y(_0525_),
    .A(_0484_));
 sg13g2_nor2_1 _3264_ (.A(_0413_),
    .B(_0263_),
    .Y(_0526_));
 sg13g2_nor4_1 _3265_ (.A(_0523_),
    .B(_0524_),
    .C(_0525_),
    .D(_0526_),
    .Y(_0527_));
 sg13g2_nor2_1 _3266_ (.A(_0316_),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_nand2_1 _3267_ (.Y(_0529_),
    .A(_0528_),
    .B(net26));
 sg13g2_nand2_1 _3268_ (.Y(_0530_),
    .A(_0527_),
    .B(_0316_));
 sg13g2_nand2_1 _3269_ (.Y(_0531_),
    .A(_0529_),
    .B(_0530_));
 sg13g2_inv_1 _3270_ (.Y(_0532_),
    .A(_0531_));
 sg13g2_nor2_1 _3271_ (.A(net30),
    .B(_0264_),
    .Y(_0533_));
 sg13g2_nor2_2 _3272_ (.A(_0377_),
    .B(_0533_),
    .Y(_0534_));
 sg13g2_inv_1 _3273_ (.Y(_0535_),
    .A(_0410_));
 sg13g2_nor2_1 _3274_ (.A(_0535_),
    .B(_0418_),
    .Y(_0536_));
 sg13g2_and3_1 _3275_ (.X(_0537_),
    .A(_0250_),
    .B(_0338_),
    .C(_0261_));
 sg13g2_inv_1 _3276_ (.Y(_0538_),
    .A(_0270_));
 sg13g2_nor2_1 _3277_ (.A(_0538_),
    .B(_0263_),
    .Y(_0539_));
 sg13g2_xnor2_1 _3278_ (.Y(_0540_),
    .A(_1804_),
    .B(_1802_));
 sg13g2_xor2_1 _3279_ (.B(_1858_),
    .A(_1859_),
    .X(_0541_));
 sg13g2_xor2_1 _3280_ (.B(_0541_),
    .A(_0540_),
    .X(_0542_));
 sg13g2_inv_1 _3281_ (.Y(_0543_),
    .A(_0347_));
 sg13g2_nand2_1 _3282_ (.Y(_0544_),
    .A(_0193_),
    .B(net65));
 sg13g2_o21ai_1 _3283_ (.B1(_0544_),
    .Y(_0545_),
    .A1(net65),
    .A2(_0543_));
 sg13g2_buf_1 _3284_ (.A(_0545_),
    .X(_0546_));
 sg13g2_inv_1 _3285_ (.Y(_0547_),
    .A(_0546_));
 sg13g2_xnor2_1 _3286_ (.Y(_0548_),
    .A(net61),
    .B(_1846_));
 sg13g2_inv_1 _3287_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_a21oi_1 _3288_ (.A1(_0549_),
    .A2(_1894_),
    .Y(_0550_),
    .B1(net44));
 sg13g2_o21ai_1 _3289_ (.B1(_0550_),
    .Y(_0551_),
    .A1(_0170_),
    .A2(_0547_));
 sg13g2_o21ai_1 _3290_ (.B1(_0551_),
    .Y(_0552_),
    .A1(net39),
    .A2(_0542_));
 sg13g2_nor2_1 _3291_ (.A(_0034_),
    .B(_0168_),
    .Y(_0553_));
 sg13g2_a21oi_1 _3292_ (.A1(_0225_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(net34));
 sg13g2_nand2_1 _3293_ (.Y(_0555_),
    .A(_0552_),
    .B(_0554_));
 sg13g2_a21oi_1 _3294_ (.A1(net23),
    .A2(_0225_),
    .Y(_0556_),
    .B1(net33));
 sg13g2_o21ai_1 _3295_ (.B1(_0556_),
    .Y(_0557_),
    .A1(_0225_),
    .A2(_0468_));
 sg13g2_nor2b_1 _3296_ (.A(net32),
    .B_N(_0557_),
    .Y(_0558_));
 sg13g2_a221oi_1 _3297_ (.B2(_0558_),
    .C1(net29),
    .B1(_0555_),
    .A1(_0225_),
    .Y(_0559_),
    .A2(net32));
 sg13g2_o21ai_1 _3298_ (.B1(net47),
    .Y(_0560_),
    .A1(_0559_),
    .A2(_0437_));
 sg13g2_a21oi_1 _3299_ (.A1(_0019_),
    .A2(net52),
    .Y(_0561_),
    .B1(_0487_));
 sg13g2_a21oi_1 _3300_ (.A1(_0560_),
    .A2(_0561_),
    .Y(_0562_),
    .B1(_0329_));
 sg13g2_nand2_1 _3301_ (.Y(_0563_),
    .A(_0482_),
    .B(_0562_));
 sg13g2_nor4_2 _3302_ (.A(_0536_),
    .B(_0537_),
    .C(_0539_),
    .Y(_0564_),
    .D(_0563_));
 sg13g2_inv_1 _3303_ (.Y(_0565_),
    .A(_0533_));
 sg13g2_nor2_1 _3304_ (.A(_0565_),
    .B(_0564_),
    .Y(_0566_));
 sg13g2_a21oi_2 _3305_ (.B1(_0566_),
    .Y(_0567_),
    .A2(_0564_),
    .A1(_0534_));
 sg13g2_nand3_1 _3306_ (.B(_0532_),
    .C(_0567_),
    .A(_0497_),
    .Y(_0568_));
 sg13g2_a22oi_1 _3307_ (.Y(_0569_),
    .B1(_0530_),
    .B2(_0566_),
    .A2(net26),
    .A1(_0528_));
 sg13g2_nand2_1 _3308_ (.Y(_0570_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_nand2b_1 _3309_ (.Y(_0571_),
    .B(_0570_),
    .A_N(_0379_));
 sg13g2_nand3_1 _3310_ (.B(_0379_),
    .C(_0569_),
    .A(_0568_),
    .Y(_0572_));
 sg13g2_buf_2 _3311_ (.A(_0572_),
    .X(_0573_));
 sg13g2_nand2_2 _3312_ (.Y(_0574_),
    .A(_0571_),
    .B(_0573_));
 sg13g2_nand3b_1 _3313_ (.B(_0493_),
    .C(_0378_),
    .Y(_0575_),
    .A_N(_0481_));
 sg13g2_inv_1 _3314_ (.Y(_0576_),
    .A(_0447_));
 sg13g2_a21oi_1 _3315_ (.A1(_0575_),
    .A2(_0576_),
    .Y(_0577_),
    .B1(_0495_));
 sg13g2_nand2b_1 _3316_ (.Y(_0578_),
    .B(_0577_),
    .A_N(_0567_));
 sg13g2_nand2_1 _3317_ (.Y(_0579_),
    .A(_0497_),
    .B(_0567_));
 sg13g2_nand3_1 _3318_ (.B(_0579_),
    .C(_1744_),
    .A(_0578_),
    .Y(_0580_));
 sg13g2_nor2_1 _3319_ (.A(_0495_),
    .B(_0492_),
    .Y(_0581_));
 sg13g2_nand2_1 _3320_ (.Y(_0582_),
    .A(_0581_),
    .B(\lfsr[9] ));
 sg13g2_nand2b_1 _3321_ (.Y(_0583_),
    .B(_0446_),
    .A_N(_0374_));
 sg13g2_a21oi_1 _3322_ (.A1(_0583_),
    .A2(\lfsr[8] ),
    .Y(_0584_),
    .B1(_0447_));
 sg13g2_nand2_1 _3323_ (.Y(_0585_),
    .A(_0581_),
    .B(_0576_));
 sg13g2_o21ai_1 _3324_ (.B1(\lfsr[9] ),
    .Y(_0586_),
    .A1(_0495_),
    .A2(_0492_));
 sg13g2_a22oi_1 _3325_ (.Y(_0587_),
    .B1(_0585_),
    .B2(_0586_),
    .A2(_0584_),
    .A1(_0582_));
 sg13g2_nand2_1 _3326_ (.Y(_0588_),
    .A(_0580_),
    .B(_0587_));
 sg13g2_nand2_1 _3327_ (.Y(_0589_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_nand2_1 _3328_ (.Y(_0590_),
    .A(_0589_),
    .B(\lfsr[10] ));
 sg13g2_nand2_1 _3329_ (.Y(_0591_),
    .A(_0588_),
    .B(_0590_));
 sg13g2_inv_1 _3330_ (.Y(_0592_),
    .A(_0021_));
 sg13g2_nand2_1 _3331_ (.Y(_0593_),
    .A(_0591_),
    .B(_0592_));
 sg13g2_nand2_1 _3332_ (.Y(_0594_),
    .A(_0564_),
    .B(_0534_));
 sg13g2_o21ai_1 _3333_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0566_),
    .A2(_0497_));
 sg13g2_xnor2_1 _3334_ (.Y(_0596_),
    .A(_0532_),
    .B(_0595_));
 sg13g2_nand2_1 _3335_ (.Y(_0597_),
    .A(_0593_),
    .B(_0596_));
 sg13g2_nand4_1 _3336_ (.B(_0576_),
    .C(_0581_),
    .A(_0567_),
    .Y(_0598_),
    .D(_0583_));
 sg13g2_nand2b_1 _3337_ (.Y(_0599_),
    .B(_0570_),
    .A_N(_0598_));
 sg13g2_nand4_1 _3338_ (.B(_0599_),
    .C(_0021_),
    .A(_0588_),
    .Y(_0600_),
    .D(_0590_));
 sg13g2_nand2_1 _3339_ (.Y(_0601_),
    .A(_0597_),
    .B(_0600_));
 sg13g2_xor2_1 _3340_ (.B(_0601_),
    .A(_0574_),
    .X(net8));
 sg13g2_nand2_1 _3341_ (.Y(_0602_),
    .A(_0493_),
    .B(_0378_));
 sg13g2_xnor2_1 _3342_ (.Y(_0603_),
    .A(_0602_),
    .B(_0573_));
 sg13g2_inv_1 _3343_ (.Y(_0604_),
    .A(_0603_));
 sg13g2_a21oi_1 _3344_ (.A1(_0601_),
    .A2(_0574_),
    .Y(_0605_),
    .B1(_0604_));
 sg13g2_nand3_1 _3345_ (.B(_0574_),
    .C(_0604_),
    .A(_0601_),
    .Y(_0606_));
 sg13g2_nor2b_1 _3346_ (.A(_0605_),
    .B_N(_0606_),
    .Y(net9));
 sg13g2_nand2_1 _3347_ (.Y(_0607_),
    .A(_0573_),
    .B(_0602_));
 sg13g2_nand2_1 _3348_ (.Y(_0608_),
    .A(_0606_),
    .B(_0607_));
 sg13g2_nor2_1 _3349_ (.A(_0565_),
    .B(_0491_),
    .Y(_0609_));
 sg13g2_inv_1 _3350_ (.Y(_0610_),
    .A(_0534_));
 sg13g2_nor2_1 _3351_ (.A(_0610_),
    .B(_0493_),
    .Y(_0611_));
 sg13g2_nor2_1 _3352_ (.A(_0609_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_inv_1 _3353_ (.Y(_0613_),
    .A(_0612_));
 sg13g2_nand2_1 _3354_ (.Y(_0614_),
    .A(_0608_),
    .B(_0613_));
 sg13g2_nand3_1 _3355_ (.B(_0607_),
    .C(_0612_),
    .A(_0606_),
    .Y(_0615_));
 sg13g2_nand2_1 _3356_ (.Y(net10),
    .A(_0614_),
    .B(_0615_));
 sg13g2_nor2_1 _3357_ (.A(_0613_),
    .B(_0603_),
    .Y(_0616_));
 sg13g2_nand3_1 _3358_ (.B(_0574_),
    .C(_0616_),
    .A(_0601_),
    .Y(_0617_));
 sg13g2_inv_1 _3359_ (.Y(_0618_),
    .A(_0602_));
 sg13g2_o21ai_1 _3360_ (.B1(_0610_),
    .Y(_0619_),
    .A1(_0618_),
    .A2(_0573_));
 sg13g2_nand2_1 _3361_ (.Y(_0620_),
    .A(_0617_),
    .B(_0619_));
 sg13g2_xnor2_1 _3362_ (.Y(_0621_),
    .A(_0418_),
    .B(_0534_));
 sg13g2_nand2_1 _3363_ (.Y(_0622_),
    .A(_0620_),
    .B(_0621_));
 sg13g2_nand2_1 _3364_ (.Y(_0623_),
    .A(_0565_),
    .B(_0316_));
 sg13g2_nand2_1 _3365_ (.Y(net11),
    .A(_0622_),
    .B(_0623_));
 sg13g2_xnor2_1 _3366_ (.Y(_0624_),
    .A(_0022_),
    .B(_0220_));
 sg13g2_xnor2_1 _3367_ (.Y(_0625_),
    .A(_1688_),
    .B(_1783_));
 sg13g2_xnor2_1 _3368_ (.Y(_0626_),
    .A(_1709_),
    .B(_1826_));
 sg13g2_nand2b_1 _3369_ (.Y(_0627_),
    .B(_0626_),
    .A_N(_0625_));
 sg13g2_xnor2_1 _3370_ (.Y(_0628_),
    .A(_1693_),
    .B(net25));
 sg13g2_inv_1 _3371_ (.Y(_0629_),
    .A(_0628_));
 sg13g2_xnor2_1 _3372_ (.Y(_0630_),
    .A(net54),
    .B(net41));
 sg13g2_nor2_1 _3373_ (.A(_1724_),
    .B(net45),
    .Y(_0631_));
 sg13g2_nand2_1 _3374_ (.Y(_0632_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_o21ai_1 _3375_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_1862_),
    .A2(net41));
 sg13g2_xnor2_1 _3376_ (.Y(_0634_),
    .A(net72),
    .B(net36));
 sg13g2_nand2_1 _3377_ (.Y(_0635_),
    .A(_0633_),
    .B(_0634_));
 sg13g2_o21ai_1 _3378_ (.B1(_0635_),
    .Y(_0636_),
    .A1(_1828_),
    .A2(net36));
 sg13g2_inv_1 _3379_ (.Y(_0637_),
    .A(_1810_));
 sg13g2_xnor2_1 _3380_ (.Y(_0638_),
    .A(_0637_),
    .B(net28));
 sg13g2_nand2_1 _3381_ (.Y(_0639_),
    .A(_0636_),
    .B(_0638_));
 sg13g2_nor2_1 _3382_ (.A(_0629_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_nand2b_1 _3383_ (.Y(_0641_),
    .B(_0640_),
    .A_N(_0627_));
 sg13g2_inv_1 _3384_ (.Y(_0642_),
    .A(_0036_));
 sg13g2_nand2_1 _3385_ (.Y(_0643_),
    .A(_0397_),
    .B(_0642_));
 sg13g2_nand2b_1 _3386_ (.Y(_0644_),
    .B(_0183_),
    .A_N(_0023_));
 sg13g2_o21ai_1 _3387_ (.B1(_0644_),
    .Y(_0645_),
    .A1(_0643_),
    .A2(_0625_));
 sg13g2_nor2_1 _3388_ (.A(_1810_),
    .B(net28),
    .Y(_0646_));
 sg13g2_a22oi_1 _3389_ (.Y(_0647_),
    .B1(_0646_),
    .B2(_0628_),
    .A2(_0356_),
    .A1(_1753_));
 sg13g2_nor2_1 _3390_ (.A(_0647_),
    .B(_0627_),
    .Y(_0648_));
 sg13g2_nor2_1 _3391_ (.A(_0645_),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_nand2_1 _3392_ (.Y(_0650_),
    .A(_0641_),
    .B(_0649_));
 sg13g2_nand2b_1 _3393_ (.Y(_0651_),
    .B(_0650_),
    .A_N(_0624_));
 sg13g2_nand3_1 _3394_ (.B(_0624_),
    .C(_0649_),
    .A(_0641_),
    .Y(_0652_));
 sg13g2_nand2_1 _3395_ (.Y(_0653_),
    .A(_0651_),
    .B(_0652_));
 sg13g2_nor2_1 _3396_ (.A(net74),
    .B(\i_project.controller_0.t[10] ),
    .Y(_0654_));
 sg13g2_nand2_1 _3397_ (.Y(_0655_),
    .A(net74),
    .B(\i_project.controller_0.t[10] ));
 sg13g2_inv_1 _3398_ (.Y(_0656_),
    .A(_0655_));
 sg13g2_nor2_1 _3399_ (.A(_0654_),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_xnor2_1 _3400_ (.Y(_0658_),
    .A(net75),
    .B(_1687_));
 sg13g2_xnor2_1 _3401_ (.Y(_0659_),
    .A(net59),
    .B(_1693_));
 sg13g2_nand2_1 _3402_ (.Y(_0660_),
    .A(_1416_),
    .B(net55));
 sg13g2_xnor2_1 _3403_ (.Y(_0661_),
    .A(net63),
    .B(_1697_));
 sg13g2_nand2_1 _3404_ (.Y(_0662_),
    .A(net63),
    .B(net54));
 sg13g2_o21ai_1 _3405_ (.B1(_0662_),
    .Y(_0663_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_xor2_1 _3406_ (.B(net72),
    .A(_1419_),
    .X(_0664_));
 sg13g2_nand2_1 _3407_ (.Y(_0665_),
    .A(_0663_),
    .B(_0664_));
 sg13g2_o21ai_1 _3408_ (.B1(_0665_),
    .Y(_0666_),
    .A1(net61),
    .A2(_1690_));
 sg13g2_xor2_1 _3409_ (.B(net71),
    .A(net57),
    .X(_0667_));
 sg13g2_nand2_1 _3410_ (.Y(_0668_),
    .A(net57),
    .B(net71));
 sg13g2_inv_1 _3411_ (.Y(_0669_),
    .A(_0668_));
 sg13g2_a21oi_2 _3412_ (.B1(_0669_),
    .Y(_0670_),
    .A2(_0667_),
    .A1(_0666_));
 sg13g2_nand2_1 _3413_ (.Y(_0671_),
    .A(net59),
    .B(_1693_));
 sg13g2_o21ai_1 _3414_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0659_),
    .A2(_0670_));
 sg13g2_xor2_1 _3415_ (.B(_1709_),
    .A(net60),
    .X(_0673_));
 sg13g2_nand2_1 _3416_ (.Y(_0674_),
    .A(net60),
    .B(_1709_));
 sg13g2_inv_1 _3417_ (.Y(_0675_),
    .A(_0674_));
 sg13g2_a21oi_1 _3418_ (.A1(_0672_),
    .A2(_0673_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_nand2_1 _3419_ (.Y(_0677_),
    .A(net75),
    .B(_1687_));
 sg13g2_o21ai_1 _3420_ (.B1(_0677_),
    .Y(_0678_),
    .A1(_0658_),
    .A2(_0676_));
 sg13g2_xnor2_1 _3421_ (.Y(_0679_),
    .A(_0657_),
    .B(_0678_));
 sg13g2_xor2_1 _3422_ (.B(_0679_),
    .A(_0653_),
    .X(_0680_));
 sg13g2_o21ai_1 _3423_ (.B1(_0294_),
    .Y(_0681_),
    .A1(_0293_),
    .A2(_0680_));
 sg13g2_a21oi_1 _3424_ (.A1(_0179_),
    .A2(net49),
    .Y(_0682_),
    .B1(net43));
 sg13g2_nand2_1 _3425_ (.Y(_0683_),
    .A(_0681_),
    .B(_0682_));
 sg13g2_xnor2_1 _3426_ (.Y(_0684_),
    .A(_0178_),
    .B(net27));
 sg13g2_a21oi_1 _3427_ (.A1(_0684_),
    .A2(_0187_),
    .Y(_0685_),
    .B1(net48));
 sg13g2_nand2_1 _3428_ (.Y(_0686_),
    .A(_0683_),
    .B(_0685_));
 sg13g2_a21oi_1 _3429_ (.A1(_0177_),
    .A2(net42),
    .Y(_0687_),
    .B1(_0207_));
 sg13g2_nand2_1 _3430_ (.Y(_0688_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_nand2_1 _3431_ (.Y(_0689_),
    .A(_0688_),
    .B(_0309_));
 sg13g2_nand2_1 _3432_ (.Y(_0690_),
    .A(_0689_),
    .B(net47));
 sg13g2_nand3_1 _3433_ (.B(_0259_),
    .C(_0261_),
    .A(_0690_),
    .Y(_0691_));
 sg13g2_inv_1 _3434_ (.Y(_0692_),
    .A(_0673_));
 sg13g2_xnor2_1 _3435_ (.Y(_0693_),
    .A(_0692_),
    .B(_0672_));
 sg13g2_inv_2 _3436_ (.Y(_0694_),
    .A(_0626_));
 sg13g2_o21ai_1 _3437_ (.B1(_0647_),
    .Y(_0695_),
    .A1(_0629_),
    .A2(_0639_));
 sg13g2_xnor2_1 _3438_ (.Y(_0696_),
    .A(_0694_),
    .B(_0695_));
 sg13g2_xnor2_1 _3439_ (.Y(_0697_),
    .A(_0693_),
    .B(_0696_));
 sg13g2_nand2_1 _3440_ (.Y(_0698_),
    .A(_0697_),
    .B(_1891_));
 sg13g2_inv_1 _3441_ (.Y(_0699_),
    .A(_0392_));
 sg13g2_nand2_1 _3442_ (.Y(_0700_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_a21oi_1 _3443_ (.A1(_0352_),
    .A2(net46),
    .Y(_0701_),
    .B1(net40));
 sg13g2_nand2_1 _3444_ (.Y(_0702_),
    .A(_0700_),
    .B(_0701_));
 sg13g2_xnor2_1 _3445_ (.Y(_0703_),
    .A(_0350_),
    .B(net24));
 sg13g2_a21oi_1 _3446_ (.A1(_0703_),
    .A2(net40),
    .Y(_0704_),
    .B1(net37));
 sg13g2_nand2_1 _3447_ (.Y(_0705_),
    .A(_0702_),
    .B(_0704_));
 sg13g2_a21oi_1 _3448_ (.A1(_0349_),
    .A2(net37),
    .Y(_0706_),
    .B1(net29));
 sg13g2_nand2_1 _3449_ (.Y(_0707_),
    .A(_0705_),
    .B(_0706_));
 sg13g2_nand2_1 _3450_ (.Y(_0708_),
    .A(_0707_),
    .B(net22));
 sg13g2_nand2_1 _3451_ (.Y(_0709_),
    .A(_0708_),
    .B(_0249_));
 sg13g2_inv_1 _3452_ (.Y(_0710_),
    .A(_0709_));
 sg13g2_nor3_1 _3453_ (.A(_0331_),
    .B(_0339_),
    .C(_0710_),
    .Y(_0711_));
 sg13g2_nor2_1 _3454_ (.A(net30),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_o21ai_1 _3455_ (.B1(_0712_),
    .Y(_0713_),
    .A1(_0538_),
    .A2(_0691_));
 sg13g2_xor2_1 _3456_ (.B(\i_project.controller_0.t[11] ),
    .A(_1434_),
    .X(_0714_));
 sg13g2_nor3_1 _3457_ (.A(_0654_),
    .B(_0656_),
    .C(_0658_),
    .Y(_0715_));
 sg13g2_nand3b_1 _3458_ (.B(_0715_),
    .C(_0673_),
    .Y(_0716_),
    .A_N(_0659_));
 sg13g2_o21ai_1 _3459_ (.B1(_0674_),
    .Y(_0717_),
    .A1(_0671_),
    .A2(_0692_));
 sg13g2_o21ai_1 _3460_ (.B1(_0655_),
    .Y(_0718_),
    .A1(_0677_),
    .A2(_0654_));
 sg13g2_a21oi_1 _3461_ (.A1(_0717_),
    .A2(_0715_),
    .Y(_0719_),
    .B1(_0718_));
 sg13g2_o21ai_1 _3462_ (.B1(_0719_),
    .Y(_0720_),
    .A1(_0716_),
    .A2(_0670_));
 sg13g2_xnor2_1 _3463_ (.Y(_0721_),
    .A(_0714_),
    .B(_0720_));
 sg13g2_xnor2_1 _3464_ (.Y(_0722_),
    .A(_0240_),
    .B(_0721_));
 sg13g2_nor2_1 _3465_ (.A(_0625_),
    .B(_0624_),
    .Y(_0723_));
 sg13g2_nand2b_1 _3466_ (.Y(_0724_),
    .B(_0639_),
    .A_N(_0646_));
 sg13g2_nand4_1 _3467_ (.B(_0626_),
    .C(_0628_),
    .A(_0723_),
    .Y(_0725_),
    .D(_0724_));
 sg13g2_nand2_1 _3468_ (.Y(_0726_),
    .A(_0356_),
    .B(_1753_));
 sg13g2_o21ai_1 _3469_ (.B1(_0643_),
    .Y(_0727_),
    .A1(_0726_),
    .A2(_0694_));
 sg13g2_nand2_1 _3470_ (.Y(_0728_),
    .A(_0220_),
    .B(_0022_));
 sg13g2_nand2b_1 _3471_ (.Y(_0729_),
    .B(_0728_),
    .A_N(_0644_));
 sg13g2_o21ai_1 _3472_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0022_),
    .A2(_0220_));
 sg13g2_a21oi_1 _3473_ (.A1(_0723_),
    .A2(_0727_),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_nand2_1 _3474_ (.Y(_0732_),
    .A(_0725_),
    .B(_0731_));
 sg13g2_nand2_1 _3475_ (.Y(_0733_),
    .A(_0732_),
    .B(\i_project.controller_0.t[11] ));
 sg13g2_nand3_1 _3476_ (.B(_1715_),
    .C(_0731_),
    .A(_0725_),
    .Y(_0734_));
 sg13g2_nand2_1 _3477_ (.Y(_0735_),
    .A(_0733_),
    .B(_0734_));
 sg13g2_nand2b_1 _3478_ (.Y(_0736_),
    .B(_0735_),
    .A_N(_0722_));
 sg13g2_nand3_1 _3479_ (.B(_0734_),
    .C(_0722_),
    .A(_0733_),
    .Y(_0737_));
 sg13g2_nand3_1 _3480_ (.B(_0737_),
    .C(net44),
    .A(_0736_),
    .Y(_0738_));
 sg13g2_xnor2_1 _3481_ (.Y(_0739_),
    .A(_1451_),
    .B(_0240_));
 sg13g2_o21ai_1 _3482_ (.B1(_0293_),
    .Y(_0740_),
    .A1(_0165_),
    .A2(_0739_));
 sg13g2_nand2_1 _3483_ (.Y(_0741_),
    .A(_0738_),
    .B(_0740_));
 sg13g2_a21oi_1 _3484_ (.A1(_0276_),
    .A2(net46),
    .Y(_0742_),
    .B1(net40));
 sg13g2_nand2_1 _3485_ (.Y(_0743_),
    .A(_0741_),
    .B(_0742_));
 sg13g2_xnor2_1 _3486_ (.Y(_0744_),
    .A(_0291_),
    .B(net24));
 sg13g2_a21oi_1 _3487_ (.A1(_0744_),
    .A2(net40),
    .Y(_0745_),
    .B1(_0367_));
 sg13g2_nand2_1 _3488_ (.Y(_0746_),
    .A(_0743_),
    .B(_0745_));
 sg13g2_a21oi_1 _3489_ (.A1(_0292_),
    .A2(_0367_),
    .Y(_0747_),
    .B1(net29));
 sg13g2_nand2_1 _3490_ (.Y(_0748_),
    .A(_0746_),
    .B(_0747_));
 sg13g2_nand2_1 _3491_ (.Y(_0749_),
    .A(_0748_),
    .B(net22));
 sg13g2_nand2_1 _3492_ (.Y(_0750_),
    .A(_0749_),
    .B(net47));
 sg13g2_nand2_1 _3493_ (.Y(_0751_),
    .A(_0750_),
    .B(_0313_));
 sg13g2_buf_8 _3494_ (.A(_0751_),
    .X(_0752_));
 sg13g2_nand2_2 _3495_ (.Y(_0753_),
    .A(_0752_),
    .B(net30));
 sg13g2_nor2_1 _3496_ (.A(_0413_),
    .B(_0752_),
    .Y(_0754_));
 sg13g2_a21oi_2 _3497_ (.B1(_0754_),
    .Y(_0755_),
    .A2(_0753_),
    .A1(_0713_));
 sg13g2_nand3_1 _3498_ (.B(_0313_),
    .C(_0479_),
    .A(_0750_),
    .Y(_0756_));
 sg13g2_xor2_1 _3499_ (.B(_0663_),
    .A(_0664_),
    .X(_0757_));
 sg13g2_xor2_1 _3500_ (.B(_0633_),
    .A(_0634_),
    .X(_0758_));
 sg13g2_xor2_1 _3501_ (.B(_0758_),
    .A(_0757_),
    .X(_0759_));
 sg13g2_inv_1 _3502_ (.Y(_0760_),
    .A(_0550_));
 sg13g2_o21ai_1 _3503_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_0340_),
    .A2(_0759_));
 sg13g2_a21oi_1 _3504_ (.A1(_0460_),
    .A2(net46),
    .Y(_0762_),
    .B1(net34));
 sg13g2_nand2_1 _3505_ (.Y(_0763_),
    .A(_0761_),
    .B(_0762_));
 sg13g2_a21oi_1 _3506_ (.A1(_0362_),
    .A2(_0458_),
    .Y(_0764_),
    .B1(net33));
 sg13g2_o21ai_1 _3507_ (.B1(_0764_),
    .Y(_0765_),
    .A1(_0362_),
    .A2(_0458_));
 sg13g2_nand3_1 _3508_ (.B(_0360_),
    .C(_0765_),
    .A(_0763_),
    .Y(_0766_));
 sg13g2_nand2b_1 _3509_ (.Y(_0767_),
    .B(net32),
    .A_N(_0458_));
 sg13g2_nand3_1 _3510_ (.B(_0420_),
    .C(_0767_),
    .A(_0766_),
    .Y(_0768_));
 sg13g2_nand2_1 _3511_ (.Y(_0769_),
    .A(_0448_),
    .B(_0768_));
 sg13g2_nand2_1 _3512_ (.Y(_0770_),
    .A(_0756_),
    .B(_0769_));
 sg13g2_nand2_1 _3513_ (.Y(_0771_),
    .A(_0690_),
    .B(_0261_));
 sg13g2_nor2_1 _3514_ (.A(_0333_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_nand2_1 _3515_ (.Y(_0773_),
    .A(_0772_),
    .B(_0410_));
 sg13g2_nand2_1 _3516_ (.Y(_0774_),
    .A(_0773_),
    .B(net26));
 sg13g2_nor2_1 _3517_ (.A(_0770_),
    .B(_0774_),
    .Y(_0775_));
 sg13g2_nand3_1 _3518_ (.B(_0313_),
    .C(_0270_),
    .A(_0750_),
    .Y(_0776_));
 sg13g2_nand2_1 _3519_ (.Y(_0777_),
    .A(_0695_),
    .B(_0626_));
 sg13g2_xnor2_1 _3520_ (.Y(_0778_),
    .A(_0179_),
    .B(_0676_));
 sg13g2_a21oi_1 _3521_ (.A1(_0777_),
    .A2(_0643_),
    .Y(_0779_),
    .B1(_0778_));
 sg13g2_nand3_1 _3522_ (.B(_0778_),
    .C(_0643_),
    .A(_0777_),
    .Y(_0780_));
 sg13g2_nand2_1 _3523_ (.Y(_0781_),
    .A(_0780_),
    .B(net44));
 sg13g2_inv_1 _3524_ (.Y(_0782_),
    .A(_0180_));
 sg13g2_o21ai_1 _3525_ (.B1(_0782_),
    .Y(_0783_),
    .A1(_0779_),
    .A2(_0781_));
 sg13g2_a21oi_1 _3526_ (.A1(_0391_),
    .A2(net49),
    .Y(_0784_),
    .B1(net43));
 sg13g2_nand2_1 _3527_ (.Y(_0785_),
    .A(_0783_),
    .B(_0784_));
 sg13g2_xnor2_1 _3528_ (.Y(_0786_),
    .A(_0390_),
    .B(net27));
 sg13g2_a21oi_1 _3529_ (.A1(_0786_),
    .A2(net43),
    .Y(_0787_),
    .B1(_0203_));
 sg13g2_nand2_1 _3530_ (.Y(_0788_),
    .A(_0785_),
    .B(_0787_));
 sg13g2_a21oi_1 _3531_ (.A1(_0389_),
    .A2(net42),
    .Y(_0789_),
    .B1(net35));
 sg13g2_nand2_1 _3532_ (.Y(_0790_),
    .A(_0788_),
    .B(_0789_));
 sg13g2_nand2_1 _3533_ (.Y(_0791_),
    .A(_0790_),
    .B(_0246_));
 sg13g2_nand2_1 _3534_ (.Y(_0792_),
    .A(_0791_),
    .B(net47));
 sg13g2_nand2_1 _3535_ (.Y(_0793_),
    .A(_0792_),
    .B(_0407_));
 sg13g2_nor2_1 _3536_ (.A(_0333_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_nand2_1 _3537_ (.Y(_0795_),
    .A(_0794_),
    .B(_0335_));
 sg13g2_nand2_1 _3538_ (.Y(_0796_),
    .A(_0776_),
    .B(_0795_));
 sg13g2_inv_2 _3539_ (.Y(_0797_),
    .A(_0796_));
 sg13g2_nand2_1 _3540_ (.Y(_0798_),
    .A(_0775_),
    .B(_0797_));
 sg13g2_nor2_1 _3541_ (.A(_0520_),
    .B(_0793_),
    .Y(_0799_));
 sg13g2_nand2_1 _3542_ (.Y(_0800_),
    .A(_0794_),
    .B(_0319_));
 sg13g2_nand2_1 _3543_ (.Y(_0801_),
    .A(_0800_),
    .B(_0375_));
 sg13g2_nor2_1 _3544_ (.A(_0799_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_nand2_1 _3545_ (.Y(_0803_),
    .A(_0797_),
    .B(_0802_));
 sg13g2_nand2_2 _3546_ (.Y(_0804_),
    .A(_0803_),
    .B(_0753_));
 sg13g2_nor2_1 _3547_ (.A(_0798_),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_nor3_1 _3548_ (.A(_0333_),
    .B(_0535_),
    .C(_0793_),
    .Y(_0806_));
 sg13g2_nand3_1 _3549_ (.B(_0330_),
    .C(_0338_),
    .A(_0709_),
    .Y(_0807_));
 sg13g2_xnor2_1 _3550_ (.Y(_0808_),
    .A(_0195_),
    .B(_0468_));
 sg13g2_xor2_1 _3551_ (.B(_0661_),
    .A(_0660_),
    .X(_0809_));
 sg13g2_xor2_1 _3552_ (.B(_0630_),
    .A(_0631_),
    .X(_0810_));
 sg13g2_xor2_1 _3553_ (.B(_0810_),
    .A(_0809_),
    .X(_0811_));
 sg13g2_inv_1 _3554_ (.Y(_0812_),
    .A(_0461_));
 sg13g2_o21ai_1 _3555_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0340_),
    .A2(_0811_));
 sg13g2_a21oi_1 _3556_ (.A1(_0426_),
    .A2(_0424_),
    .Y(_0814_),
    .B1(_0433_));
 sg13g2_a221oi_1 _3557_ (.B2(_0814_),
    .C1(net32),
    .B1(_0813_),
    .A1(_0433_),
    .Y(_0815_),
    .A2(_0808_));
 sg13g2_nand2b_1 _3558_ (.Y(_0816_),
    .B(net32),
    .A_N(_0195_));
 sg13g2_nand2_1 _3559_ (.Y(_0817_),
    .A(_0816_),
    .B(_0420_));
 sg13g2_inv_1 _3560_ (.Y(_0818_),
    .A(_0439_));
 sg13g2_o21ai_1 _3561_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0815_),
    .A2(_0817_));
 sg13g2_nand2_1 _3562_ (.Y(_0820_),
    .A(_0807_),
    .B(_0819_));
 sg13g2_nor2_1 _3563_ (.A(_0806_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_inv_2 _3564_ (.Y(_0822_),
    .A(_0771_));
 sg13g2_nand2_1 _3565_ (.Y(_0823_),
    .A(_0822_),
    .B(_0485_));
 sg13g2_nand2_1 _3566_ (.Y(_0824_),
    .A(_0821_),
    .B(_0823_));
 sg13g2_nand2_1 _3567_ (.Y(_0825_),
    .A(_0772_),
    .B(_0319_));
 sg13g2_nor2b_1 _3568_ (.A(_0824_),
    .B_N(_0825_),
    .Y(_0826_));
 sg13g2_nor2_1 _3569_ (.A(_0538_),
    .B(_0691_),
    .Y(_0827_));
 sg13g2_nor2_1 _3570_ (.A(net30),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_inv_1 _3571_ (.Y(_0829_),
    .A(_0752_));
 sg13g2_nand2_1 _3572_ (.Y(_0830_),
    .A(_0829_),
    .B(_0324_));
 sg13g2_nand3_1 _3573_ (.B(_0828_),
    .C(_0830_),
    .A(_0826_),
    .Y(_0831_));
 sg13g2_nor2_1 _3574_ (.A(_0755_),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_nor2_1 _3575_ (.A(_0775_),
    .B(_0803_),
    .Y(_0833_));
 sg13g2_inv_1 _3576_ (.Y(_0834_),
    .A(_0833_));
 sg13g2_o21ai_1 _3577_ (.B1(_0834_),
    .Y(_0835_),
    .A1(_0805_),
    .A2(_0832_));
 sg13g2_inv_1 _3578_ (.Y(_0836_),
    .A(_0487_));
 sg13g2_a21oi_1 _3579_ (.A1(_0259_),
    .A2(_0321_),
    .Y(_0837_),
    .B1(_0836_));
 sg13g2_nand2b_1 _3580_ (.Y(_0838_),
    .B(_0822_),
    .A_N(_0837_));
 sg13g2_nand3_1 _3581_ (.B(_0838_),
    .C(net26),
    .A(_0773_),
    .Y(_0839_));
 sg13g2_nand2_2 _3582_ (.Y(_0840_),
    .A(_0839_),
    .B(_0753_));
 sg13g2_a21oi_1 _3583_ (.A1(_0535_),
    .A2(_0376_),
    .Y(_0841_),
    .B1(_0752_));
 sg13g2_nand2_1 _3584_ (.Y(_0842_),
    .A(_0822_),
    .B(_0338_));
 sg13g2_xor2_1 _3585_ (.B(_0666_),
    .A(_0667_),
    .X(_0843_));
 sg13g2_xnor2_1 _3586_ (.Y(_0844_),
    .A(_0638_),
    .B(_0636_));
 sg13g2_xnor2_1 _3587_ (.Y(_0845_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_inv_1 _3588_ (.Y(_0846_),
    .A(_0509_));
 sg13g2_o21ai_1 _3589_ (.B1(_0846_),
    .Y(_0847_),
    .A1(net39),
    .A2(_0845_));
 sg13g2_a21oi_1 _3590_ (.A1(_0549_),
    .A2(net46),
    .Y(_0848_),
    .B1(net34));
 sg13g2_nand2_1 _3591_ (.Y(_0849_),
    .A(_0847_),
    .B(_0848_));
 sg13g2_a21oi_1 _3592_ (.A1(_0361_),
    .A2(_0546_),
    .Y(_0850_),
    .B1(_0469_));
 sg13g2_o21ai_1 _3593_ (.B1(_0850_),
    .Y(_0851_),
    .A1(net23),
    .A2(_0546_));
 sg13g2_nand3_1 _3594_ (.B(net38),
    .C(_0851_),
    .A(_0849_),
    .Y(_0852_));
 sg13g2_a21oi_1 _3595_ (.A1(_0546_),
    .A2(_0473_),
    .Y(_0853_),
    .B1(_0368_));
 sg13g2_a21oi_1 _3596_ (.A1(_0852_),
    .A2(_0853_),
    .Y(_0854_),
    .B1(_0437_));
 sg13g2_nand2b_1 _3597_ (.Y(_0855_),
    .B(net47),
    .A_N(_0854_));
 sg13g2_nand2_1 _3598_ (.Y(_0856_),
    .A(_0855_),
    .B(_0561_));
 sg13g2_nand3_1 _3599_ (.B(_0800_),
    .C(_0856_),
    .A(_0842_),
    .Y(_0857_));
 sg13g2_nor3_1 _3600_ (.A(_0827_),
    .B(_0841_),
    .C(_0857_),
    .Y(_0858_));
 sg13g2_xnor2_1 _3601_ (.Y(_0859_),
    .A(_0840_),
    .B(_0858_));
 sg13g2_inv_2 _3602_ (.Y(_0860_),
    .A(_0859_));
 sg13g2_a21oi_1 _3603_ (.A1(net23),
    .A2(_0505_),
    .Y(_0861_),
    .B1(net33));
 sg13g2_o21ai_1 _3604_ (.B1(_0861_),
    .Y(_0862_),
    .A1(net23),
    .A2(_0505_));
 sg13g2_nand2_1 _3605_ (.Y(_0863_),
    .A(_0862_),
    .B(net38));
 sg13g2_xnor2_1 _3606_ (.Y(_0864_),
    .A(_0670_),
    .B(_0351_));
 sg13g2_a21oi_1 _3607_ (.A1(_0724_),
    .A2(_0864_),
    .Y(_0865_),
    .B1(net39));
 sg13g2_o21ai_1 _3608_ (.B1(_0865_),
    .Y(_0866_),
    .A1(_0724_),
    .A2(_0864_));
 sg13g2_inv_1 _3609_ (.Y(_0867_),
    .A(_0353_));
 sg13g2_a221oi_1 _3610_ (.B2(_0867_),
    .C1(net34),
    .B1(_0866_),
    .A1(_0424_),
    .Y(_0868_),
    .A2(_0508_));
 sg13g2_a21oi_1 _3611_ (.A1(_0505_),
    .A2(_0473_),
    .Y(_0869_),
    .B1(_0368_));
 sg13g2_o21ai_1 _3612_ (.B1(_0869_),
    .Y(_0870_),
    .A1(_0863_),
    .A2(_0868_));
 sg13g2_a21o_1 _3613_ (.A2(net22),
    .A1(_0870_),
    .B1(net52),
    .X(_0871_));
 sg13g2_a21oi_1 _3614_ (.A1(_0871_),
    .A2(_0521_),
    .Y(_0872_),
    .B1(net30));
 sg13g2_nand2_1 _3615_ (.Y(_0873_),
    .A(_0776_),
    .B(_0872_));
 sg13g2_o21ai_1 _3616_ (.B1(_0825_),
    .Y(_0874_),
    .A1(_0336_),
    .A2(_0752_));
 sg13g2_nor3_1 _3617_ (.A(_0752_),
    .B(_0873_),
    .C(_0874_),
    .Y(_0875_));
 sg13g2_nand2_1 _3618_ (.Y(_0876_),
    .A(_0752_),
    .B(_0376_));
 sg13g2_nor2_1 _3619_ (.A(_0873_),
    .B(_0874_),
    .Y(_0877_));
 sg13g2_nor2_1 _3620_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_nor2_1 _3621_ (.A(_0875_),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_nor2b_1 _3622_ (.A(_0860_),
    .B_N(_0879_),
    .Y(_0880_));
 sg13g2_nand2_1 _3623_ (.Y(_0881_),
    .A(_0835_),
    .B(_0880_));
 sg13g2_inv_1 _3624_ (.Y(_0882_),
    .A(_0840_));
 sg13g2_nor2_1 _3625_ (.A(_0858_),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_a21oi_1 _3626_ (.A1(_0879_),
    .A2(_0883_),
    .Y(_0884_),
    .B1(_0878_));
 sg13g2_nand2_1 _3627_ (.Y(_0885_),
    .A(_0881_),
    .B(_0884_));
 sg13g2_xor2_1 _3628_ (.B(_0885_),
    .A(_0755_),
    .X(_0886_));
 sg13g2_nor2_1 _3629_ (.A(_0833_),
    .B(_0805_),
    .Y(_0887_));
 sg13g2_inv_1 _3630_ (.Y(_0888_),
    .A(_0832_));
 sg13g2_inv_1 _3631_ (.Y(_0889_),
    .A(_0828_));
 sg13g2_nor3_1 _3632_ (.A(_0754_),
    .B(_0711_),
    .C(_0889_),
    .Y(_0890_));
 sg13g2_nand2_1 _3633_ (.Y(_0891_),
    .A(_0831_),
    .B(_0890_));
 sg13g2_nand4_1 _3634_ (.B(_0859_),
    .C(_0888_),
    .A(_0887_),
    .Y(_0892_),
    .D(_0891_));
 sg13g2_nand2b_1 _3635_ (.Y(_0893_),
    .B(_0885_),
    .A_N(_0892_));
 sg13g2_nand2_1 _3636_ (.Y(_0894_),
    .A(_0893_),
    .B(_1747_));
 sg13g2_a21oi_1 _3637_ (.A1(_0859_),
    .A2(_0833_),
    .Y(_0895_),
    .B1(_0883_));
 sg13g2_nand3_1 _3638_ (.B(_0859_),
    .C(_0888_),
    .A(_0887_),
    .Y(_0896_));
 sg13g2_nand2_1 _3639_ (.Y(_0897_),
    .A(_0895_),
    .B(_0896_));
 sg13g2_xnor2_1 _3640_ (.Y(_0898_),
    .A(_0879_),
    .B(_0897_));
 sg13g2_nand2_1 _3641_ (.Y(_0899_),
    .A(_0894_),
    .B(_0898_));
 sg13g2_o21ai_1 _3642_ (.B1(\lfsr[17] ),
    .Y(_0900_),
    .A1(_0833_),
    .A2(_0805_));
 sg13g2_nand2_1 _3643_ (.Y(_0901_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_nand2_1 _3644_ (.Y(_0902_),
    .A(_0900_),
    .B(_0901_));
 sg13g2_a21oi_1 _3645_ (.A1(_0891_),
    .A2(\lfsr[16] ),
    .Y(_0903_),
    .B1(_0832_));
 sg13g2_nand2_1 _3646_ (.Y(_0904_),
    .A(_0887_),
    .B(\lfsr[17] ));
 sg13g2_nand2_1 _3647_ (.Y(_0905_),
    .A(_0903_),
    .B(_0904_));
 sg13g2_nand2_1 _3648_ (.Y(_0906_),
    .A(_0902_),
    .B(_0905_));
 sg13g2_nand2_1 _3649_ (.Y(_0907_),
    .A(_0906_),
    .B(_1746_));
 sg13g2_xnor2_1 _3650_ (.Y(_0908_),
    .A(_0859_),
    .B(_0835_));
 sg13g2_nor2_1 _3651_ (.A(_1746_),
    .B(_0906_),
    .Y(_0909_));
 sg13g2_a21oi_1 _3652_ (.A1(_0907_),
    .A2(_0908_),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_nand2_1 _3653_ (.Y(_0911_),
    .A(_0899_),
    .B(_0910_));
 sg13g2_nand2b_1 _3654_ (.Y(_0912_),
    .B(_1747_),
    .A_N(_0898_));
 sg13g2_nand2_1 _3655_ (.Y(_0913_),
    .A(_0911_),
    .B(_0912_));
 sg13g2_xor2_1 _3656_ (.B(_0913_),
    .A(_0886_),
    .X(net14));
 sg13g2_nand3_1 _3657_ (.B(_0755_),
    .C(_0884_),
    .A(_0881_),
    .Y(_0914_));
 sg13g2_xnor2_1 _3658_ (.Y(_0915_),
    .A(_0804_),
    .B(_0914_));
 sg13g2_inv_1 _3659_ (.Y(_0916_),
    .A(_0915_));
 sg13g2_a21oi_1 _3660_ (.A1(_0913_),
    .A2(_0886_),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_nand3_1 _3661_ (.B(_0886_),
    .C(_0916_),
    .A(_0913_),
    .Y(_0918_));
 sg13g2_nor2b_1 _3662_ (.A(_0917_),
    .B_N(_0918_),
    .Y(net15));
 sg13g2_nand2_1 _3663_ (.Y(_0919_),
    .A(_0914_),
    .B(_0804_));
 sg13g2_nand2_1 _3664_ (.Y(_0920_),
    .A(_0918_),
    .B(_0919_));
 sg13g2_nor2_1 _3665_ (.A(_0803_),
    .B(_0840_),
    .Y(_0921_));
 sg13g2_nor2_1 _3666_ (.A(_0839_),
    .B(_0804_),
    .Y(_0922_));
 sg13g2_nor2_1 _3667_ (.A(_0921_),
    .B(_0922_),
    .Y(_0923_));
 sg13g2_inv_1 _3668_ (.Y(_0924_),
    .A(_0923_));
 sg13g2_nand2_1 _3669_ (.Y(_0925_),
    .A(_0920_),
    .B(_0924_));
 sg13g2_nand3_1 _3670_ (.B(_0919_),
    .C(_0923_),
    .A(_0918_),
    .Y(_0926_));
 sg13g2_nand2_1 _3671_ (.Y(net16),
    .A(_0925_),
    .B(_0926_));
 sg13g2_nor2_1 _3672_ (.A(_0924_),
    .B(_0915_),
    .Y(_0927_));
 sg13g2_nand3_1 _3673_ (.B(_0886_),
    .C(_0927_),
    .A(_0913_),
    .Y(_0928_));
 sg13g2_inv_1 _3674_ (.Y(_0929_),
    .A(_0804_));
 sg13g2_o21ai_1 _3675_ (.B1(_0840_),
    .Y(_0930_),
    .A1(_0929_),
    .A2(_0914_));
 sg13g2_nand2_1 _3676_ (.Y(_0931_),
    .A(_0928_),
    .B(_0930_));
 sg13g2_xnor2_1 _3677_ (.Y(_0932_),
    .A(_0829_),
    .B(_0840_));
 sg13g2_nand2_1 _3678_ (.Y(_0933_),
    .A(_0931_),
    .B(_0932_));
 sg13g2_nand2_1 _3679_ (.Y(_0934_),
    .A(_0839_),
    .B(_0829_));
 sg13g2_nand2_1 _3680_ (.Y(net17),
    .A(_0933_),
    .B(_0934_));
 sg13g2_nand2_1 _3681_ (.Y(_0935_),
    .A(_1783_),
    .B(_1810_));
 sg13g2_nand3_1 _3682_ (.B(_1781_),
    .C(_0637_),
    .A(_1779_),
    .Y(_0936_));
 sg13g2_nand2_1 _3683_ (.Y(_0937_),
    .A(_0935_),
    .B(_0936_));
 sg13g2_nand2_1 _3684_ (.Y(_0938_),
    .A(_0937_),
    .B(net75));
 sg13g2_o21ai_1 _3685_ (.B1(_0938_),
    .Y(_0939_),
    .A1(_1692_),
    .A2(_0183_));
 sg13g2_xnor2_1 _3686_ (.Y(_0940_),
    .A(_1752_),
    .B(_0939_));
 sg13g2_xnor2_1 _3687_ (.Y(_0941_),
    .A(_0277_),
    .B(_0940_));
 sg13g2_inv_1 _3688_ (.Y(_0942_),
    .A(_1828_));
 sg13g2_nand2_1 _3689_ (.Y(_0943_),
    .A(_1826_),
    .B(_0942_));
 sg13g2_nand2_1 _3690_ (.Y(_0944_),
    .A(_0397_),
    .B(_1828_));
 sg13g2_nand2_1 _3691_ (.Y(_0945_),
    .A(_0943_),
    .B(_0944_));
 sg13g2_nand2_1 _3692_ (.Y(_0946_),
    .A(_0945_),
    .B(_1579_));
 sg13g2_nand3_1 _3693_ (.B(_0944_),
    .C(_1428_),
    .A(_0943_),
    .Y(_0947_));
 sg13g2_nand2_1 _3694_ (.Y(_0948_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_nand2_1 _3695_ (.Y(_0949_),
    .A(_1835_),
    .B(_1862_));
 sg13g2_nand3_1 _3696_ (.B(_1834_),
    .C(_1863_),
    .A(_1833_),
    .Y(_0950_));
 sg13g2_nand2_1 _3697_ (.Y(_0951_),
    .A(_0949_),
    .B(_0950_));
 sg13g2_nand2_1 _3698_ (.Y(_0952_),
    .A(_0951_),
    .B(net59));
 sg13g2_nand2_1 _3699_ (.Y(_0953_),
    .A(_1835_),
    .B(_1698_));
 sg13g2_nand2_1 _3700_ (.Y(_0954_),
    .A(_0952_),
    .B(_0953_));
 sg13g2_inv_1 _3701_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_nand2_1 _3702_ (.Y(_0956_),
    .A(_0948_),
    .B(_0955_));
 sg13g2_nand3_1 _3703_ (.B(_0947_),
    .C(_0954_),
    .A(_0946_),
    .Y(_0957_));
 sg13g2_nand2_1 _3704_ (.Y(_0958_),
    .A(_0956_),
    .B(_0957_));
 sg13g2_inv_1 _3705_ (.Y(_0959_),
    .A(_0943_));
 sg13g2_a21oi_1 _3706_ (.A1(_0944_),
    .A2(_1428_),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_inv_1 _3707_ (.Y(_0961_),
    .A(_0960_));
 sg13g2_nand3_1 _3708_ (.B(_0936_),
    .C(_1425_),
    .A(_0935_),
    .Y(_0962_));
 sg13g2_nand3_1 _3709_ (.B(_0938_),
    .C(_0962_),
    .A(_0961_),
    .Y(_0963_));
 sg13g2_nand2_1 _3710_ (.Y(_0964_),
    .A(_0938_),
    .B(_0962_));
 sg13g2_nand2_1 _3711_ (.Y(_0965_),
    .A(_0964_),
    .B(_0960_));
 sg13g2_nand2_1 _3712_ (.Y(_0966_),
    .A(_0963_),
    .B(_0965_));
 sg13g2_nor2_1 _3713_ (.A(_0958_),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_inv_1 _3714_ (.Y(_0968_),
    .A(_0041_));
 sg13g2_nand2_1 _3715_ (.Y(_0969_),
    .A(_1878_),
    .B(_0968_));
 sg13g2_nand3_1 _3716_ (.B(_1877_),
    .C(_0041_),
    .A(_1876_),
    .Y(_0970_));
 sg13g2_nand2_1 _3717_ (.Y(_0971_),
    .A(_0969_),
    .B(_0970_));
 sg13g2_nand2_1 _3718_ (.Y(_0972_),
    .A(_0971_),
    .B(net57));
 sg13g2_nand3_1 _3719_ (.B(_0970_),
    .C(_1422_),
    .A(_0969_),
    .Y(_0973_));
 sg13g2_xnor2_1 _3720_ (.Y(_0974_),
    .A(_0042_),
    .B(net36));
 sg13g2_nand2_1 _3721_ (.Y(_0975_),
    .A(_0974_),
    .B(net58));
 sg13g2_nand2_1 _3722_ (.Y(_0976_),
    .A(net36),
    .B(net70));
 sg13g2_nand2_1 _3723_ (.Y(_0977_),
    .A(_0975_),
    .B(_0976_));
 sg13g2_nand3_1 _3724_ (.B(_0973_),
    .C(_0977_),
    .A(_0972_),
    .Y(_0978_));
 sg13g2_buf_1 _3725_ (.A(_0978_),
    .X(_0979_));
 sg13g2_inv_1 _3726_ (.Y(_0980_),
    .A(_0979_));
 sg13g2_nand3_1 _3727_ (.B(_0950_),
    .C(_1445_),
    .A(_0949_),
    .Y(_0981_));
 sg13g2_nand2_1 _3728_ (.Y(_0982_),
    .A(_0952_),
    .B(_0981_));
 sg13g2_nor2_1 _3729_ (.A(_1724_),
    .B(_1878_),
    .Y(_0983_));
 sg13g2_a21oi_1 _3730_ (.A1(_0971_),
    .A2(net57),
    .Y(_0984_),
    .B1(_0983_));
 sg13g2_nand2_1 _3731_ (.Y(_0985_),
    .A(_0982_),
    .B(_0984_));
 sg13g2_xnor2_1 _3732_ (.Y(_0986_),
    .A(_1445_),
    .B(_0951_));
 sg13g2_nand2b_1 _3733_ (.Y(_0987_),
    .B(_0972_),
    .A_N(_0983_));
 sg13g2_nand2_1 _3734_ (.Y(_0988_),
    .A(_0986_),
    .B(_0987_));
 sg13g2_inv_1 _3735_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_a21oi_1 _3736_ (.A1(_0980_),
    .A2(_0985_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_inv_1 _3737_ (.Y(_0991_),
    .A(_0990_));
 sg13g2_inv_1 _3738_ (.Y(_0992_),
    .A(_0965_));
 sg13g2_o21ai_1 _3739_ (.B1(_0963_),
    .Y(_0993_),
    .A1(_0957_),
    .A2(_0992_));
 sg13g2_a21oi_1 _3740_ (.A1(_0967_),
    .A2(_0991_),
    .Y(_0994_),
    .B1(_0993_));
 sg13g2_nand2_1 _3741_ (.Y(_0995_),
    .A(_1851_),
    .B(_0024_));
 sg13g2_inv_1 _3742_ (.Y(_0996_),
    .A(_0024_));
 sg13g2_nand3_1 _3743_ (.B(_1849_),
    .C(_0996_),
    .A(_1848_),
    .Y(_0997_));
 sg13g2_nand2_1 _3744_ (.Y(_0998_),
    .A(_0995_),
    .B(_0997_));
 sg13g2_nand2_1 _3745_ (.Y(_0999_),
    .A(_0998_),
    .B(_1414_));
 sg13g2_o21ai_1 _3746_ (.B1(_0999_),
    .Y(_1000_),
    .A1(_1719_),
    .A2(_0464_));
 sg13g2_xnor2_1 _3747_ (.Y(_1001_),
    .A(net61),
    .B(_0974_));
 sg13g2_nor2_1 _3748_ (.A(_1000_),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_nand3_1 _3749_ (.B(_0997_),
    .C(_1460_),
    .A(_0995_),
    .Y(_1003_));
 sg13g2_nand2_1 _3750_ (.Y(_1004_),
    .A(_0999_),
    .B(_1003_));
 sg13g2_nor2_1 _3751_ (.A(_1559_),
    .B(_1855_),
    .Y(_1005_));
 sg13g2_nand2_1 _3752_ (.Y(_1006_),
    .A(_1004_),
    .B(_1005_));
 sg13g2_nor2b_2 _3753_ (.A(_1720_),
    .B_N(_0426_),
    .Y(_1007_));
 sg13g2_nor2_1 _3754_ (.A(_1005_),
    .B(_1004_),
    .Y(_1008_));
 sg13g2_a21oi_1 _3755_ (.A1(_1006_),
    .A2(_1007_),
    .Y(_1009_),
    .B1(_1008_));
 sg13g2_nand2_1 _3756_ (.Y(_1010_),
    .A(_1001_),
    .B(_1000_));
 sg13g2_o21ai_1 _3757_ (.B1(_1010_),
    .Y(_1011_),
    .A1(_1002_),
    .A2(_1009_));
 sg13g2_nand2_1 _3758_ (.Y(_1012_),
    .A(_0972_),
    .B(_0973_));
 sg13g2_nand2b_1 _3759_ (.Y(_1013_),
    .B(_1012_),
    .A_N(_0977_));
 sg13g2_nand2_1 _3760_ (.Y(_1014_),
    .A(_1013_),
    .B(_0979_));
 sg13g2_nand2_1 _3761_ (.Y(_1015_),
    .A(_0988_),
    .B(_0985_));
 sg13g2_nor2_1 _3762_ (.A(_1014_),
    .B(_1015_),
    .Y(_1016_));
 sg13g2_nand3_1 _3763_ (.B(_1011_),
    .C(_1016_),
    .A(_0967_),
    .Y(_1017_));
 sg13g2_nand2_1 _3764_ (.Y(_1018_),
    .A(_0994_),
    .B(_1017_));
 sg13g2_nand2b_1 _3765_ (.Y(_1019_),
    .B(_1018_),
    .A_N(_0941_));
 sg13g2_nand3_1 _3766_ (.B(_1017_),
    .C(_0941_),
    .A(_0994_),
    .Y(_1020_));
 sg13g2_nand3_1 _3767_ (.B(_1020_),
    .C(net49),
    .A(_1019_),
    .Y(_1021_));
 sg13g2_nor2_1 _3768_ (.A(_1752_),
    .B(_1826_),
    .Y(_1022_));
 sg13g2_nor2_1 _3769_ (.A(_1810_),
    .B(net25),
    .Y(_1023_));
 sg13g2_inv_1 _3770_ (.Y(_1024_),
    .A(_1023_));
 sg13g2_xnor2_1 _3771_ (.Y(_1025_),
    .A(_1753_),
    .B(_0397_));
 sg13g2_nor2_1 _3772_ (.A(_1024_),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_xnor2_1 _3773_ (.Y(_1027_),
    .A(_1692_),
    .B(net25));
 sg13g2_nand2_1 _3774_ (.Y(_1028_),
    .A(net28),
    .B(_1828_));
 sg13g2_nor2_1 _3775_ (.A(_1862_),
    .B(net36),
    .Y(_1029_));
 sg13g2_nor2_1 _3776_ (.A(_1828_),
    .B(net28),
    .Y(_1030_));
 sg13g2_a21oi_1 _3777_ (.A1(_1028_),
    .A2(_1029_),
    .Y(_1031_),
    .B1(_1030_));
 sg13g2_nor3_1 _3778_ (.A(_1027_),
    .B(_1031_),
    .C(_1025_),
    .Y(_1032_));
 sg13g2_nor3_1 _3779_ (.A(_1022_),
    .B(_1026_),
    .C(_1032_),
    .Y(_1033_));
 sg13g2_nor2_1 _3780_ (.A(_1027_),
    .B(_1025_),
    .Y(_1034_));
 sg13g2_xnor2_1 _3781_ (.Y(_1035_),
    .A(net55),
    .B(net41));
 sg13g2_nor2_1 _3782_ (.A(_1730_),
    .B(net45),
    .Y(_1036_));
 sg13g2_nand2_1 _3783_ (.Y(_1037_),
    .A(_1035_),
    .B(_1036_));
 sg13g2_o21ai_1 _3784_ (.B1(_1037_),
    .Y(_1038_),
    .A1(_0041_),
    .A2(net41));
 sg13g2_buf_1 _3785_ (.A(_1038_),
    .X(_1039_));
 sg13g2_nand2b_1 _3786_ (.Y(_1040_),
    .B(_1028_),
    .A_N(_1030_));
 sg13g2_xnor2_1 _3787_ (.Y(_1041_),
    .A(net54),
    .B(net36));
 sg13g2_nor2b_1 _3788_ (.A(_1040_),
    .B_N(_1041_),
    .Y(_1042_));
 sg13g2_nand3_1 _3789_ (.B(_1039_),
    .C(_1042_),
    .A(_1034_),
    .Y(_1043_));
 sg13g2_xnor2_1 _3790_ (.Y(_1044_),
    .A(_0642_),
    .B(_1783_));
 sg13g2_xor2_1 _3791_ (.B(_1693_),
    .A(net75),
    .X(_1045_));
 sg13g2_nand2_1 _3792_ (.Y(_1046_),
    .A(net63),
    .B(net70));
 sg13g2_xnor2_1 _3793_ (.Y(_1047_),
    .A(_1419_),
    .B(_1695_));
 sg13g2_nand2_1 _3794_ (.Y(_1048_),
    .A(net58),
    .B(net55));
 sg13g2_o21ai_1 _3795_ (.B1(_1048_),
    .Y(_1049_),
    .A1(_1046_),
    .A2(_1047_));
 sg13g2_xnor2_1 _3796_ (.Y(_1050_),
    .A(_1430_),
    .B(net72));
 sg13g2_xor2_1 _3797_ (.B(_1697_),
    .A(_1421_),
    .X(_1051_));
 sg13g2_inv_1 _3798_ (.Y(_1052_),
    .A(_1051_));
 sg13g2_nor2_1 _3799_ (.A(_1050_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_nand2_1 _3800_ (.Y(_1054_),
    .A(net57),
    .B(net54));
 sg13g2_nand2_1 _3801_ (.Y(_1055_),
    .A(_1430_),
    .B(net72));
 sg13g2_o21ai_1 _3802_ (.B1(_1055_),
    .Y(_1056_),
    .A1(_1054_),
    .A2(_1050_));
 sg13g2_a21oi_1 _3803_ (.A1(_1049_),
    .A2(_1053_),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_nand2_1 _3804_ (.Y(_1058_),
    .A(_1416_),
    .B(_1701_));
 sg13g2_inv_1 _3805_ (.Y(_1059_),
    .A(_1058_));
 sg13g2_xnor2_1 _3806_ (.Y(_1060_),
    .A(net63),
    .B(net70));
 sg13g2_nor2_1 _3807_ (.A(_1060_),
    .B(_1047_),
    .Y(_1061_));
 sg13g2_nand3_1 _3808_ (.B(_1059_),
    .C(_1061_),
    .A(_1053_),
    .Y(_1062_));
 sg13g2_nand2_1 _3809_ (.Y(_1063_),
    .A(_1057_),
    .B(_1062_));
 sg13g2_xor2_1 _3810_ (.B(net71),
    .A(_1428_),
    .X(_1064_));
 sg13g2_nand2_1 _3811_ (.Y(_1065_),
    .A(_1063_),
    .B(_1064_));
 sg13g2_o21ai_1 _3812_ (.B1(_1065_),
    .Y(_1066_),
    .A1(_1579_),
    .A2(_1692_));
 sg13g2_xnor2_1 _3813_ (.Y(_1067_),
    .A(_1045_),
    .B(_1066_));
 sg13g2_xnor2_1 _3814_ (.Y(_1068_),
    .A(_1044_),
    .B(_1067_));
 sg13g2_a21oi_1 _3815_ (.A1(_1033_),
    .A2(_1043_),
    .Y(_1069_),
    .B1(_1068_));
 sg13g2_nand3_1 _3816_ (.B(_1033_),
    .C(_1043_),
    .A(_1068_),
    .Y(_1070_));
 sg13g2_nand3b_1 _3817_ (.B(net44),
    .C(_1070_),
    .Y(_1071_),
    .A_N(_1069_));
 sg13g2_a21oi_1 _3818_ (.A1(_1071_),
    .A2(_0782_),
    .Y(_1072_),
    .B1(_0186_));
 sg13g2_nand2_1 _3819_ (.Y(_1073_),
    .A(_1021_),
    .B(_1072_));
 sg13g2_xnor2_1 _3820_ (.Y(_1074_),
    .A(_1694_),
    .B(net27));
 sg13g2_a21oi_1 _3821_ (.A1(_1074_),
    .A2(net43),
    .Y(_1075_),
    .B1(net48));
 sg13g2_nand2_1 _3822_ (.Y(_1076_),
    .A(_1073_),
    .B(_1075_));
 sg13g2_a21oi_1 _3823_ (.A1(_1753_),
    .A2(net48),
    .Y(_1077_),
    .B1(net35));
 sg13g2_nand2_1 _3824_ (.Y(_1078_),
    .A(_1076_),
    .B(_1077_));
 sg13g2_nand2_1 _3825_ (.Y(_1079_),
    .A(_1078_),
    .B(_0246_));
 sg13g2_nand2_1 _3826_ (.Y(_1080_),
    .A(_1079_),
    .B(_0248_));
 sg13g2_nand2_2 _3827_ (.Y(_1081_),
    .A(_1080_),
    .B(_0313_));
 sg13g2_nand2_1 _3828_ (.Y(_1082_),
    .A(_1081_),
    .B(_0328_));
 sg13g2_inv_1 _3829_ (.Y(_1083_),
    .A(_1082_));
 sg13g2_nor2_1 _3830_ (.A(_1015_),
    .B(_0958_),
    .Y(_1084_));
 sg13g2_xnor2_1 _3831_ (.Y(_1085_),
    .A(_0977_),
    .B(_1012_));
 sg13g2_nand2_1 _3832_ (.Y(_1086_),
    .A(_1011_),
    .B(_1085_));
 sg13g2_nand2_1 _3833_ (.Y(_1087_),
    .A(_1086_),
    .B(_0979_));
 sg13g2_nand2_1 _3834_ (.Y(_1088_),
    .A(_1084_),
    .B(_1087_));
 sg13g2_inv_1 _3835_ (.Y(_1089_),
    .A(_0957_));
 sg13g2_a21oi_1 _3836_ (.A1(_0956_),
    .A2(_0989_),
    .Y(_1090_),
    .B1(_1089_));
 sg13g2_nand2_1 _3837_ (.Y(_1091_),
    .A(_1088_),
    .B(_1090_));
 sg13g2_inv_1 _3838_ (.Y(_1092_),
    .A(_0966_));
 sg13g2_nand2_1 _3839_ (.Y(_1093_),
    .A(_1091_),
    .B(_1092_));
 sg13g2_nand3_1 _3840_ (.B(_0966_),
    .C(_1090_),
    .A(_1088_),
    .Y(_1094_));
 sg13g2_nand3_1 _3841_ (.B(_1094_),
    .C(net49),
    .A(_1093_),
    .Y(_1095_));
 sg13g2_xor2_1 _3842_ (.B(_1063_),
    .A(_1064_),
    .X(_1096_));
 sg13g2_xnor2_1 _3843_ (.Y(_1097_),
    .A(_1096_),
    .B(_1025_));
 sg13g2_nand2_1 _3844_ (.Y(_1098_),
    .A(_1042_),
    .B(_1039_));
 sg13g2_nand2_1 _3845_ (.Y(_1099_),
    .A(_1098_),
    .B(_1031_));
 sg13g2_nand2b_1 _3846_ (.Y(_1100_),
    .B(_1099_),
    .A_N(_1027_));
 sg13g2_nand2_1 _3847_ (.Y(_1101_),
    .A(_1100_),
    .B(_1024_));
 sg13g2_nand2b_1 _3848_ (.Y(_1102_),
    .B(_1101_),
    .A_N(_1097_));
 sg13g2_nand3_1 _3849_ (.B(_1024_),
    .C(_1097_),
    .A(_1100_),
    .Y(_1103_));
 sg13g2_nand3_1 _3850_ (.B(_1103_),
    .C(_1890_),
    .A(_1102_),
    .Y(_1104_));
 sg13g2_a21oi_1 _3851_ (.A1(_1104_),
    .A2(_0699_),
    .Y(_1105_),
    .B1(_0186_));
 sg13g2_nand2_1 _3852_ (.Y(_1106_),
    .A(_1095_),
    .B(_1105_));
 sg13g2_xnor2_1 _3853_ (.Y(_1107_),
    .A(_1692_),
    .B(_0199_));
 sg13g2_a21oi_1 _3854_ (.A1(_1107_),
    .A2(_0186_),
    .Y(_1108_),
    .B1(_0202_));
 sg13g2_nand2_1 _3855_ (.Y(_1109_),
    .A(_1106_),
    .B(_1108_));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net80),
    .D(_0000_),
    .Q_N(_1979_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net81),
    .D(_0001_),
    .Q_N(_1980_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net82),
    .D(_0002_),
    .Q_N(_1978_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net83),
    .D(_0052_),
    .Q_N(_1981_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net84),
    .D(_0003_),
    .Q_N(_1977_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net85),
    .D(_0004_),
    .Q_N(_1976_),
    .Q(_0164_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _3856__80 (.L_HI(net80));
 sg13g2_buf_1 _3864_ (.A(net86),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3865_ (.A(net87),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3866_ (.A(net88),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3867_ (.A(net89),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3868_ (.A(net90),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3869_ (.A(net91),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3870_ (.A(net92),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3871_ (.A(net93),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3872_ (.A(hsync),
    .X(net12));
 sg13g2_buf_1 _3873_ (.A(\i_project.controller_0.vga_sync.o_vsync ),
    .X(net13));
 sg13g2_buf_1 _3874_ (.A(net78),
    .X(uio_out[6]));
 sg13g2_buf_1 _3875_ (.A(net79),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net94),
    .D(_0053_),
    .Q_N(_0050_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[10]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net95),
    .D(_0054_),
    .Q_N(_1975_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 \counter[11]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net96),
    .D(_0055_),
    .Q_N(_1974_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 \counter[12]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net97),
    .D(_0056_),
    .Q_N(_1973_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 \counter[13]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net98),
    .D(_0057_),
    .Q_N(_1972_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 \counter[14]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net99),
    .D(_0058_),
    .Q_N(_1971_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 \counter[15]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net100),
    .D(_0059_),
    .Q_N(_1970_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 \counter[16]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net101),
    .D(_0060_),
    .Q_N(_1969_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 \counter[17]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net102),
    .D(_0061_),
    .Q_N(_1968_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 \counter[18]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net103),
    .D(_0062_),
    .Q_N(_1967_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 \counter[19]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net104),
    .D(_0063_),
    .Q_N(_1966_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net105),
    .D(_0064_),
    .Q_N(_1965_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[20]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net106),
    .D(_0065_),
    .Q_N(_1964_),
    .Q(\counter[20] ));
 sg13g2_dfrbp_1 \counter[21]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net107),
    .D(_0066_),
    .Q_N(_1963_),
    .Q(\counter[21] ));
 sg13g2_dfrbp_1 \counter[22]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net108),
    .D(_0067_),
    .Q_N(_1962_),
    .Q(\counter[22] ));
 sg13g2_dfrbp_1 \counter[23]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net109),
    .D(_0068_),
    .Q_N(_1961_),
    .Q(\counter[23] ));
 sg13g2_dfrbp_1 \counter[24]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net110),
    .D(_0069_),
    .Q_N(_1960_),
    .Q(\counter[24] ));
 sg13g2_dfrbp_1 \counter[25]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net111),
    .D(_0070_),
    .Q_N(_1959_),
    .Q(\counter[25] ));
 sg13g2_dfrbp_1 \counter[26]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net112),
    .D(_0071_),
    .Q_N(_1958_),
    .Q(\counter[26] ));
 sg13g2_dfrbp_1 \counter[27]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net113),
    .D(_0072_),
    .Q_N(_1957_),
    .Q(\counter[27] ));
 sg13g2_dfrbp_1 \counter[28]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net114),
    .D(_0073_),
    .Q_N(_1956_),
    .Q(\counter[28] ));
 sg13g2_dfrbp_1 \counter[29]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net115),
    .D(_0074_),
    .Q_N(_1955_),
    .Q(\counter[29] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net116),
    .D(_0075_),
    .Q_N(_1954_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[30]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net117),
    .D(_0076_),
    .Q_N(_1953_),
    .Q(\counter[30] ));
 sg13g2_dfrbp_1 \counter[31]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net118),
    .D(_0077_),
    .Q_N(_1952_),
    .Q(\counter[31] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net119),
    .D(_0078_),
    .Q_N(_1951_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net120),
    .D(_0079_),
    .Q_N(_1950_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net121),
    .D(_0080_),
    .Q_N(_1949_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net122),
    .D(_0081_),
    .Q_N(_1948_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net123),
    .D(_0082_),
    .Q_N(_1947_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net124),
    .D(_0083_),
    .Q_N(_1946_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \counter[9]$_SDFF_PN0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net125),
    .D(_0084_),
    .Q_N(_1982_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 \depth[0]$_DFF_P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net126),
    .D(_0005_),
    .Q_N(_1983_),
    .Q(\depth[0] ));
 sg13g2_dfrbp_1 \depth[1]$_DFF_P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net127),
    .D(_0006_),
    .Q_N(_1984_),
    .Q(\depth[1] ));
 sg13g2_dfrbp_1 \depth[2]$_DFF_P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net128),
    .D(_0007_),
    .Q_N(_0043_),
    .Q(\depth[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[2]$_DFFE_PN_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net129),
    .D(_0003_),
    .Q_N(_1945_),
    .Q(\i_project.controller_0.divider[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[3]$_DFFE_PN_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net130),
    .D(_0004_),
    .Q_N(_1944_),
    .Q(\i_project.controller_0.divider[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[4]$_DFFE_PN_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net131),
    .D(_0085_),
    .Q_N(_1943_),
    .Q(\i_project.controller_0.mode[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[5]$_DFFE_PN_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net132),
    .D(_0086_),
    .Q_N(_1942_),
    .Q(\i_project.controller_0.mode[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[6]$_DFFE_PN_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net133),
    .D(_0087_),
    .Q_N(_0029_),
    .Q(\i_project.controller_0.mode[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[7]$_DFFE_PN_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net134),
    .D(_0088_),
    .Q_N(_0027_),
    .Q(\i_project.controller_0.vga_sync.mode ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[0]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net135),
    .D(_0089_),
    .Q_N(_0051_),
    .Q(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[10]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net136),
    .D(_0090_),
    .Q_N(_0022_),
    .Q(\i_project.controller_0.t[10] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[11]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net137),
    .D(_0091_),
    .Q_N(_1941_),
    .Q(\i_project.controller_0.t[11] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[1]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net138),
    .D(_0092_),
    .Q_N(_0024_),
    .Q(\i_project.controller_0.mode_ramp_base[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[2]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net139),
    .D(_0093_),
    .Q_N(_0042_),
    .Q(\i_project.controller_0.mode_ramp_base[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[3]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net140),
    .D(_0094_),
    .Q_N(_0041_),
    .Q(\i_project.controller_0.mode_ramp_base[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[4]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net141),
    .D(_0095_),
    .Q_N(_0040_),
    .Q(\i_project.controller_0.mode_ramp_base[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[5]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net142),
    .D(_0096_),
    .Q_N(_0039_),
    .Q(\i_project.controller_0.mode_ramp_base[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[6]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_0097_),
    .Q_N(_0038_),
    .Q(\i_project.controller_0.mode_ramp_base[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[7]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net144),
    .D(_0098_),
    .Q_N(_0037_),
    .Q(\i_project.controller_0.mode_ramp_base[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[8]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net145),
    .D(_0099_),
    .Q_N(_0036_),
    .Q(\i_project.controller_0.t[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[9]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net146),
    .D(_0100_),
    .Q_N(_0023_),
    .Q(\i_project.controller_0.t[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net147),
    .D(_0101_),
    .Q_N(_0049_),
    .Q(\i_project.controller_0.h[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net148),
    .D(_0102_),
    .Q_N(_0035_),
    .Q(\i_project.controller_0.h[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net149),
    .D(_0103_),
    .Q_N(_0034_),
    .Q(\i_project.controller_0.h[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net150),
    .D(_0104_),
    .Q_N(_0025_),
    .Q(\i_project.controller_0.h[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net151),
    .D(_0105_),
    .Q_N(_0045_),
    .Q(\i_project.controller_0.h[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net152),
    .D(_0106_),
    .Q_N(_0046_),
    .Q(\i_project.controller_0.h[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net153),
    .D(_0107_),
    .Q_N(_0047_),
    .Q(\i_project.controller_0.h[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net154),
    .D(_0108_),
    .Q_N(_0028_),
    .Q(\i_project.controller_0.h[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net155),
    .D(_0109_),
    .Q_N(_0026_),
    .Q(\i_project.controller_0.h[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net156),
    .D(_0110_),
    .Q_N(_0017_),
    .Q(\i_project.controller_0.h[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hsync$_DFFE_PP_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net157),
    .D(_0111_),
    .Q_N(hsync),
    .Q(\i_project.controller_0.vga_sync.hsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net158),
    .D(_0112_),
    .Q_N(_1940_),
    .Q(\i_project.controller_0.v[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net159),
    .D(_0113_),
    .Q_N(_1939_),
    .Q(\i_project.controller_0.v[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net160),
    .D(_0114_),
    .Q_N(_1938_),
    .Q(\i_project.controller_0.v[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net161),
    .D(_0115_),
    .Q_N(_1937_),
    .Q(\i_project.controller_0.v[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net162),
    .D(_0116_),
    .Q_N(_1936_),
    .Q(\i_project.controller_0.v[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net163),
    .D(_0117_),
    .Q_N(_0031_),
    .Q(\i_project.controller_0.v[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net164),
    .D(_0118_),
    .Q_N(_1935_),
    .Q(\i_project.controller_0.v[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net165),
    .D(_0119_),
    .Q_N(_1934_),
    .Q(\i_project.controller_0.v[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net166),
    .D(_0120_),
    .Q_N(_0032_),
    .Q(\i_project.controller_0.v[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net167),
    .D(_0121_),
    .Q_N(_0030_),
    .Q(\i_project.controller_0.v[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vsync$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net168),
    .D(_0122_),
    .Q_N(_1933_),
    .Q(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[0]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net169),
    .D(_0123_),
    .Q_N(_1932_),
    .Q(\i_project.controller_0.voffset[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[1]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net170),
    .D(_0124_),
    .Q_N(_1931_),
    .Q(\i_project.controller_0.voffset[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[2]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net171),
    .D(_0125_),
    .Q_N(_1930_),
    .Q(\i_project.controller_0.voffset[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[3]$_SDFFCE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net172),
    .D(_0126_),
    .Q_N(_1929_),
    .Q(\i_project.controller_0.voffset[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[4]$_SDFFCE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net173),
    .D(_0127_),
    .Q_N(_1928_),
    .Q(\i_project.controller_0.voffset[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[5]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net174),
    .D(_0128_),
    .Q_N(_1927_),
    .Q(\i_project.controller_0.voffset[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[6]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net175),
    .D(_0129_),
    .Q_N(_1926_),
    .Q(\i_project.controller_0.voffset[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[7]$_SDFFCE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net176),
    .D(_0130_),
    .Q_N(_1925_),
    .Q(\i_project.controller_0.voffset[7] ));
 sg13g2_dfrbp_1 \lfsr[0]$_SDFF_PN1_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net177),
    .D(_0131_),
    .Q_N(_1924_),
    .Q(\lfsr[0] ));
 sg13g2_dfrbp_1 \lfsr[10]$_SDFF_PN1_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net178),
    .D(_0132_),
    .Q_N(_1923_),
    .Q(\lfsr[10] ));
 sg13g2_dfrbp_1 \lfsr[11]$_SDFF_PN1_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net179),
    .D(_0133_),
    .Q_N(_0021_),
    .Q(\lfsr[11] ));
 sg13g2_dfrbp_1 \lfsr[12]$_SDFF_PN1_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net180),
    .D(_0134_),
    .Q_N(_1922_),
    .Q(\lfsr[12] ));
 sg13g2_dfrbp_1 \lfsr[13]$_SDFF_PN1_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net181),
    .D(_0135_),
    .Q_N(_1921_),
    .Q(\lfsr[13] ));
 sg13g2_dfrbp_1 \lfsr[14]$_SDFF_PN1_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net182),
    .D(_0136_),
    .Q_N(_1920_),
    .Q(\lfsr[14] ));
 sg13g2_dfrbp_1 \lfsr[15]$_SDFF_PN1_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net183),
    .D(_0137_),
    .Q_N(_1919_),
    .Q(\lfsr[15] ));
 sg13g2_dfrbp_1 \lfsr[16]$_SDFF_PN1_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net184),
    .D(_0138_),
    .Q_N(_1918_),
    .Q(\lfsr[16] ));
 sg13g2_dfrbp_1 \lfsr[17]$_SDFF_PN1_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net185),
    .D(_0139_),
    .Q_N(_1917_),
    .Q(\lfsr[17] ));
 sg13g2_dfrbp_1 \lfsr[18]$_SDFF_PN1_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net186),
    .D(_0140_),
    .Q_N(_1916_),
    .Q(\lfsr[18] ));
 sg13g2_dfrbp_1 \lfsr[19]$_SDFF_PN1_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net187),
    .D(_0141_),
    .Q_N(_1915_),
    .Q(\lfsr[19] ));
 sg13g2_dfrbp_1 \lfsr[1]$_SDFF_PN1_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net188),
    .D(_0142_),
    .Q_N(_1914_),
    .Q(\lfsr[1] ));
 sg13g2_dfrbp_1 \lfsr[20]$_SDFF_PN1_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net189),
    .D(_0143_),
    .Q_N(_1913_),
    .Q(\lfsr[20] ));
 sg13g2_dfrbp_1 \lfsr[21]$_SDFF_PN1_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net190),
    .D(_0144_),
    .Q_N(_1912_),
    .Q(\lfsr[21] ));
 sg13g2_dfrbp_1 \lfsr[22]$_SDFF_PN1_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net191),
    .D(_0145_),
    .Q_N(_1911_),
    .Q(\lfsr[22] ));
 sg13g2_dfrbp_1 \lfsr[23]$_SDFF_PN1_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net192),
    .D(_0146_),
    .Q_N(_1910_),
    .Q(\lfsr[23] ));
 sg13g2_dfrbp_1 \lfsr[24]$_SDFF_PN1_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net193),
    .D(_0147_),
    .Q_N(_1909_),
    .Q(\lfsr[24] ));
 sg13g2_dfrbp_1 \lfsr[25]$_SDFF_PN1_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net194),
    .D(_0148_),
    .Q_N(_1908_),
    .Q(\lfsr[25] ));
 sg13g2_dfrbp_1 \lfsr[26]$_SDFF_PN1_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net195),
    .D(_0149_),
    .Q_N(_1907_),
    .Q(\lfsr[26] ));
 sg13g2_dfrbp_1 \lfsr[27]$_SDFF_PN1_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net196),
    .D(_0150_),
    .Q_N(_1906_),
    .Q(\lfsr[27] ));
 sg13g2_dfrbp_1 \lfsr[28]$_SDFF_PN1_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net197),
    .D(_0151_),
    .Q_N(_1905_),
    .Q(\lfsr[28] ));
 sg13g2_dfrbp_1 \lfsr[29]$_SDFF_PN1_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net198),
    .D(_0152_),
    .Q_N(_1904_),
    .Q(\lfsr[29] ));
 sg13g2_dfrbp_1 \lfsr[2]$_SDFF_PN1_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net199),
    .D(_0153_),
    .Q_N(_1903_),
    .Q(\lfsr[2] ));
 sg13g2_dfrbp_1 \lfsr[30]$_SDFF_PN1_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net200),
    .D(_0154_),
    .Q_N(_1902_),
    .Q(\lfsr[30] ));
 sg13g2_dfrbp_1 \lfsr[31]$_SDFF_PN1_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net201),
    .D(_0155_),
    .Q_N(_1901_),
    .Q(\lfsr[31] ));
 sg13g2_dfrbp_1 \lfsr[3]$_SDFF_PN1_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net202),
    .D(_0156_),
    .Q_N(_1900_),
    .Q(\lfsr[3] ));
 sg13g2_dfrbp_1 \lfsr[4]$_SDFF_PN1_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net203),
    .D(_0157_),
    .Q_N(_1899_),
    .Q(\lfsr[4] ));
 sg13g2_dfrbp_1 \lfsr[5]$_SDFF_PN1_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net204),
    .D(_0158_),
    .Q_N(_1898_),
    .Q(\lfsr[5] ));
 sg13g2_dfrbp_1 \lfsr[6]$_SDFF_PN1_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net205),
    .D(_0159_),
    .Q_N(_1897_),
    .Q(\lfsr[6] ));
 sg13g2_dfrbp_1 \lfsr[7]$_SDFF_PN1_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net206),
    .D(_0160_),
    .Q_N(_1896_),
    .Q(\lfsr[7] ));
 sg13g2_dfrbp_1 \lfsr[8]$_SDFF_PN1_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net207),
    .D(_0161_),
    .Q_N(_1895_),
    .Q(\lfsr[8] ));
 sg13g2_dfrbp_1 \lfsr[9]$_SDFF_PN1_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net208),
    .D(_0162_),
    .Q_N(_1985_),
    .Q(\lfsr[9] ));
 sg13g2_dfrbp_1 \project_rst_n$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net209),
    .D(_0008_),
    .Q_N(_1986_),
    .Q(\i_project.controller_0.rst_n ));
 sg13g2_dfrbp_1 \project_ui_in[2]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net210),
    .D(\counter[30] ),
    .Q_N(_0019_),
    .Q(\i_project.controller_0.grey_pass[10] ));
 sg13g2_dfrbp_1 \project_ui_in[3]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net211),
    .D(\counter[31] ),
    .Q_N(_0018_),
    .Q(\i_project.controller_0.grey_pass[11] ));
 sg13g2_dfrbp_1 \project_ui_in[4]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net212),
    .D(_0009_),
    .Q_N(_0044_),
    .Q(\i_project.controller_0.grey_pass[12] ));
 sg13g2_dfrbp_1 \project_ui_in[5]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net213),
    .D(_0010_),
    .Q_N(_0020_),
    .Q(\i_project.controller_0.grey_pass[13] ));
 sg13g2_dfrbp_1 \project_ui_in[6]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net214),
    .D(_0011_),
    .Q_N(_0048_),
    .Q(\i_project.controller_0.grey_pass[14] ));
 sg13g2_dfrbp_1 \project_ui_in[7]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net215),
    .D(_0163_),
    .Q_N(_0033_),
    .Q(\i_project.controller_0.grey_pass[15] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout22 (.A(_0309_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0468_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0361_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1836_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0376_),
    .X(net26));
 sg13g2_buf_4 fanout27 (.X(net27),
    .A(_0200_));
 sg13g2_buf_2 fanout28 (.A(_1873_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0368_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0329_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1569_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0473_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0469_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0433_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0207_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1846_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0367_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0360_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0340_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0303_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1851_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0304_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0187_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1891_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1855_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0424_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0249_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0203_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0167_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1653_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1637_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1527_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0172_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1698_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1696_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1547_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1454_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1453_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1431_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1429_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1420_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1417_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1415_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1360_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1356_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1354_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1748_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1745_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1743_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1700_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1691_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1689_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1486_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1426_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1424_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1355_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1358_),
    .X(net77));
 sg13g2_tielo _3874__78 (.L_LO(net78));
 sg13g2_tielo _3875__79 (.L_LO(net79));
 sg13g2_tiehi _3857__81 (.L_HI(net81));
 sg13g2_tiehi _3858__82 (.L_HI(net82));
 sg13g2_tiehi _3859__83 (.L_HI(net83));
 sg13g2_tiehi _3860__84 (.L_HI(net84));
 sg13g2_tiehi _3861__85 (.L_HI(net85));
 sg13g2_tiehi _3864__86 (.L_HI(net86));
 sg13g2_tiehi _3865__87 (.L_HI(net87));
 sg13g2_tiehi _3866__88 (.L_HI(net88));
 sg13g2_tiehi _3867__89 (.L_HI(net89));
 sg13g2_tiehi _3868__90 (.L_HI(net90));
 sg13g2_tiehi _3869__91 (.L_HI(net91));
 sg13g2_tiehi _3870__92 (.L_HI(net92));
 sg13g2_tiehi _3871__93 (.L_HI(net93));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__94  (.L_HI(net94));
 sg13g2_tiehi \counter[10]$_SDFF_PN0__95  (.L_HI(net95));
 sg13g2_tiehi \counter[11]$_SDFF_PN0__96  (.L_HI(net96));
 sg13g2_tiehi \counter[12]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \counter[13]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \counter[14]$_SDFF_PN0__99  (.L_HI(net99));
 sg13g2_tiehi \counter[15]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \counter[16]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \counter[17]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter[18]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter[19]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \counter[20]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \counter[21]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \counter[22]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \counter[23]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \counter[24]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \counter[25]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \counter[26]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \counter[27]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \counter[28]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \counter[29]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \counter[30]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \counter[31]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \counter[9]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \depth[0]$_DFF_P__126  (.L_HI(net126));
 sg13g2_tiehi \depth[1]$_DFF_P__127  (.L_HI(net127));
 sg13g2_tiehi \depth[2]$_DFF_P__128  (.L_HI(net128));
 sg13g2_tiehi \i_project.controller_0.mode_params[2]$_DFFE_PN__129  (.L_HI(net129));
 sg13g2_tiehi \i_project.controller_0.mode_params[3]$_DFFE_PN__130  (.L_HI(net130));
 sg13g2_tiehi \i_project.controller_0.mode_params[4]$_DFFE_PN__131  (.L_HI(net131));
 sg13g2_tiehi \i_project.controller_0.mode_params[5]$_DFFE_PN__132  (.L_HI(net132));
 sg13g2_tiehi \i_project.controller_0.mode_params[6]$_DFFE_PN__133  (.L_HI(net133));
 sg13g2_tiehi \i_project.controller_0.mode_params[7]$_DFFE_PN__134  (.L_HI(net134));
 sg13g2_tiehi \i_project.controller_0.t[0]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \i_project.controller_0.t[10]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \i_project.controller_0.t[11]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \i_project.controller_0.t[1]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \i_project.controller_0.t[2]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \i_project.controller_0.t[3]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \i_project.controller_0.t[4]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \i_project.controller_0.t[5]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \i_project.controller_0.t[6]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \i_project.controller_0.t[7]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \i_project.controller_0.t[8]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \i_project.controller_0.t[9]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0__147  (.L_HI(net147));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0__148  (.L_HI(net148));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0__149  (.L_HI(net149));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0__150  (.L_HI(net150));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0__151  (.L_HI(net151));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0__152  (.L_HI(net152));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0__153  (.L_HI(net153));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0__154  (.L_HI(net154));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0__155  (.L_HI(net155));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0__156  (.L_HI(net156));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hsync$_DFFE_PP__157  (.L_HI(net157));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P__158  (.L_HI(net158));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P__159  (.L_HI(net159));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P__160  (.L_HI(net160));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P__161  (.L_HI(net161));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P__162  (.L_HI(net162));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P__163  (.L_HI(net163));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P__164  (.L_HI(net164));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P__165  (.L_HI(net165));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P__166  (.L_HI(net166));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P__167  (.L_HI(net167));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vsync$_DFFE_PP__168  (.L_HI(net168));
 sg13g2_tiehi \i_project.controller_0.voffset[0]$_DFFE_PP__169  (.L_HI(net169));
 sg13g2_tiehi \i_project.controller_0.voffset[1]$_DFFE_PP__170  (.L_HI(net170));
 sg13g2_tiehi \i_project.controller_0.voffset[2]$_DFFE_PP__171  (.L_HI(net171));
 sg13g2_tiehi \i_project.controller_0.voffset[3]$_SDFFCE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \i_project.controller_0.voffset[4]$_SDFFCE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \i_project.controller_0.voffset[5]$_DFFE_PP__174  (.L_HI(net174));
 sg13g2_tiehi \i_project.controller_0.voffset[6]$_DFFE_PP__175  (.L_HI(net175));
 sg13g2_tiehi \i_project.controller_0.voffset[7]$_SDFFCE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \lfsr[0]$_SDFF_PN1__177  (.L_HI(net177));
 sg13g2_tiehi \lfsr[10]$_SDFF_PN1__178  (.L_HI(net178));
 sg13g2_tiehi \lfsr[11]$_SDFF_PN1__179  (.L_HI(net179));
 sg13g2_tiehi \lfsr[12]$_SDFF_PN1__180  (.L_HI(net180));
 sg13g2_tiehi \lfsr[13]$_SDFF_PN1__181  (.L_HI(net181));
 sg13g2_tiehi \lfsr[14]$_SDFF_PN1__182  (.L_HI(net182));
 sg13g2_tiehi \lfsr[15]$_SDFF_PN1__183  (.L_HI(net183));
 sg13g2_tiehi \lfsr[16]$_SDFF_PN1__184  (.L_HI(net184));
 sg13g2_tiehi \lfsr[17]$_SDFF_PN1__185  (.L_HI(net185));
 sg13g2_tiehi \lfsr[18]$_SDFF_PN1__186  (.L_HI(net186));
 sg13g2_tiehi \lfsr[19]$_SDFF_PN1__187  (.L_HI(net187));
 sg13g2_tiehi \lfsr[1]$_SDFF_PN1__188  (.L_HI(net188));
 sg13g2_tiehi \lfsr[20]$_SDFF_PN1__189  (.L_HI(net189));
 sg13g2_tiehi \lfsr[21]$_SDFF_PN1__190  (.L_HI(net190));
 sg13g2_tiehi \lfsr[22]$_SDFF_PN1__191  (.L_HI(net191));
 sg13g2_tiehi \lfsr[23]$_SDFF_PN1__192  (.L_HI(net192));
 sg13g2_tiehi \lfsr[24]$_SDFF_PN1__193  (.L_HI(net193));
 sg13g2_tiehi \lfsr[25]$_SDFF_PN1__194  (.L_HI(net194));
 sg13g2_tiehi \lfsr[26]$_SDFF_PN1__195  (.L_HI(net195));
 sg13g2_tiehi \lfsr[27]$_SDFF_PN1__196  (.L_HI(net196));
 sg13g2_tiehi \lfsr[28]$_SDFF_PN1__197  (.L_HI(net197));
 sg13g2_tiehi \lfsr[29]$_SDFF_PN1__198  (.L_HI(net198));
 sg13g2_tiehi \lfsr[2]$_SDFF_PN1__199  (.L_HI(net199));
 sg13g2_tiehi \lfsr[30]$_SDFF_PN1__200  (.L_HI(net200));
 sg13g2_tiehi \lfsr[31]$_SDFF_PN1__201  (.L_HI(net201));
 sg13g2_tiehi \lfsr[3]$_SDFF_PN1__202  (.L_HI(net202));
 sg13g2_tiehi \lfsr[4]$_SDFF_PN1__203  (.L_HI(net203));
 sg13g2_tiehi \lfsr[5]$_SDFF_PN1__204  (.L_HI(net204));
 sg13g2_tiehi \lfsr[6]$_SDFF_PN1__205  (.L_HI(net205));
 sg13g2_tiehi \lfsr[7]$_SDFF_PN1__206  (.L_HI(net206));
 sg13g2_tiehi \lfsr[8]$_SDFF_PN1__207  (.L_HI(net207));
 sg13g2_tiehi \lfsr[9]$_SDFF_PN1__208  (.L_HI(net208));
 sg13g2_tiehi \project_rst_n$_DFF_P__209  (.L_HI(net209));
 sg13g2_tiehi \project_ui_in[2]$_DFF_P__210  (.L_HI(net210));
 sg13g2_tiehi \project_ui_in[3]$_DFF_P__211  (.L_HI(net211));
 sg13g2_tiehi \project_ui_in[4]$_DFF_P__212  (.L_HI(net212));
 sg13g2_tiehi \project_ui_in[5]$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \project_ui_in[6]$_DFF_P__214  (.L_HI(net214));
 sg13g2_tiehi \project_ui_in[7]$_SDFF_PN0__215  (.L_HI(net215));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_35 ();
 sg13g2_fill_1 FILLER_0_37 ();
 sg13g2_fill_2 FILLER_0_64 ();
 sg13g2_fill_1 FILLER_0_66 ();
 sg13g2_decap_4 FILLER_0_71 ();
 sg13g2_fill_1 FILLER_0_106 ();
 sg13g2_fill_2 FILLER_0_111 ();
 sg13g2_fill_2 FILLER_0_121 ();
 sg13g2_fill_2 FILLER_0_127 ();
 sg13g2_decap_4 FILLER_0_142 ();
 sg13g2_fill_2 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_4 FILLER_0_201 ();
 sg13g2_fill_2 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_fill_1 FILLER_0_240 ();
 sg13g2_decap_4 FILLER_0_271 ();
 sg13g2_decap_4 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_fill_2 FILLER_0_315 ();
 sg13g2_fill_1 FILLER_0_326 ();
 sg13g2_fill_2 FILLER_0_331 ();
 sg13g2_fill_2 FILLER_0_359 ();
 sg13g2_fill_2 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_decap_8 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_30 ();
 sg13g2_decap_4 FILLER_1_48 ();
 sg13g2_decap_4 FILLER_1_76 ();
 sg13g2_fill_1 FILLER_1_80 ();
 sg13g2_fill_2 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_94 ();
 sg13g2_decap_8 FILLER_1_101 ();
 sg13g2_decap_4 FILLER_1_108 ();
 sg13g2_fill_1 FILLER_1_117 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_fill_2 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_fill_2 FILLER_1_158 ();
 sg13g2_fill_1 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_165 ();
 sg13g2_fill_1 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_173 ();
 sg13g2_fill_2 FILLER_1_179 ();
 sg13g2_fill_2 FILLER_1_185 ();
 sg13g2_decap_4 FILLER_1_195 ();
 sg13g2_fill_2 FILLER_1_199 ();
 sg13g2_decap_4 FILLER_1_222 ();
 sg13g2_fill_1 FILLER_1_234 ();
 sg13g2_fill_1 FILLER_1_243 ();
 sg13g2_fill_1 FILLER_1_249 ();
 sg13g2_fill_1 FILLER_1_254 ();
 sg13g2_fill_2 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_260 ();
 sg13g2_fill_1 FILLER_1_266 ();
 sg13g2_fill_1 FILLER_1_272 ();
 sg13g2_fill_1 FILLER_1_277 ();
 sg13g2_fill_1 FILLER_1_304 ();
 sg13g2_fill_1 FILLER_1_348 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_4 FILLER_1_364 ();
 sg13g2_fill_1 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_51 ();
 sg13g2_fill_2 FILLER_2_58 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_decap_4 FILLER_2_73 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_decap_4 FILLER_2_94 ();
 sg13g2_fill_2 FILLER_2_98 ();
 sg13g2_fill_2 FILLER_2_129 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_fill_2 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_4 FILLER_2_154 ();
 sg13g2_fill_2 FILLER_2_158 ();
 sg13g2_fill_2 FILLER_2_165 ();
 sg13g2_fill_1 FILLER_2_167 ();
 sg13g2_fill_2 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_197 ();
 sg13g2_decap_4 FILLER_2_204 ();
 sg13g2_decap_4 FILLER_2_226 ();
 sg13g2_fill_1 FILLER_2_230 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_fill_1 FILLER_2_244 ();
 sg13g2_fill_1 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_292 ();
 sg13g2_fill_1 FILLER_2_298 ();
 sg13g2_fill_1 FILLER_2_319 ();
 sg13g2_fill_1 FILLER_2_325 ();
 sg13g2_fill_2 FILLER_2_331 ();
 sg13g2_fill_1 FILLER_2_338 ();
 sg13g2_fill_2 FILLER_2_342 ();
 sg13g2_fill_2 FILLER_2_387 ();
 sg13g2_fill_1 FILLER_2_389 ();
 sg13g2_fill_2 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_22 ();
 sg13g2_decap_4 FILLER_3_30 ();
 sg13g2_fill_2 FILLER_3_34 ();
 sg13g2_fill_2 FILLER_3_74 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_87 ();
 sg13g2_fill_1 FILLER_3_89 ();
 sg13g2_decap_4 FILLER_3_97 ();
 sg13g2_fill_1 FILLER_3_101 ();
 sg13g2_decap_4 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_167 ();
 sg13g2_fill_2 FILLER_3_178 ();
 sg13g2_decap_4 FILLER_3_186 ();
 sg13g2_fill_2 FILLER_3_190 ();
 sg13g2_decap_4 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_208 ();
 sg13g2_decap_8 FILLER_3_227 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_2 FILLER_3_246 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_279 ();
 sg13g2_fill_1 FILLER_3_284 ();
 sg13g2_fill_1 FILLER_3_311 ();
 sg13g2_fill_1 FILLER_3_338 ();
 sg13g2_fill_2 FILLER_3_398 ();
 sg13g2_fill_1 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_4 FILLER_4_26 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_fill_1 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_48 ();
 sg13g2_fill_2 FILLER_4_57 ();
 sg13g2_decap_4 FILLER_4_67 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_decap_8 FILLER_4_111 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_154 ();
 sg13g2_fill_1 FILLER_4_166 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_fill_2 FILLER_4_189 ();
 sg13g2_fill_1 FILLER_4_191 ();
 sg13g2_decap_4 FILLER_4_200 ();
 sg13g2_decap_4 FILLER_4_232 ();
 sg13g2_fill_2 FILLER_4_240 ();
 sg13g2_fill_1 FILLER_4_242 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_fill_1 FILLER_4_273 ();
 sg13g2_fill_2 FILLER_4_277 ();
 sg13g2_fill_1 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_decap_4 FILLER_4_316 ();
 sg13g2_fill_1 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_fill_1 FILLER_4_332 ();
 sg13g2_fill_1 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_347 ();
 sg13g2_fill_1 FILLER_4_352 ();
 sg13g2_fill_1 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_fill_1 FILLER_4_368 ();
 sg13g2_fill_2 FILLER_4_381 ();
 sg13g2_fill_1 FILLER_4_383 ();
 sg13g2_fill_1 FILLER_4_387 ();
 sg13g2_fill_2 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_fill_1 FILLER_5_6 ();
 sg13g2_decap_4 FILLER_5_11 ();
 sg13g2_fill_1 FILLER_5_19 ();
 sg13g2_fill_2 FILLER_5_37 ();
 sg13g2_fill_1 FILLER_5_52 ();
 sg13g2_decap_4 FILLER_5_57 ();
 sg13g2_fill_2 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_1 FILLER_5_83 ();
 sg13g2_decap_8 FILLER_5_89 ();
 sg13g2_fill_2 FILLER_5_96 ();
 sg13g2_fill_1 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_fill_1 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_144 ();
 sg13g2_fill_1 FILLER_5_149 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_1 FILLER_5_166 ();
 sg13g2_fill_2 FILLER_5_181 ();
 sg13g2_fill_2 FILLER_5_188 ();
 sg13g2_fill_1 FILLER_5_193 ();
 sg13g2_fill_2 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_decap_4 FILLER_5_233 ();
 sg13g2_decap_4 FILLER_5_251 ();
 sg13g2_fill_2 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_293 ();
 sg13g2_decap_4 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_fill_2 FILLER_5_333 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_365 ();
 sg13g2_fill_1 FILLER_5_399 ();
 sg13g2_decap_4 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_5_412 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_31 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_2 FILLER_6_44 ();
 sg13g2_fill_1 FILLER_6_46 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_decap_4 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_72 ();
 sg13g2_fill_1 FILLER_6_120 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_135 ();
 sg13g2_fill_2 FILLER_6_169 ();
 sg13g2_fill_1 FILLER_6_171 ();
 sg13g2_fill_2 FILLER_6_181 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_decap_4 FILLER_6_232 ();
 sg13g2_fill_2 FILLER_6_241 ();
 sg13g2_fill_1 FILLER_6_243 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_fill_2 FILLER_6_279 ();
 sg13g2_fill_1 FILLER_6_300 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_336 ();
 sg13g2_fill_2 FILLER_6_390 ();
 sg13g2_fill_1 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_fill_1 FILLER_7_19 ();
 sg13g2_fill_2 FILLER_7_36 ();
 sg13g2_fill_1 FILLER_7_38 ();
 sg13g2_fill_1 FILLER_7_45 ();
 sg13g2_decap_4 FILLER_7_50 ();
 sg13g2_fill_1 FILLER_7_57 ();
 sg13g2_fill_2 FILLER_7_72 ();
 sg13g2_fill_1 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_131 ();
 sg13g2_decap_8 FILLER_7_138 ();
 sg13g2_decap_4 FILLER_7_153 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_fill_1 FILLER_7_208 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_decap_4 FILLER_7_284 ();
 sg13g2_fill_2 FILLER_7_292 ();
 sg13g2_decap_4 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_fill_2 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_decap_4 FILLER_7_321 ();
 sg13g2_fill_1 FILLER_7_325 ();
 sg13g2_fill_2 FILLER_7_331 ();
 sg13g2_decap_4 FILLER_7_362 ();
 sg13g2_fill_1 FILLER_7_366 ();
 sg13g2_fill_1 FILLER_7_373 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_fill_1 FILLER_7_404 ();
 sg13g2_decap_8 FILLER_7_418 ();
 sg13g2_decap_4 FILLER_7_425 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_57 ();
 sg13g2_decap_4 FILLER_8_75 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_103 ();
 sg13g2_fill_2 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_decap_8 FILLER_8_134 ();
 sg13g2_fill_1 FILLER_8_141 ();
 sg13g2_decap_4 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_fill_2 FILLER_8_232 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_fill_1 FILLER_8_264 ();
 sg13g2_decap_4 FILLER_8_287 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_decap_4 FILLER_8_340 ();
 sg13g2_fill_2 FILLER_8_387 ();
 sg13g2_fill_2 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_40 ();
 sg13g2_fill_1 FILLER_9_45 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_fill_1 FILLER_9_80 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_fill_1 FILLER_9_116 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_200 ();
 sg13g2_fill_2 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_291 ();
 sg13g2_fill_1 FILLER_9_293 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_318 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_2 FILLER_9_343 ();
 sg13g2_fill_2 FILLER_9_348 ();
 sg13g2_fill_1 FILLER_9_350 ();
 sg13g2_fill_1 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_fill_1 FILLER_9_391 ();
 sg13g2_fill_2 FILLER_9_397 ();
 sg13g2_fill_1 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_9 ();
 sg13g2_fill_2 FILLER_10_13 ();
 sg13g2_decap_4 FILLER_10_32 ();
 sg13g2_fill_2 FILLER_10_64 ();
 sg13g2_fill_1 FILLER_10_66 ();
 sg13g2_fill_2 FILLER_10_83 ();
 sg13g2_fill_1 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_94 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_4 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_2 FILLER_10_227 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_2 FILLER_10_329 ();
 sg13g2_fill_2 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_9 ();
 sg13g2_fill_2 FILLER_11_30 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_1 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_55 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_fill_2 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_69 ();
 sg13g2_decap_4 FILLER_11_102 ();
 sg13g2_decap_4 FILLER_11_110 ();
 sg13g2_fill_2 FILLER_11_130 ();
 sg13g2_decap_4 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_171 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_fill_2 FILLER_11_193 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_220 ();
 sg13g2_fill_2 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_fill_1 FILLER_11_237 ();
 sg13g2_fill_2 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_262 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_decap_4 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_decap_4 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_4 FILLER_11_356 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_395 ();
 sg13g2_fill_1 FILLER_11_399 ();
 sg13g2_fill_1 FILLER_11_409 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_25 ();
 sg13g2_fill_2 FILLER_12_34 ();
 sg13g2_fill_1 FILLER_12_36 ();
 sg13g2_fill_2 FILLER_12_88 ();
 sg13g2_decap_4 FILLER_12_107 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_150 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_fill_2 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_fill_1 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_313 ();
 sg13g2_decap_4 FILLER_12_318 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_333 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_decap_4 FILLER_12_351 ();
 sg13g2_fill_1 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_4 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_422 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_4 ();
 sg13g2_fill_1 FILLER_13_19 ();
 sg13g2_fill_1 FILLER_13_34 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_fill_2 FILLER_13_107 ();
 sg13g2_decap_4 FILLER_13_113 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_fill_1 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_126 ();
 sg13g2_decap_4 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_fill_2 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_1 FILLER_13_162 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_178 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_fill_2 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_206 ();
 sg13g2_fill_1 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_227 ();
 sg13g2_decap_4 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_decap_4 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_363 ();
 sg13g2_decap_4 FILLER_13_373 ();
 sg13g2_fill_2 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_fill_1 FILLER_13_397 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_22 ();
 sg13g2_fill_1 FILLER_14_24 ();
 sg13g2_decap_4 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_fill_2 FILLER_14_80 ();
 sg13g2_fill_1 FILLER_14_82 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_1 FILLER_14_115 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_fill_1 FILLER_14_247 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_2 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_4 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_365 ();
 sg13g2_decap_4 FILLER_14_370 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_17 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_37 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_2 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_decap_4 FILLER_15_130 ();
 sg13g2_fill_1 FILLER_15_134 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_decap_4 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_262 ();
 sg13g2_decap_4 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_351 ();
 sg13g2_fill_2 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_fill_1 FILLER_15_397 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_fill_2 FILLER_15_418 ();
 sg13g2_decap_8 FILLER_15_423 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_44 ();
 sg13g2_decap_4 FILLER_16_55 ();
 sg13g2_fill_2 FILLER_16_99 ();
 sg13g2_fill_2 FILLER_16_104 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_152 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_197 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_2 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_1 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_4 FILLER_16_375 ();
 sg13g2_fill_2 FILLER_16_379 ();
 sg13g2_fill_1 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_9 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_1 FILLER_17_27 ();
 sg13g2_fill_2 FILLER_17_36 ();
 sg13g2_fill_2 FILLER_17_43 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_71 ();
 sg13g2_fill_1 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_86 ();
 sg13g2_decap_8 FILLER_17_92 ();
 sg13g2_decap_4 FILLER_17_99 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_160 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_decap_4 FILLER_17_395 ();
 sg13g2_fill_1 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_370 ();
 sg13g2_fill_2 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_377 ();
 sg13g2_fill_2 FILLER_18_404 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_16 ();
 sg13g2_fill_1 FILLER_19_18 ();
 sg13g2_fill_1 FILLER_19_23 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_51 ();
 sg13g2_fill_1 FILLER_19_60 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_100 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_fill_2 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_396 ();
 sg13g2_fill_1 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_fill_1 FILLER_20_89 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_decap_4 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_decap_4 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_fill_2 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_decap_4 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_decap_4 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_decap_4 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_decap_4 FILLER_21_424 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_37 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_decap_4 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_decap_4 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_fill_2 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_decap_8 FILLER_23_87 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_decap_4 FILLER_23_101 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_125 ();
 sg13g2_decap_8 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_decap_4 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_288 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_415 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_2 FILLER_24_31 ();
 sg13g2_fill_2 FILLER_24_37 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_4 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_13 ();
 sg13g2_fill_1 FILLER_25_19 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_fill_2 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_decap_4 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_fill_2 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_174 ();
 sg13g2_fill_2 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_decap_4 FILLER_25_242 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_fill_2 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_decap_4 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_30 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_287 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_fill_1 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_4 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_decap_4 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_decap_4 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_417 ();
 sg13g2_decap_4 FILLER_27_424 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_30 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_122 ();
 sg13g2_decap_4 FILLER_28_128 ();
 sg13g2_decap_4 FILLER_28_137 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_decap_4 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_decap_4 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_decap_4 FILLER_29_196 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_350 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_4 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_417 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_15 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_31_31 ();
 sg13g2_fill_1 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_38 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_2 FILLER_31_57 ();
 sg13g2_fill_2 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_78 ();
 sg13g2_fill_1 FILLER_31_89 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_decap_4 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_decap_4 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_fill_1 FILLER_31_420 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_27 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_4 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_4 FILLER_32_227 ();
 sg13g2_decap_4 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_20 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_145 ();
 sg13g2_decap_4 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_1 FILLER_33_401 ();
 sg13g2_fill_2 FILLER_33_419 ();
 sg13g2_fill_1 FILLER_33_421 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_5 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_fill_2 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_decap_4 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_35_31 ();
 sg13g2_fill_1 FILLER_35_33 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_fill_2 FILLER_35_86 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_fill_2 FILLER_35_421 ();
 sg13g2_fill_2 FILLER_35_427 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_fill_2 FILLER_36_59 ();
 sg13g2_fill_1 FILLER_36_65 ();
 sg13g2_fill_2 FILLER_36_71 ();
 sg13g2_decap_4 FILLER_36_82 ();
 sg13g2_decap_4 FILLER_36_90 ();
 sg13g2_fill_2 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_114 ();
 sg13g2_decap_8 FILLER_36_121 ();
 sg13g2_decap_4 FILLER_36_128 ();
 sg13g2_decap_4 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_160 ();
 sg13g2_decap_4 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_decap_4 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_2 FILLER_36_374 ();
 sg13g2_decap_4 FILLER_36_384 ();
 sg13g2_fill_2 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_144 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_219 ();
 sg13g2_decap_4 FILLER_37_228 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_341 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_2 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_33 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_45 ();
 sg13g2_fill_2 FILLER_38_51 ();
 sg13g2_fill_1 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_62 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_decap_4 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_decap_4 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_401 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
