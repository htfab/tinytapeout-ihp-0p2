module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_inv ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_cc ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_set_cc ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _14849_ (.A(\cpu.ex.pc[1] ),
    .X(_08141_));
 sg13g2_buf_1 _14850_ (.A(net1117),
    .X(_08142_));
 sg13g2_buf_1 _14851_ (.A(net1060),
    .X(_08143_));
 sg13g2_buf_2 _14852_ (.A(_00190_),
    .X(_08144_));
 sg13g2_buf_1 _14853_ (.A(_08144_),
    .X(_08145_));
 sg13g2_buf_1 _14854_ (.A(\cpu.ex.pc[2] ),
    .X(_08146_));
 sg13g2_buf_2 _14855_ (.A(_08146_),
    .X(_08147_));
 sg13g2_buf_1 _14856_ (.A(\cpu.ex.pc[3] ),
    .X(_08148_));
 sg13g2_inv_1 _14857_ (.Y(_08149_),
    .A(_08148_));
 sg13g2_buf_2 _14858_ (.A(_08149_),
    .X(_08150_));
 sg13g2_buf_2 _14859_ (.A(\cpu.ex.pc[4] ),
    .X(_08151_));
 sg13g2_nor2_1 _14860_ (.A(net918),
    .B(net1116),
    .Y(_08152_));
 sg13g2_nand2_1 _14861_ (.Y(_08153_),
    .A(net918),
    .B(net1116));
 sg13g2_o21ai_1 _14862_ (.B1(_08153_),
    .Y(_08154_),
    .A1(net1058),
    .A2(_08152_));
 sg13g2_and2_1 _14863_ (.A(net1059),
    .B(_08154_),
    .X(_08155_));
 sg13g2_buf_1 _14864_ (.A(_08155_),
    .X(_08156_));
 sg13g2_buf_1 _14865_ (.A(_08156_),
    .X(_08157_));
 sg13g2_buf_1 _14866_ (.A(_08157_),
    .X(_08158_));
 sg13g2_inv_2 _14867_ (.Y(_08159_),
    .A(_08146_));
 sg13g2_buf_1 _14868_ (.A(_08148_),
    .X(_08160_));
 sg13g2_nor3_1 _14869_ (.A(_08159_),
    .B(net1057),
    .C(net1116),
    .Y(_08161_));
 sg13g2_buf_2 _14870_ (.A(_08161_),
    .X(_08162_));
 sg13g2_buf_1 _14871_ (.A(_08162_),
    .X(_08163_));
 sg13g2_buf_1 _14872_ (.A(net694),
    .X(_08164_));
 sg13g2_buf_1 _14873_ (.A(net625),
    .X(_08165_));
 sg13g2_buf_1 _14874_ (.A(net560),
    .X(_08166_));
 sg13g2_nand2_1 _14875_ (.Y(_08167_),
    .A(\cpu.icache.r_data[1][16] ),
    .B(net505));
 sg13g2_nor3_1 _14876_ (.A(net1058),
    .B(net918),
    .C(_08151_),
    .Y(_08168_));
 sg13g2_buf_2 _14877_ (.A(_08168_),
    .X(_08169_));
 sg13g2_buf_1 _14878_ (.A(_08169_),
    .X(_08170_));
 sg13g2_buf_2 _14879_ (.A(net624),
    .X(_08171_));
 sg13g2_buf_1 _14880_ (.A(net559),
    .X(_08172_));
 sg13g2_buf_1 _14881_ (.A(net504),
    .X(_08173_));
 sg13g2_nor3_1 _14882_ (.A(_08159_),
    .B(net918),
    .C(net1059),
    .Y(_08174_));
 sg13g2_buf_2 _14883_ (.A(_08174_),
    .X(_08175_));
 sg13g2_buf_1 _14884_ (.A(_08175_),
    .X(_08176_));
 sg13g2_buf_1 _14885_ (.A(net623),
    .X(_08177_));
 sg13g2_buf_1 _14886_ (.A(net558),
    .X(_08178_));
 sg13g2_a22oi_1 _14887_ (.Y(_08179_),
    .B1(net503),
    .B2(\cpu.icache.r_data[7][16] ),
    .A2(net451),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_nor3_1 _14888_ (.A(_08146_),
    .B(net1057),
    .C(_08144_),
    .Y(_08180_));
 sg13g2_buf_2 _14889_ (.A(_08180_),
    .X(_08181_));
 sg13g2_buf_1 _14890_ (.A(_08181_),
    .X(_08182_));
 sg13g2_buf_1 _14891_ (.A(net693),
    .X(_08183_));
 sg13g2_nor2_1 _14892_ (.A(_08160_),
    .B(_08144_),
    .Y(_08184_));
 sg13g2_buf_2 _14893_ (.A(_08184_),
    .X(_08185_));
 sg13g2_and2_1 _14894_ (.A(net1058),
    .B(_08185_),
    .X(_08186_));
 sg13g2_buf_2 _14895_ (.A(_08186_),
    .X(_08187_));
 sg13g2_buf_1 _14896_ (.A(_08187_),
    .X(_08188_));
 sg13g2_buf_2 _14897_ (.A(_08188_),
    .X(_08189_));
 sg13g2_a22oi_1 _14898_ (.Y(_08190_),
    .B1(net502),
    .B2(\cpu.icache.r_data[5][16] ),
    .A2(net622),
    .A1(\cpu.icache.r_data[4][16] ));
 sg13g2_nor2_1 _14899_ (.A(_08146_),
    .B(_08144_),
    .Y(_08191_));
 sg13g2_and2_1 _14900_ (.A(_08160_),
    .B(_08191_),
    .X(_08192_));
 sg13g2_buf_1 _14901_ (.A(_08192_),
    .X(_08193_));
 sg13g2_buf_1 _14902_ (.A(_08193_),
    .X(_08194_));
 sg13g2_buf_1 _14903_ (.A(net692),
    .X(_08195_));
 sg13g2_nor2_2 _14904_ (.A(_08159_),
    .B(net918),
    .Y(_08196_));
 sg13g2_and2_1 _14905_ (.A(net1059),
    .B(_08196_),
    .X(_08197_));
 sg13g2_buf_2 _14906_ (.A(_08197_),
    .X(_08198_));
 sg13g2_buf_1 _14907_ (.A(_08198_),
    .X(_08199_));
 sg13g2_buf_1 _14908_ (.A(net556),
    .X(_08200_));
 sg13g2_buf_1 _14909_ (.A(net501),
    .X(_08201_));
 sg13g2_a22oi_1 _14910_ (.Y(_08202_),
    .B1(net450),
    .B2(\cpu.icache.r_data[3][16] ),
    .A2(net621),
    .A1(\cpu.icache.r_data[6][16] ));
 sg13g2_nand4_1 _14911_ (.B(_08179_),
    .C(_08190_),
    .A(_08167_),
    .Y(_08203_),
    .D(_08202_));
 sg13g2_a21o_1 _14912_ (.A2(net452),
    .A1(\cpu.icache.r_data[0][16] ),
    .B1(_08203_),
    .X(_08204_));
 sg13g2_nand2_1 _14913_ (.Y(_08205_),
    .A(net1059),
    .B(_08154_));
 sg13g2_buf_1 _14914_ (.A(_08205_),
    .X(_08206_));
 sg13g2_buf_1 _14915_ (.A(net555),
    .X(_08207_));
 sg13g2_buf_2 _14916_ (.A(net500),
    .X(_08208_));
 sg13g2_buf_1 _14917_ (.A(_08208_),
    .X(_08209_));
 sg13g2_buf_1 _14918_ (.A(net388),
    .X(_08210_));
 sg13g2_buf_1 _14919_ (.A(net500),
    .X(_08211_));
 sg13g2_buf_1 _14920_ (.A(net448),
    .X(_08212_));
 sg13g2_a22oi_1 _14921_ (.Y(_08213_),
    .B1(net450),
    .B2(\cpu.icache.r_data[3][0] ),
    .A2(net622),
    .A1(\cpu.icache.r_data[4][0] ));
 sg13g2_buf_1 _14922_ (.A(net504),
    .X(_08214_));
 sg13g2_and2_1 _14923_ (.A(\cpu.icache.r_data[6][0] ),
    .B(net692),
    .X(_08215_));
 sg13g2_a221oi_1 _14924_ (.B2(\cpu.icache.r_data[7][0] ),
    .C1(_08215_),
    .B1(net503),
    .A1(\cpu.icache.r_data[2][0] ),
    .Y(_08216_),
    .A2(net447));
 sg13g2_buf_1 _14925_ (.A(_08165_),
    .X(_08217_));
 sg13g2_a22oi_1 _14926_ (.Y(_08218_),
    .B1(net502),
    .B2(\cpu.icache.r_data[5][0] ),
    .A2(net499),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_nand4_1 _14927_ (.B(_08213_),
    .C(_08216_),
    .A(net387),
    .Y(_08219_),
    .D(_08218_));
 sg13g2_o21ai_1 _14928_ (.B1(_08219_),
    .Y(_08220_),
    .A1(\cpu.icache.r_data[0][0] ),
    .A2(net349));
 sg13g2_nor2_1 _14929_ (.A(net1060),
    .B(_08220_),
    .Y(_08221_));
 sg13g2_a21o_1 _14930_ (.A2(_08204_),
    .A1(net919),
    .B1(_08221_),
    .X(_08222_));
 sg13g2_buf_2 _14931_ (.A(_08222_),
    .X(_08223_));
 sg13g2_buf_1 _14932_ (.A(_08145_),
    .X(_08224_));
 sg13g2_buf_1 _14933_ (.A(net917),
    .X(_08225_));
 sg13g2_buf_1 _14934_ (.A(net800),
    .X(_08226_));
 sg13g2_buf_1 _14935_ (.A(net1058),
    .X(_08227_));
 sg13g2_buf_1 _14936_ (.A(net1057),
    .X(_08228_));
 sg13g2_nor2_2 _14937_ (.A(net916),
    .B(net915),
    .Y(_08229_));
 sg13g2_buf_1 _14938_ (.A(net915),
    .X(_08230_));
 sg13g2_buf_1 _14939_ (.A(_08230_),
    .X(_08231_));
 sg13g2_mux2_1 _14940_ (.A0(\cpu.icache.r_data[5][17] ),
    .A1(\cpu.icache.r_data[7][17] ),
    .S(net690),
    .X(_08232_));
 sg13g2_buf_1 _14941_ (.A(net916),
    .X(_08233_));
 sg13g2_a22oi_1 _14942_ (.Y(_08234_),
    .B1(_08232_),
    .B2(net798),
    .A2(_08229_),
    .A1(\cpu.icache.r_data[4][17] ));
 sg13g2_a22oi_1 _14943_ (.Y(_08235_),
    .B1(net450),
    .B2(\cpu.icache.r_data[3][17] ),
    .A2(net621),
    .A1(\cpu.icache.r_data[6][17] ));
 sg13g2_a22oi_1 _14944_ (.Y(_08236_),
    .B1(net505),
    .B2(\cpu.icache.r_data[1][17] ),
    .A2(net451),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_nand2_1 _14945_ (.Y(_08237_),
    .A(_08235_),
    .B(_08236_));
 sg13g2_a21oi_1 _14946_ (.A1(\cpu.icache.r_data[0][17] ),
    .A2(_08158_),
    .Y(_08238_),
    .B1(_08237_));
 sg13g2_o21ai_1 _14947_ (.B1(_08238_),
    .Y(_08239_),
    .A1(net691),
    .A2(_08234_));
 sg13g2_a22oi_1 _14948_ (.Y(_08240_),
    .B1(net450),
    .B2(\cpu.icache.r_data[3][1] ),
    .A2(net622),
    .A1(\cpu.icache.r_data[4][1] ));
 sg13g2_and2_1 _14949_ (.A(\cpu.icache.r_data[7][1] ),
    .B(net558),
    .X(_08241_));
 sg13g2_a221oi_1 _14950_ (.B2(\cpu.icache.r_data[2][1] ),
    .C1(_08241_),
    .B1(_08214_),
    .A1(\cpu.icache.r_data[6][1] ),
    .Y(_08242_),
    .A2(net621));
 sg13g2_a22oi_1 _14951_ (.Y(_08243_),
    .B1(_08189_),
    .B2(\cpu.icache.r_data[5][1] ),
    .A2(net505),
    .A1(\cpu.icache.r_data[1][1] ));
 sg13g2_nand4_1 _14952_ (.B(_08240_),
    .C(_08242_),
    .A(_08212_),
    .Y(_08244_),
    .D(_08243_));
 sg13g2_o21ai_1 _14953_ (.B1(_08244_),
    .Y(_08245_),
    .A1(\cpu.icache.r_data[0][1] ),
    .A2(net349));
 sg13g2_nor2_1 _14954_ (.A(net1060),
    .B(_08245_),
    .Y(_08246_));
 sg13g2_a21oi_1 _14955_ (.A1(net919),
    .A2(_08239_),
    .Y(_08247_),
    .B1(_08246_));
 sg13g2_buf_1 _14956_ (.A(_08247_),
    .X(_08248_));
 sg13g2_buf_1 _14957_ (.A(_08248_),
    .X(_08249_));
 sg13g2_nand2_1 _14958_ (.Y(_08250_),
    .A(_08223_),
    .B(_08249_));
 sg13g2_buf_1 _14959_ (.A(_08250_),
    .X(_08251_));
 sg13g2_inv_1 _14960_ (.Y(_08252_),
    .A(\cpu.ex.pc[1] ));
 sg13g2_buf_2 _14961_ (.A(_08252_),
    .X(_08253_));
 sg13g2_nand2_1 _14962_ (.Y(_08254_),
    .A(\cpu.icache.r_data[7][15] ),
    .B(net623));
 sg13g2_a22oi_1 _14963_ (.Y(_08255_),
    .B1(net625),
    .B2(\cpu.icache.r_data[1][15] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][15] ));
 sg13g2_a22oi_1 _14964_ (.Y(_08256_),
    .B1(net556),
    .B2(\cpu.icache.r_data[3][15] ),
    .A2(net693),
    .A1(\cpu.icache.r_data[4][15] ));
 sg13g2_a22oi_1 _14965_ (.Y(_08257_),
    .B1(_08188_),
    .B2(\cpu.icache.r_data[5][15] ),
    .A2(net692),
    .A1(\cpu.icache.r_data[6][15] ));
 sg13g2_nand4_1 _14966_ (.B(_08255_),
    .C(_08256_),
    .A(_08254_),
    .Y(_08258_),
    .D(_08257_));
 sg13g2_nand2_1 _14967_ (.Y(_08259_),
    .A(_00203_),
    .B(net506));
 sg13g2_o21ai_1 _14968_ (.B1(_08259_),
    .Y(_08260_),
    .A1(net506),
    .A2(_08258_));
 sg13g2_a22oi_1 _14969_ (.Y(_08261_),
    .B1(net623),
    .B2(\cpu.icache.r_data[7][31] ),
    .A2(net625),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_a22oi_1 _14970_ (.Y(_08262_),
    .B1(_08171_),
    .B2(\cpu.icache.r_data[2][31] ),
    .A2(_08182_),
    .A1(\cpu.icache.r_data[4][31] ));
 sg13g2_and2_1 _14971_ (.A(net1057),
    .B(net1059),
    .X(_08263_));
 sg13g2_buf_2 _14972_ (.A(_08263_),
    .X(_08264_));
 sg13g2_a22oi_1 _14973_ (.Y(_08265_),
    .B1(_08264_),
    .B2(\cpu.icache.r_data[3][31] ),
    .A2(_08185_),
    .A1(\cpu.icache.r_data[5][31] ));
 sg13g2_nand2b_1 _14974_ (.Y(_08266_),
    .B(_08227_),
    .A_N(_08265_));
 sg13g2_a21oi_1 _14975_ (.A1(\cpu.icache.r_data[6][31] ),
    .A2(net692),
    .Y(_08267_),
    .B1(net1056));
 sg13g2_and4_1 _14976_ (.A(_08261_),
    .B(_08262_),
    .C(_08266_),
    .D(_08267_),
    .X(_08268_));
 sg13g2_nand2b_1 _14977_ (.Y(_08269_),
    .B(net506),
    .A_N(_00204_));
 sg13g2_a22oi_1 _14978_ (.Y(_08270_),
    .B1(_08268_),
    .B2(_08269_),
    .A2(_08260_),
    .A1(net1056));
 sg13g2_buf_1 _14979_ (.A(_08270_),
    .X(_08271_));
 sg13g2_nor2_1 _14980_ (.A(_00202_),
    .B(net555),
    .Y(_08272_));
 sg13g2_buf_1 _14981_ (.A(_08191_),
    .X(_08273_));
 sg13g2_mux2_1 _14982_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(net1059),
    .X(_08274_));
 sg13g2_a22oi_1 _14983_ (.Y(_08275_),
    .B1(_08274_),
    .B2(_08147_),
    .A2(_08273_),
    .A1(\cpu.icache.r_data[6][30] ));
 sg13g2_nor2_1 _14984_ (.A(_08150_),
    .B(_08275_),
    .Y(_08276_));
 sg13g2_a22oi_1 _14985_ (.Y(_08277_),
    .B1(_08187_),
    .B2(\cpu.icache.r_data[5][30] ),
    .A2(_08162_),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_a22oi_1 _14986_ (.Y(_08278_),
    .B1(_08169_),
    .B2(\cpu.icache.r_data[2][30] ),
    .A2(_08181_),
    .A1(\cpu.icache.r_data[4][30] ));
 sg13g2_nand2_1 _14987_ (.Y(_08279_),
    .A(_08277_),
    .B(_08278_));
 sg13g2_nor3_1 _14988_ (.A(_08272_),
    .B(_08276_),
    .C(_08279_),
    .Y(_08280_));
 sg13g2_nand2_1 _14989_ (.Y(_08281_),
    .A(_00201_),
    .B(_08156_));
 sg13g2_a22oi_1 _14990_ (.Y(_08282_),
    .B1(_08162_),
    .B2(\cpu.icache.r_data[1][14] ),
    .A2(_08169_),
    .A1(\cpu.icache.r_data[2][14] ));
 sg13g2_a22oi_1 _14991_ (.Y(_08283_),
    .B1(_08175_),
    .B2(\cpu.icache.r_data[7][14] ),
    .A2(_08198_),
    .A1(\cpu.icache.r_data[3][14] ));
 sg13g2_nor2_1 _14992_ (.A(_08159_),
    .B(net1057),
    .Y(_08284_));
 sg13g2_buf_2 _14993_ (.A(_08284_),
    .X(_08285_));
 sg13g2_mux2_1 _14994_ (.A0(\cpu.icache.r_data[4][14] ),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(net1057),
    .X(_08286_));
 sg13g2_a22oi_1 _14995_ (.Y(_08287_),
    .B1(_08286_),
    .B2(_08159_),
    .A2(_08285_),
    .A1(\cpu.icache.r_data[5][14] ));
 sg13g2_or2_1 _14996_ (.X(_08288_),
    .B(_08287_),
    .A(net917));
 sg13g2_nand4_1 _14997_ (.B(_08282_),
    .C(_08283_),
    .A(net555),
    .Y(_08289_),
    .D(_08288_));
 sg13g2_a21oi_1 _14998_ (.A1(_08281_),
    .A2(_08289_),
    .Y(_08290_),
    .B1(net1117));
 sg13g2_a21oi_1 _14999_ (.A1(net1117),
    .A2(_08280_),
    .Y(_08291_),
    .B1(_08290_));
 sg13g2_buf_1 _15000_ (.A(_08291_),
    .X(_08292_));
 sg13g2_inv_1 _15001_ (.Y(_08293_),
    .A(_08292_));
 sg13g2_a22oi_1 _15002_ (.Y(_08294_),
    .B1(net556),
    .B2(\cpu.icache.r_data[3][13] ),
    .A2(_08181_),
    .A1(\cpu.icache.r_data[4][13] ));
 sg13g2_and2_1 _15003_ (.A(\cpu.icache.r_data[6][13] ),
    .B(_08193_),
    .X(_08295_));
 sg13g2_a221oi_1 _15004_ (.B2(\cpu.icache.r_data[7][13] ),
    .C1(_08295_),
    .B1(_08175_),
    .A1(\cpu.icache.r_data[2][13] ),
    .Y(_08296_),
    .A2(net624));
 sg13g2_a22oi_1 _15005_ (.Y(_08297_),
    .B1(_08187_),
    .B2(\cpu.icache.r_data[5][13] ),
    .A2(net694),
    .A1(\cpu.icache.r_data[1][13] ));
 sg13g2_nand4_1 _15006_ (.B(_08294_),
    .C(_08296_),
    .A(_08206_),
    .Y(_08298_),
    .D(_08297_));
 sg13g2_o21ai_1 _15007_ (.B1(_08298_),
    .Y(_08299_),
    .A1(\cpu.icache.r_data[0][13] ),
    .A2(_08207_));
 sg13g2_nand2_1 _15008_ (.Y(_08300_),
    .A(\cpu.icache.r_data[1][29] ),
    .B(_08163_));
 sg13g2_a22oi_1 _15009_ (.Y(_08301_),
    .B1(_08175_),
    .B2(\cpu.icache.r_data[7][29] ),
    .A2(net624),
    .A1(\cpu.icache.r_data[2][29] ));
 sg13g2_a22oi_1 _15010_ (.Y(_08302_),
    .B1(net557),
    .B2(\cpu.icache.r_data[5][29] ),
    .A2(_08181_),
    .A1(\cpu.icache.r_data[4][29] ));
 sg13g2_a22oi_1 _15011_ (.Y(_08303_),
    .B1(_08198_),
    .B2(\cpu.icache.r_data[3][29] ),
    .A2(_08194_),
    .A1(\cpu.icache.r_data[6][29] ));
 sg13g2_nand4_1 _15012_ (.B(_08301_),
    .C(_08302_),
    .A(_08300_),
    .Y(_08304_),
    .D(_08303_));
 sg13g2_a21oi_1 _15013_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(net506),
    .Y(_08305_),
    .B1(_08304_));
 sg13g2_mux2_1 _15014_ (.A0(_08299_),
    .A1(_08305_),
    .S(_08142_),
    .X(_08306_));
 sg13g2_buf_1 _15015_ (.A(_08306_),
    .X(_08307_));
 sg13g2_and2_1 _15016_ (.A(_08293_),
    .B(_08307_),
    .X(_08308_));
 sg13g2_buf_2 _15017_ (.A(_08308_),
    .X(_08309_));
 sg13g2_nand2_1 _15018_ (.Y(_08310_),
    .A(_08271_),
    .B(_08309_));
 sg13g2_buf_2 _15019_ (.A(_08310_),
    .X(_08311_));
 sg13g2_buf_1 _15020_ (.A(net1056),
    .X(_08312_));
 sg13g2_inv_1 _15021_ (.Y(_08313_),
    .A(_00205_));
 sg13g2_a22oi_1 _15022_ (.Y(_08314_),
    .B1(net499),
    .B2(\cpu.icache.r_data[1][10] ),
    .A2(net447),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_a22oi_1 _15023_ (.Y(_08315_),
    .B1(net558),
    .B2(\cpu.icache.r_data[7][10] ),
    .A2(net501),
    .A1(\cpu.icache.r_data[3][10] ));
 sg13g2_buf_1 _15024_ (.A(_08285_),
    .X(_08316_));
 sg13g2_buf_1 _15025_ (.A(_08228_),
    .X(_08317_));
 sg13g2_mux2_1 _15026_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(net797),
    .X(_08318_));
 sg13g2_buf_1 _15027_ (.A(_08159_),
    .X(_08319_));
 sg13g2_buf_1 _15028_ (.A(net912),
    .X(_08320_));
 sg13g2_a22oi_1 _15029_ (.Y(_08321_),
    .B1(_08318_),
    .B2(net796),
    .A2(_08316_),
    .A1(\cpu.icache.r_data[5][10] ));
 sg13g2_or2_1 _15030_ (.X(_08322_),
    .B(_08321_),
    .A(net691));
 sg13g2_nand4_1 _15031_ (.B(_08314_),
    .C(_08315_),
    .A(_08209_),
    .Y(_08323_),
    .D(_08322_));
 sg13g2_o21ai_1 _15032_ (.B1(_08323_),
    .Y(_08324_),
    .A1(_08313_),
    .A2(_08210_));
 sg13g2_nor2_1 _15033_ (.A(_00206_),
    .B(_08209_),
    .Y(_08325_));
 sg13g2_mux2_1 _15034_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(net799),
    .X(_08326_));
 sg13g2_a22oi_1 _15035_ (.Y(_08327_),
    .B1(_08326_),
    .B2(net796),
    .A2(net689),
    .A1(\cpu.icache.r_data[5][26] ));
 sg13g2_nor2_1 _15036_ (.A(net691),
    .B(_08327_),
    .Y(_08328_));
 sg13g2_a22oi_1 _15037_ (.Y(_08329_),
    .B1(net499),
    .B2(\cpu.icache.r_data[1][26] ),
    .A2(net451),
    .A1(\cpu.icache.r_data[2][26] ));
 sg13g2_a22oi_1 _15038_ (.Y(_08330_),
    .B1(net503),
    .B2(\cpu.icache.r_data[7][26] ),
    .A2(net450),
    .A1(\cpu.icache.r_data[3][26] ));
 sg13g2_nand2_1 _15039_ (.Y(_08331_),
    .A(_08329_),
    .B(_08330_));
 sg13g2_nor4_1 _15040_ (.A(net913),
    .B(_08325_),
    .C(_08328_),
    .D(_08331_),
    .Y(_08332_));
 sg13g2_a21oi_1 _15041_ (.A1(net913),
    .A2(_08324_),
    .Y(_08333_),
    .B1(_08332_));
 sg13g2_buf_1 _15042_ (.A(_08333_),
    .X(_08334_));
 sg13g2_inv_2 _15043_ (.Y(_08335_),
    .A(_08334_));
 sg13g2_nor2_1 _15044_ (.A(_00208_),
    .B(net349),
    .Y(_08336_));
 sg13g2_mux2_1 _15045_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(net690),
    .X(_08337_));
 sg13g2_a22oi_1 _15046_ (.Y(_08338_),
    .B1(_08337_),
    .B2(net796),
    .A2(net689),
    .A1(\cpu.icache.r_data[5][27] ));
 sg13g2_nor2_1 _15047_ (.A(net691),
    .B(_08338_),
    .Y(_08339_));
 sg13g2_a22oi_1 _15048_ (.Y(_08340_),
    .B1(net505),
    .B2(\cpu.icache.r_data[1][27] ),
    .A2(net451),
    .A1(\cpu.icache.r_data[2][27] ));
 sg13g2_buf_1 _15049_ (.A(_08201_),
    .X(_08341_));
 sg13g2_a22oi_1 _15050_ (.Y(_08342_),
    .B1(net503),
    .B2(\cpu.icache.r_data[7][27] ),
    .A2(net386),
    .A1(\cpu.icache.r_data[3][27] ));
 sg13g2_nand2_1 _15051_ (.Y(_08343_),
    .A(_08340_),
    .B(_08342_));
 sg13g2_nor3_1 _15052_ (.A(_08336_),
    .B(_08339_),
    .C(_08343_),
    .Y(_08344_));
 sg13g2_nand2_1 _15053_ (.Y(_08345_),
    .A(_00207_),
    .B(net452));
 sg13g2_buf_2 _15054_ (.A(net502),
    .X(_08346_));
 sg13g2_a22oi_1 _15055_ (.Y(_08347_),
    .B1(net446),
    .B2(\cpu.icache.r_data[5][11] ),
    .A2(_08166_),
    .A1(\cpu.icache.r_data[1][11] ));
 sg13g2_a22oi_1 _15056_ (.Y(_08348_),
    .B1(_08173_),
    .B2(\cpu.icache.r_data[2][11] ),
    .A2(net622),
    .A1(\cpu.icache.r_data[4][11] ));
 sg13g2_mux2_1 _15057_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(\cpu.icache.r_data[3][11] ),
    .S(_08225_),
    .X(_08349_));
 sg13g2_a22oi_1 _15058_ (.Y(_08350_),
    .B1(_08349_),
    .B2(net798),
    .A2(net914),
    .A1(\cpu.icache.r_data[6][11] ));
 sg13g2_nand2b_1 _15059_ (.Y(_08351_),
    .B(net690),
    .A_N(_08350_));
 sg13g2_nand4_1 _15060_ (.B(_08347_),
    .C(_08348_),
    .A(_08210_),
    .Y(_08352_),
    .D(_08351_));
 sg13g2_a21oi_1 _15061_ (.A1(_08345_),
    .A2(_08352_),
    .Y(_08353_),
    .B1(net1060));
 sg13g2_a21oi_1 _15062_ (.A1(net919),
    .A2(_08344_),
    .Y(_08354_),
    .B1(_08353_));
 sg13g2_buf_1 _15063_ (.A(_08354_),
    .X(_08355_));
 sg13g2_nor4_1 _15064_ (.A(net125),
    .B(_08311_),
    .C(_08335_),
    .D(net191),
    .Y(_08356_));
 sg13g2_buf_1 _15065_ (.A(\cpu.dec.r_op[5] ),
    .X(_08357_));
 sg13g2_buf_1 _15066_ (.A(_08357_),
    .X(_08358_));
 sg13g2_buf_2 _15067_ (.A(\cpu.ex.pc[12] ),
    .X(_08359_));
 sg13g2_buf_1 _15068_ (.A(_08359_),
    .X(_08360_));
 sg13g2_buf_4 _15069_ (.X(_08361_),
    .A(net1054));
 sg13g2_buf_2 _15070_ (.A(_08361_),
    .X(_08362_));
 sg13g2_buf_1 _15071_ (.A(net795),
    .X(_08363_));
 sg13g2_buf_1 _15072_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08364_));
 sg13g2_buf_1 _15073_ (.A(net1115),
    .X(_08365_));
 sg13g2_buf_1 _15074_ (.A(\cpu.dec.supmode ),
    .X(_08366_));
 sg13g2_buf_1 _15075_ (.A(net1114),
    .X(_08367_));
 sg13g2_buf_1 _15076_ (.A(net1052),
    .X(_08368_));
 sg13g2_buf_2 _15077_ (.A(_08361_),
    .X(_08369_));
 sg13g2_buf_2 _15078_ (.A(net794),
    .X(_08370_));
 sg13g2_buf_4 _15079_ (.X(_08371_),
    .A(\cpu.ex.pc[13] ));
 sg13g2_buf_1 _15080_ (.A(_08371_),
    .X(_08372_));
 sg13g2_buf_1 _15081_ (.A(net1051),
    .X(_08373_));
 sg13g2_buf_1 _15082_ (.A(net910),
    .X(_08374_));
 sg13g2_mux4_1 _15083_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net793),
    .X(_08375_));
 sg13g2_mux4_1 _15084_ (.S0(_08370_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net793),
    .X(_08376_));
 sg13g2_mux4_1 _15085_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net793),
    .X(_08377_));
 sg13g2_mux4_1 _15086_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net793),
    .X(_08378_));
 sg13g2_buf_4 _15087_ (.X(_08379_),
    .A(\cpu.ex.pc[15] ));
 sg13g2_inv_4 _15088_ (.A(_08379_),
    .Y(_08380_));
 sg13g2_buf_2 _15089_ (.A(_08380_),
    .X(_08381_));
 sg13g2_buf_2 _15090_ (.A(net909),
    .X(_08382_));
 sg13g2_buf_8 _15091_ (.A(\cpu.ex.pc[14] ),
    .X(_08383_));
 sg13g2_buf_1 _15092_ (.A(_08383_),
    .X(_08384_));
 sg13g2_buf_1 _15093_ (.A(net1050),
    .X(_08385_));
 sg13g2_buf_1 _15094_ (.A(net908),
    .X(_08386_));
 sg13g2_mux4_1 _15095_ (.S0(net792),
    .A0(_08375_),
    .A1(_08376_),
    .A2(_08377_),
    .A3(_08378_),
    .S1(net791),
    .X(_08387_));
 sg13g2_nand2_1 _15096_ (.Y(_08388_),
    .A(net911),
    .B(_08387_));
 sg13g2_mux4_1 _15097_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(_08374_),
    .X(_08389_));
 sg13g2_mux4_1 _15098_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net793),
    .X(_08390_));
 sg13g2_buf_2 _15099_ (.A(_08361_),
    .X(_08391_));
 sg13g2_buf_2 _15100_ (.A(net790),
    .X(_08392_));
 sg13g2_buf_1 _15101_ (.A(net1051),
    .X(_08393_));
 sg13g2_buf_1 _15102_ (.A(net907),
    .X(_08394_));
 sg13g2_mux4_1 _15103_ (.S0(_08392_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(_08394_),
    .X(_08395_));
 sg13g2_mux4_1 _15104_ (.S0(_08392_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(_08374_),
    .X(_08396_));
 sg13g2_mux4_1 _15105_ (.S0(net792),
    .A0(_08389_),
    .A1(_08390_),
    .A2(_08395_),
    .A3(_08396_),
    .S1(net791),
    .X(_08397_));
 sg13g2_nand2b_1 _15106_ (.Y(_08398_),
    .B(_08397_),
    .A_N(net911));
 sg13g2_nand3_1 _15107_ (.B(_08388_),
    .C(_08398_),
    .A(net1053),
    .Y(_08399_));
 sg13g2_o21ai_1 _15108_ (.B1(_08399_),
    .Y(_08400_),
    .A1(net688),
    .A2(net1053));
 sg13g2_buf_2 _15109_ (.A(_08400_),
    .X(_08401_));
 sg13g2_a22oi_1 _15110_ (.Y(_08402_),
    .B1(net621),
    .B2(\cpu.icache.r_tag[6][12] ),
    .A2(net622),
    .A1(\cpu.icache.r_tag[4][12] ));
 sg13g2_a22oi_1 _15111_ (.Y(_08403_),
    .B1(net505),
    .B2(\cpu.icache.r_tag[1][12] ),
    .A2(net451),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_mux2_1 _15112_ (.A0(\cpu.icache.r_tag[7][12] ),
    .A1(\cpu.icache.r_tag[3][12] ),
    .S(net800),
    .X(_08404_));
 sg13g2_a22oi_1 _15113_ (.Y(_08405_),
    .B1(_08185_),
    .B2(\cpu.icache.r_tag[5][12] ),
    .A2(_08404_),
    .A1(net690));
 sg13g2_nand2b_1 _15114_ (.Y(_08406_),
    .B(net798),
    .A_N(_08405_));
 sg13g2_nand4_1 _15115_ (.B(_08402_),
    .C(_08403_),
    .A(net387),
    .Y(_08407_),
    .D(_08406_));
 sg13g2_o21ai_1 _15116_ (.B1(_08407_),
    .Y(_08408_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net349));
 sg13g2_xor2_1 _15117_ (.B(_08408_),
    .A(net348),
    .X(_08409_));
 sg13g2_buf_1 _15118_ (.A(net1051),
    .X(_08410_));
 sg13g2_buf_1 _15119_ (.A(net906),
    .X(_08411_));
 sg13g2_mux4_1 _15120_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net788),
    .X(_08412_));
 sg13g2_mux4_1 _15121_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net788),
    .X(_08413_));
 sg13g2_mux4_1 _15122_ (.S0(_08370_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(net788),
    .X(_08414_));
 sg13g2_mux4_1 _15123_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net788),
    .X(_08415_));
 sg13g2_mux4_1 _15124_ (.S0(net792),
    .A0(_08412_),
    .A1(_08413_),
    .A2(_08414_),
    .A3(_08415_),
    .S1(net791),
    .X(_08416_));
 sg13g2_mux4_1 _15125_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net788),
    .X(_08417_));
 sg13g2_mux4_1 _15126_ (.S0(net688),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net788),
    .X(_08418_));
 sg13g2_mux4_1 _15127_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net793),
    .X(_08419_));
 sg13g2_mux4_1 _15128_ (.S0(net687),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(net788),
    .X(_08420_));
 sg13g2_mux4_1 _15129_ (.S0(_08382_),
    .A0(_08417_),
    .A1(_08418_),
    .A2(_08419_),
    .A3(_08420_),
    .S1(_08386_),
    .X(_08421_));
 sg13g2_mux2_1 _15130_ (.A0(_08416_),
    .A1(_08421_),
    .S(net911),
    .X(_08422_));
 sg13g2_inv_2 _15131_ (.Y(_08423_),
    .A(_08371_));
 sg13g2_nor2_1 _15132_ (.A(_08423_),
    .B(net1053),
    .Y(_08424_));
 sg13g2_a21oi_1 _15133_ (.A1(net1053),
    .A2(_08422_),
    .Y(_08425_),
    .B1(_08424_));
 sg13g2_buf_2 _15134_ (.A(_08425_),
    .X(_08426_));
 sg13g2_a22oi_1 _15135_ (.Y(_08427_),
    .B1(net450),
    .B2(\cpu.icache.r_tag[3][13] ),
    .A2(net505),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_a22oi_1 _15136_ (.Y(_08428_),
    .B1(net503),
    .B2(\cpu.icache.r_tag[7][13] ),
    .A2(net451),
    .A1(\cpu.icache.r_tag[2][13] ));
 sg13g2_mux2_1 _15137_ (.A0(\cpu.icache.r_tag[4][13] ),
    .A1(\cpu.icache.r_tag[6][13] ),
    .S(net799),
    .X(_08429_));
 sg13g2_a22oi_1 _15138_ (.Y(_08430_),
    .B1(_08429_),
    .B2(net796),
    .A2(net689),
    .A1(\cpu.icache.r_tag[5][13] ));
 sg13g2_or2_1 _15139_ (.X(_08431_),
    .B(_08430_),
    .A(_08226_));
 sg13g2_nand4_1 _15140_ (.B(_08427_),
    .C(_08428_),
    .A(net349),
    .Y(_08432_),
    .D(_08431_));
 sg13g2_o21ai_1 _15141_ (.B1(_08432_),
    .Y(_08433_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net349));
 sg13g2_xor2_1 _15142_ (.B(_08433_),
    .A(net385),
    .X(_08434_));
 sg13g2_buf_2 _15143_ (.A(_00192_),
    .X(_08435_));
 sg13g2_buf_1 _15144_ (.A(_08435_),
    .X(_08436_));
 sg13g2_buf_1 _15145_ (.A(_08371_),
    .X(_08437_));
 sg13g2_mux4_1 _15146_ (.S0(_08361_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net1048),
    .X(_08438_));
 sg13g2_mux4_1 _15147_ (.S0(_08361_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net1048),
    .X(_08439_));
 sg13g2_mux4_1 _15148_ (.S0(net1054),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1048),
    .X(_08440_));
 sg13g2_mux4_1 _15149_ (.S0(net1054),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(_08437_),
    .X(_08441_));
 sg13g2_mux4_1 _15150_ (.S0(_08380_),
    .A0(_08438_),
    .A1(_08439_),
    .A2(_08440_),
    .A3(_08441_),
    .S1(net1050),
    .X(_08442_));
 sg13g2_mux4_1 _15151_ (.S0(net1054),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net1048),
    .X(_08443_));
 sg13g2_mux4_1 _15152_ (.S0(net1054),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net1048),
    .X(_08444_));
 sg13g2_mux4_1 _15153_ (.S0(net1054),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1048),
    .X(_08445_));
 sg13g2_mux4_1 _15154_ (.S0(net1054),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net1048),
    .X(_08446_));
 sg13g2_mux4_1 _15155_ (.S0(_08380_),
    .A0(_08443_),
    .A1(_08444_),
    .A2(_08445_),
    .A3(_08446_),
    .S1(net1050),
    .X(_08447_));
 sg13g2_mux2_1 _15156_ (.A0(_08442_),
    .A1(_08447_),
    .S(net1114),
    .X(_08448_));
 sg13g2_nand2b_1 _15157_ (.Y(_08449_),
    .B(_08448_),
    .A_N(net1049));
 sg13g2_buf_2 _15158_ (.A(_08449_),
    .X(_08450_));
 sg13g2_a22oi_1 _15159_ (.Y(_08451_),
    .B1(net501),
    .B2(\cpu.icache.r_tag[3][23] ),
    .A2(net499),
    .A1(\cpu.icache.r_tag[1][23] ));
 sg13g2_a22oi_1 _15160_ (.Y(_08452_),
    .B1(net558),
    .B2(\cpu.icache.r_tag[7][23] ),
    .A2(net447),
    .A1(\cpu.icache.r_tag[2][23] ));
 sg13g2_mux2_1 _15161_ (.A0(\cpu.icache.r_tag[4][23] ),
    .A1(\cpu.icache.r_tag[6][23] ),
    .S(net797),
    .X(_08453_));
 sg13g2_a22oi_1 _15162_ (.Y(_08454_),
    .B1(_08453_),
    .B2(net912),
    .A2(net689),
    .A1(\cpu.icache.r_tag[5][23] ));
 sg13g2_or2_1 _15163_ (.X(_08455_),
    .B(_08454_),
    .A(net800));
 sg13g2_nand4_1 _15164_ (.B(_08451_),
    .C(_08452_),
    .A(net388),
    .Y(_08456_),
    .D(_08455_));
 sg13g2_o21ai_1 _15165_ (.B1(_08456_),
    .Y(_08457_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(net387));
 sg13g2_xnor2_1 _15166_ (.Y(_08458_),
    .A(net498),
    .B(_08457_));
 sg13g2_buf_1 _15167_ (.A(_08361_),
    .X(_08459_));
 sg13g2_buf_2 _15168_ (.A(net787),
    .X(_08460_));
 sg13g2_buf_1 _15169_ (.A(net1051),
    .X(_08461_));
 sg13g2_mux4_1 _15170_ (.S0(_08460_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net905),
    .X(_08462_));
 sg13g2_buf_1 _15171_ (.A(net1048),
    .X(_08463_));
 sg13g2_buf_1 _15172_ (.A(net904),
    .X(_08464_));
 sg13g2_mux4_1 _15173_ (.S0(_08460_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(_08464_),
    .X(_08465_));
 sg13g2_buf_2 _15174_ (.A(_08361_),
    .X(_08466_));
 sg13g2_mux4_1 _15175_ (.S0(_08466_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(_08461_),
    .X(_08467_));
 sg13g2_mux4_1 _15176_ (.S0(_08466_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(_08461_),
    .X(_08468_));
 sg13g2_mux4_1 _15177_ (.S0(net909),
    .A0(_08462_),
    .A1(_08465_),
    .A2(_08467_),
    .A3(_08468_),
    .S1(net908),
    .X(_08469_));
 sg13g2_mux4_1 _15178_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net905),
    .X(_08470_));
 sg13g2_mux4_1 _15179_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(net905),
    .X(_08471_));
 sg13g2_mux4_1 _15180_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(_08410_),
    .X(_08472_));
 sg13g2_mux4_1 _15181_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(_08410_),
    .X(_08473_));
 sg13g2_mux4_1 _15182_ (.S0(net909),
    .A0(_08470_),
    .A1(_08471_),
    .A2(_08472_),
    .A3(_08473_),
    .S1(_08385_),
    .X(_08474_));
 sg13g2_mux2_1 _15183_ (.A0(_08469_),
    .A1(_08474_),
    .S(net1052),
    .X(_08475_));
 sg13g2_nand2b_1 _15184_ (.Y(_08476_),
    .B(_08475_),
    .A_N(net1049));
 sg13g2_buf_1 _15185_ (.A(_08476_),
    .X(_08477_));
 sg13g2_a22oi_1 _15186_ (.Y(_08478_),
    .B1(net447),
    .B2(\cpu.icache.r_tag[2][21] ),
    .A2(net621),
    .A1(\cpu.icache.r_tag[6][21] ));
 sg13g2_a22oi_1 _15187_ (.Y(_08479_),
    .B1(net501),
    .B2(\cpu.icache.r_tag[3][21] ),
    .A2(net560),
    .A1(\cpu.icache.r_tag[1][21] ));
 sg13g2_mux2_1 _15188_ (.A0(\cpu.icache.r_tag[5][21] ),
    .A1(\cpu.icache.r_tag[7][21] ),
    .S(net797),
    .X(_08480_));
 sg13g2_a22oi_1 _15189_ (.Y(_08481_),
    .B1(_08480_),
    .B2(net916),
    .A2(_08229_),
    .A1(\cpu.icache.r_tag[4][21] ));
 sg13g2_or2_1 _15190_ (.X(_08482_),
    .B(_08481_),
    .A(net800));
 sg13g2_nand4_1 _15191_ (.B(_08478_),
    .C(_08479_),
    .A(net388),
    .Y(_08483_),
    .D(_08482_));
 sg13g2_o21ai_1 _15192_ (.B1(_08483_),
    .Y(_08484_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(net387));
 sg13g2_xnor2_1 _15193_ (.Y(_08485_),
    .A(net384),
    .B(_08484_));
 sg13g2_mux4_1 _15194_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net905),
    .X(_08486_));
 sg13g2_mux4_1 _15195_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net905),
    .X(_08487_));
 sg13g2_mux4_1 _15196_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net906),
    .X(_08488_));
 sg13g2_mux4_1 _15197_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(net906),
    .X(_08489_));
 sg13g2_mux4_1 _15198_ (.S0(net909),
    .A0(_08486_),
    .A1(_08487_),
    .A2(_08488_),
    .A3(_08489_),
    .S1(net908),
    .X(_08490_));
 sg13g2_mux4_1 _15199_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net906),
    .X(_08491_));
 sg13g2_mux4_1 _15200_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net905),
    .X(_08492_));
 sg13g2_mux4_1 _15201_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net906),
    .X(_08493_));
 sg13g2_mux4_1 _15202_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net906),
    .X(_08494_));
 sg13g2_mux4_1 _15203_ (.S0(net909),
    .A0(_08491_),
    .A1(_08492_),
    .A2(_08493_),
    .A3(_08494_),
    .S1(net908),
    .X(_08495_));
 sg13g2_mux2_1 _15204_ (.A0(_08490_),
    .A1(_08495_),
    .S(net1052),
    .X(_08496_));
 sg13g2_nand2b_1 _15205_ (.Y(_08497_),
    .B(_08496_),
    .A_N(net1049));
 sg13g2_buf_2 _15206_ (.A(_08497_),
    .X(_08498_));
 sg13g2_a22oi_1 _15207_ (.Y(_08499_),
    .B1(net558),
    .B2(\cpu.icache.r_tag[7][16] ),
    .A2(net504),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_a22oi_1 _15208_ (.Y(_08500_),
    .B1(net501),
    .B2(\cpu.icache.r_tag[3][16] ),
    .A2(net560),
    .A1(\cpu.icache.r_tag[1][16] ));
 sg13g2_mux2_1 _15209_ (.A0(\cpu.icache.r_tag[4][16] ),
    .A1(\cpu.icache.r_tag[6][16] ),
    .S(net797),
    .X(_08501_));
 sg13g2_a22oi_1 _15210_ (.Y(_08502_),
    .B1(_08501_),
    .B2(net912),
    .A2(net689),
    .A1(\cpu.icache.r_tag[5][16] ));
 sg13g2_or2_1 _15211_ (.X(_08503_),
    .B(_08502_),
    .A(net800));
 sg13g2_nand4_1 _15212_ (.B(_08499_),
    .C(_08500_),
    .A(net388),
    .Y(_08504_),
    .D(_08503_));
 sg13g2_o21ai_1 _15213_ (.B1(_08504_),
    .Y(_08505_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net387));
 sg13g2_xnor2_1 _15214_ (.Y(_08506_),
    .A(_08498_),
    .B(_08505_));
 sg13g2_mux4_1 _15215_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(net905),
    .X(_08507_));
 sg13g2_mux4_1 _15216_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net905),
    .X(_08508_));
 sg13g2_mux4_1 _15217_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net906),
    .X(_08509_));
 sg13g2_mux4_1 _15218_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net906),
    .X(_08510_));
 sg13g2_mux4_1 _15219_ (.S0(net908),
    .A0(_08507_),
    .A1(_08508_),
    .A2(_08509_),
    .A3(_08510_),
    .S1(net1052),
    .X(_08511_));
 sg13g2_a21oi_1 _15220_ (.A1(net1053),
    .A2(_08511_),
    .Y(_08512_),
    .B1(_08379_));
 sg13g2_inv_2 _15221_ (.Y(_08513_),
    .A(net1115));
 sg13g2_mux4_1 _15222_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(_08394_),
    .X(_08514_));
 sg13g2_mux4_1 _15223_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net789),
    .X(_08515_));
 sg13g2_buf_2 _15224_ (.A(net787),
    .X(_08516_));
 sg13g2_mux4_1 _15225_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net786),
    .X(_08517_));
 sg13g2_mux4_1 _15226_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net786),
    .X(_08518_));
 sg13g2_mux4_1 _15227_ (.S0(net908),
    .A0(_08514_),
    .A1(_08515_),
    .A2(_08517_),
    .A3(_08518_),
    .S1(net1052),
    .X(_08519_));
 sg13g2_nor3_1 _15228_ (.A(net792),
    .B(_08513_),
    .C(_08519_),
    .Y(_08520_));
 sg13g2_or2_1 _15229_ (.X(_08521_),
    .B(_08520_),
    .A(_08512_));
 sg13g2_buf_2 _15230_ (.A(_08521_),
    .X(_08522_));
 sg13g2_mux2_1 _15231_ (.A0(\cpu.icache.r_tag[4][15] ),
    .A1(\cpu.icache.r_tag[6][15] ),
    .S(net799),
    .X(_08523_));
 sg13g2_a22oi_1 _15232_ (.Y(_08524_),
    .B1(_08523_),
    .B2(net914),
    .A2(net501),
    .A1(\cpu.icache.r_tag[3][15] ));
 sg13g2_a22oi_1 _15233_ (.Y(_08525_),
    .B1(net502),
    .B2(\cpu.icache.r_tag[5][15] ),
    .A2(net558),
    .A1(\cpu.icache.r_tag[7][15] ));
 sg13g2_a22oi_1 _15234_ (.Y(_08526_),
    .B1(net560),
    .B2(\cpu.icache.r_tag[1][15] ),
    .A2(net504),
    .A1(\cpu.icache.r_tag[2][15] ));
 sg13g2_nand4_1 _15235_ (.B(_08524_),
    .C(_08525_),
    .A(net388),
    .Y(_08527_),
    .D(_08526_));
 sg13g2_o21ai_1 _15236_ (.B1(_08527_),
    .Y(_08528_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net387));
 sg13g2_xnor2_1 _15237_ (.Y(_08529_),
    .A(net382),
    .B(_08528_));
 sg13g2_nand4_1 _15238_ (.B(_08485_),
    .C(_08506_),
    .A(_08458_),
    .Y(_08530_),
    .D(_08529_));
 sg13g2_mux4_1 _15239_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net793),
    .X(_08531_));
 sg13g2_mux4_1 _15240_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net793),
    .X(_08532_));
 sg13g2_mux4_1 _15241_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(net789),
    .X(_08533_));
 sg13g2_mux4_1 _15242_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(net789),
    .X(_08534_));
 sg13g2_mux4_1 _15243_ (.S0(net792),
    .A0(_08531_),
    .A1(_08532_),
    .A2(_08533_),
    .A3(_08534_),
    .S1(net791),
    .X(_08535_));
 sg13g2_mux4_1 _15244_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net789),
    .X(_08536_));
 sg13g2_mux4_1 _15245_ (.S0(net686),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net789),
    .X(_08537_));
 sg13g2_mux4_1 _15246_ (.S0(_08516_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net786),
    .X(_08538_));
 sg13g2_mux4_1 _15247_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net789),
    .X(_08539_));
 sg13g2_mux4_1 _15248_ (.S0(net792),
    .A0(_08536_),
    .A1(_08537_),
    .A2(_08538_),
    .A3(_08539_),
    .S1(net791),
    .X(_08540_));
 sg13g2_mux2_1 _15249_ (.A0(_08535_),
    .A1(_08540_),
    .S(net1052),
    .X(_08541_));
 sg13g2_nand2b_1 _15250_ (.Y(_08542_),
    .B(_08541_),
    .A_N(net1049));
 sg13g2_buf_2 _15251_ (.A(_08542_),
    .X(_08543_));
 sg13g2_a22oi_1 _15252_ (.Y(_08544_),
    .B1(net558),
    .B2(\cpu.icache.r_tag[7][17] ),
    .A2(net447),
    .A1(\cpu.icache.r_tag[2][17] ));
 sg13g2_a22oi_1 _15253_ (.Y(_08545_),
    .B1(net450),
    .B2(\cpu.icache.r_tag[3][17] ),
    .A2(net499),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_mux2_1 _15254_ (.A0(\cpu.icache.r_tag[4][17] ),
    .A1(\cpu.icache.r_tag[6][17] ),
    .S(net799),
    .X(_08546_));
 sg13g2_a22oi_1 _15255_ (.Y(_08547_),
    .B1(_08546_),
    .B2(net796),
    .A2(net689),
    .A1(\cpu.icache.r_tag[5][17] ));
 sg13g2_or2_1 _15256_ (.X(_08548_),
    .B(_08547_),
    .A(net691));
 sg13g2_nand4_1 _15257_ (.B(_08544_),
    .C(_08545_),
    .A(net388),
    .Y(_08549_),
    .D(_08548_));
 sg13g2_o21ai_1 _15258_ (.B1(_08549_),
    .Y(_08550_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(net349));
 sg13g2_xnor2_1 _15259_ (.Y(_08551_),
    .A(net381),
    .B(_08550_));
 sg13g2_mux4_1 _15260_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(net789),
    .X(_08552_));
 sg13g2_mux4_1 _15261_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net789),
    .X(_08553_));
 sg13g2_mux4_1 _15262_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net786),
    .X(_08554_));
 sg13g2_mux4_1 _15263_ (.S0(_08516_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net786),
    .X(_08555_));
 sg13g2_mux4_1 _15264_ (.S0(net792),
    .A0(_08552_),
    .A1(_08553_),
    .A2(_08554_),
    .A3(_08555_),
    .S1(net791),
    .X(_08556_));
 sg13g2_mux4_1 _15265_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net786),
    .X(_08557_));
 sg13g2_mux4_1 _15266_ (.S0(net684),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net786),
    .X(_08558_));
 sg13g2_mux4_1 _15267_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(_08464_),
    .X(_08559_));
 sg13g2_mux4_1 _15268_ (.S0(net685),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net786),
    .X(_08560_));
 sg13g2_mux4_1 _15269_ (.S0(net792),
    .A0(_08557_),
    .A1(_08558_),
    .A2(_08559_),
    .A3(_08560_),
    .S1(net791),
    .X(_08561_));
 sg13g2_mux2_1 _15270_ (.A0(_08556_),
    .A1(_08561_),
    .S(net1052),
    .X(_08562_));
 sg13g2_nand2b_1 _15271_ (.Y(_08563_),
    .B(_08562_),
    .A_N(net1049));
 sg13g2_buf_2 _15272_ (.A(_08563_),
    .X(_08564_));
 sg13g2_a22oi_1 _15273_ (.Y(_08565_),
    .B1(net502),
    .B2(\cpu.icache.r_tag[5][18] ),
    .A2(net447),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_a22oi_1 _15274_ (.Y(_08566_),
    .B1(net501),
    .B2(\cpu.icache.r_tag[3][18] ),
    .A2(net499),
    .A1(\cpu.icache.r_tag[1][18] ));
 sg13g2_mux2_1 _15275_ (.A0(\cpu.icache.r_tag[4][18] ),
    .A1(\cpu.icache.r_tag[6][18] ),
    .S(net797),
    .X(_08567_));
 sg13g2_a22oi_1 _15276_ (.Y(_08568_),
    .B1(_08567_),
    .B2(net912),
    .A2(_08196_),
    .A1(\cpu.icache.r_tag[7][18] ));
 sg13g2_or2_1 _15277_ (.X(_08569_),
    .B(_08568_),
    .A(net800));
 sg13g2_nand4_1 _15278_ (.B(_08565_),
    .C(_08566_),
    .A(net388),
    .Y(_08570_),
    .D(_08569_));
 sg13g2_o21ai_1 _15279_ (.B1(_08570_),
    .Y(_08571_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net387));
 sg13g2_xnor2_1 _15280_ (.Y(_08572_),
    .A(net380),
    .B(_08571_));
 sg13g2_mux4_1 _15281_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(net907),
    .X(_08573_));
 sg13g2_mux4_1 _15282_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net907),
    .X(_08574_));
 sg13g2_mux4_1 _15283_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(_08463_),
    .X(_08575_));
 sg13g2_mux4_1 _15284_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net904),
    .X(_08576_));
 sg13g2_mux4_1 _15285_ (.S0(net909),
    .A0(_08573_),
    .A1(_08574_),
    .A2(_08575_),
    .A3(_08576_),
    .S1(net1050),
    .X(_08577_));
 sg13g2_mux4_1 _15286_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net904),
    .X(_08578_));
 sg13g2_mux4_1 _15287_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net904),
    .X(_08579_));
 sg13g2_mux4_1 _15288_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net1051),
    .X(_08580_));
 sg13g2_mux4_1 _15289_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net904),
    .X(_08581_));
 sg13g2_mux4_1 _15290_ (.S0(net909),
    .A0(_08578_),
    .A1(_08579_),
    .A2(_08580_),
    .A3(_08581_),
    .S1(net1050),
    .X(_08582_));
 sg13g2_mux2_1 _15291_ (.A0(_08577_),
    .A1(_08582_),
    .S(net1052),
    .X(_08583_));
 sg13g2_nand2b_1 _15292_ (.Y(_08584_),
    .B(_08583_),
    .A_N(net1049));
 sg13g2_buf_1 _15293_ (.A(_08584_),
    .X(_08585_));
 sg13g2_a22oi_1 _15294_ (.Y(_08586_),
    .B1(net560),
    .B2(\cpu.icache.r_tag[1][22] ),
    .A2(net504),
    .A1(\cpu.icache.r_tag[2][22] ));
 sg13g2_a22oi_1 _15295_ (.Y(_08587_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][22] ),
    .A2(net558),
    .A1(\cpu.icache.r_tag[7][22] ));
 sg13g2_mux2_1 _15296_ (.A0(\cpu.icache.r_tag[4][22] ),
    .A1(\cpu.icache.r_tag[6][22] ),
    .S(net797),
    .X(_08588_));
 sg13g2_a22oi_1 _15297_ (.Y(_08589_),
    .B1(_08588_),
    .B2(net914),
    .A2(net556),
    .A1(\cpu.icache.r_tag[3][22] ));
 sg13g2_nand4_1 _15298_ (.B(_08586_),
    .C(_08587_),
    .A(net448),
    .Y(_08590_),
    .D(_08589_));
 sg13g2_o21ai_1 _15299_ (.B1(_08590_),
    .Y(_08591_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(net448));
 sg13g2_xor2_1 _15300_ (.B(_08591_),
    .A(net445),
    .X(_08592_));
 sg13g2_mux4_1 _15301_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net907),
    .X(_08593_));
 sg13g2_mux4_1 _15302_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net910),
    .X(_08594_));
 sg13g2_mux4_1 _15303_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net907),
    .X(_08595_));
 sg13g2_mux4_1 _15304_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net907),
    .X(_08596_));
 sg13g2_mux4_1 _15305_ (.S0(_08379_),
    .A0(_08593_),
    .A1(_08594_),
    .A2(_08595_),
    .A3(_08596_),
    .S1(net1114),
    .X(_08597_));
 sg13g2_a21oi_1 _15306_ (.A1(net1053),
    .A2(_08597_),
    .Y(_08598_),
    .B1(net791));
 sg13g2_inv_1 _15307_ (.Y(_08599_),
    .A(net908));
 sg13g2_mux4_1 _15308_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(net910),
    .X(_08600_));
 sg13g2_mux4_1 _15309_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net910),
    .X(_08601_));
 sg13g2_mux4_1 _15310_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net910),
    .X(_08602_));
 sg13g2_mux4_1 _15311_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net910),
    .X(_08603_));
 sg13g2_mux4_1 _15312_ (.S0(_08379_),
    .A0(_08600_),
    .A1(_08601_),
    .A2(_08602_),
    .A3(_08603_),
    .S1(net1114),
    .X(_08604_));
 sg13g2_nor3_1 _15313_ (.A(_08599_),
    .B(_08513_),
    .C(_08604_),
    .Y(_08605_));
 sg13g2_or2_1 _15314_ (.X(_08606_),
    .B(_08605_),
    .A(_08598_));
 sg13g2_buf_2 _15315_ (.A(_08606_),
    .X(_08607_));
 sg13g2_a22oi_1 _15316_ (.Y(_08608_),
    .B1(net692),
    .B2(\cpu.icache.r_tag[6][14] ),
    .A2(net693),
    .A1(\cpu.icache.r_tag[4][14] ));
 sg13g2_a22oi_1 _15317_ (.Y(_08609_),
    .B1(net560),
    .B2(\cpu.icache.r_tag[1][14] ),
    .A2(net504),
    .A1(\cpu.icache.r_tag[2][14] ));
 sg13g2_mux2_1 _15318_ (.A0(\cpu.icache.r_tag[7][14] ),
    .A1(\cpu.icache.r_tag[3][14] ),
    .S(net917),
    .X(_08610_));
 sg13g2_a22oi_1 _15319_ (.Y(_08611_),
    .B1(_08610_),
    .B2(_08230_),
    .A2(_08185_),
    .A1(\cpu.icache.r_tag[5][14] ));
 sg13g2_nand2b_1 _15320_ (.Y(_08612_),
    .B(net798),
    .A_N(_08611_));
 sg13g2_nand4_1 _15321_ (.B(_08608_),
    .C(_08609_),
    .A(_08211_),
    .Y(_08613_),
    .D(_08612_));
 sg13g2_o21ai_1 _15322_ (.B1(_08613_),
    .Y(_08614_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(net448));
 sg13g2_xor2_1 _15323_ (.B(_08614_),
    .A(net444),
    .X(_08615_));
 sg13g2_mux4_1 _15324_ (.S0(_08362_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(_08373_),
    .X(_08616_));
 sg13g2_mux4_1 _15325_ (.S0(_08362_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(_08373_),
    .X(_08617_));
 sg13g2_mux4_1 _15326_ (.S0(_08369_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(_08393_),
    .X(_08618_));
 sg13g2_mux4_1 _15327_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net907),
    .X(_08619_));
 sg13g2_mux4_1 _15328_ (.S0(_08381_),
    .A0(_08616_),
    .A1(_08617_),
    .A2(_08618_),
    .A3(_08619_),
    .S1(net908),
    .X(_08620_));
 sg13g2_mux4_1 _15329_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(net910),
    .X(_08621_));
 sg13g2_mux4_1 _15330_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(net910),
    .X(_08622_));
 sg13g2_mux4_1 _15331_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net907),
    .X(_08623_));
 sg13g2_mux4_1 _15332_ (.S0(_08369_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(_08393_),
    .X(_08624_));
 sg13g2_mux4_1 _15333_ (.S0(net909),
    .A0(_08621_),
    .A1(_08622_),
    .A2(_08623_),
    .A3(_08624_),
    .S1(_08385_),
    .X(_08625_));
 sg13g2_mux2_1 _15334_ (.A0(_08620_),
    .A1(_08625_),
    .S(_08367_),
    .X(_08626_));
 sg13g2_nand2b_1 _15335_ (.Y(_08627_),
    .B(_08626_),
    .A_N(net1049));
 sg13g2_buf_1 _15336_ (.A(_08627_),
    .X(_08628_));
 sg13g2_a22oi_1 _15337_ (.Y(_08629_),
    .B1(net504),
    .B2(\cpu.icache.r_tag[2][20] ),
    .A2(net692),
    .A1(\cpu.icache.r_tag[6][20] ));
 sg13g2_a22oi_1 _15338_ (.Y(_08630_),
    .B1(net556),
    .B2(\cpu.icache.r_tag[3][20] ),
    .A2(net560),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_mux2_1 _15339_ (.A0(\cpu.icache.r_tag[5][20] ),
    .A1(\cpu.icache.r_tag[7][20] ),
    .S(net915),
    .X(_08631_));
 sg13g2_a22oi_1 _15340_ (.Y(_08632_),
    .B1(_08631_),
    .B2(net916),
    .A2(_08229_),
    .A1(\cpu.icache.r_tag[4][20] ));
 sg13g2_or2_1 _15341_ (.X(_08633_),
    .B(_08632_),
    .A(net800));
 sg13g2_nand4_1 _15342_ (.B(_08629_),
    .C(_08630_),
    .A(net448),
    .Y(_08634_),
    .D(_08633_));
 sg13g2_o21ai_1 _15343_ (.B1(_08634_),
    .Y(_08635_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(net388));
 sg13g2_xor2_1 _15344_ (.B(_08635_),
    .A(net443),
    .X(_08636_));
 sg13g2_nor3_1 _15345_ (.A(_08592_),
    .B(_08615_),
    .C(_08636_),
    .Y(_08637_));
 sg13g2_mux4_1 _15346_ (.S0(_08391_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(net904),
    .X(_08638_));
 sg13g2_mux4_1 _15347_ (.S0(_08391_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(_08463_),
    .X(_08639_));
 sg13g2_mux4_1 _15348_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net1051),
    .X(_08640_));
 sg13g2_mux4_1 _15349_ (.S0(_08459_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(_08372_),
    .X(_08641_));
 sg13g2_mux4_1 _15350_ (.S0(_08381_),
    .A0(_08638_),
    .A1(_08639_),
    .A2(_08640_),
    .A3(_08641_),
    .S1(net1050),
    .X(_08642_));
 sg13g2_mux4_1 _15351_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net904),
    .X(_08643_));
 sg13g2_mux4_1 _15352_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net904),
    .X(_08644_));
 sg13g2_mux4_1 _15353_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net1051),
    .X(_08645_));
 sg13g2_mux4_1 _15354_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net1051),
    .X(_08646_));
 sg13g2_mux4_1 _15355_ (.S0(_08380_),
    .A0(_08643_),
    .A1(_08644_),
    .A2(_08645_),
    .A3(_08646_),
    .S1(net1050),
    .X(_08647_));
 sg13g2_mux2_1 _15356_ (.A0(_08642_),
    .A1(_08647_),
    .S(_08367_),
    .X(_08648_));
 sg13g2_nand2b_1 _15357_ (.Y(_08649_),
    .B(_08648_),
    .A_N(net1049));
 sg13g2_buf_2 _15358_ (.A(_08649_),
    .X(_08650_));
 sg13g2_mux2_1 _15359_ (.A0(\cpu.icache.r_tag[7][19] ),
    .A1(\cpu.icache.r_tag[3][19] ),
    .S(net917),
    .X(_08651_));
 sg13g2_a22oi_1 _15360_ (.Y(_08652_),
    .B1(_08196_),
    .B2(_08651_),
    .A2(net693),
    .A1(\cpu.icache.r_tag[4][19] ));
 sg13g2_a22oi_1 _15361_ (.Y(_08653_),
    .B1(net560),
    .B2(\cpu.icache.r_tag[1][19] ),
    .A2(net504),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_a22oi_1 _15362_ (.Y(_08654_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][19] ),
    .A2(net692),
    .A1(\cpu.icache.r_tag[6][19] ));
 sg13g2_nand4_1 _15363_ (.B(_08652_),
    .C(_08653_),
    .A(net448),
    .Y(_08655_),
    .D(_08654_));
 sg13g2_o21ai_1 _15364_ (.B1(_08655_),
    .Y(_08656_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(net448));
 sg13g2_xor2_1 _15365_ (.B(_08656_),
    .A(_08650_),
    .X(_08657_));
 sg13g2_inv_1 _15366_ (.Y(_08658_),
    .A(\cpu.ex.pc[11] ));
 sg13g2_buf_1 _15367_ (.A(_08658_),
    .X(_08659_));
 sg13g2_a22oi_1 _15368_ (.Y(_08660_),
    .B1(net556),
    .B2(\cpu.icache.r_tag[3][11] ),
    .A2(net693),
    .A1(\cpu.icache.r_tag[4][11] ));
 sg13g2_a22oi_1 _15369_ (.Y(_08661_),
    .B1(net625),
    .B2(\cpu.icache.r_tag[1][11] ),
    .A2(net559),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_mux2_1 _15370_ (.A0(\cpu.icache.r_tag[5][11] ),
    .A1(\cpu.icache.r_tag[7][11] ),
    .S(net915),
    .X(_08662_));
 sg13g2_nor2_1 _15371_ (.A(net1058),
    .B(_08150_),
    .Y(_08663_));
 sg13g2_a22oi_1 _15372_ (.Y(_08664_),
    .B1(_08663_),
    .B2(\cpu.icache.r_tag[6][11] ),
    .A2(_08662_),
    .A1(net916));
 sg13g2_or2_1 _15373_ (.X(_08665_),
    .B(_08664_),
    .A(net917));
 sg13g2_nand4_1 _15374_ (.B(_08660_),
    .C(_08661_),
    .A(net500),
    .Y(_08666_),
    .D(_08665_));
 sg13g2_o21ai_1 _15375_ (.B1(_08666_),
    .Y(_08667_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net449));
 sg13g2_xnor2_1 _15376_ (.Y(_08668_),
    .A(net1047),
    .B(_08667_));
 sg13g2_buf_2 _15377_ (.A(\cpu.ex.pc[6] ),
    .X(_08669_));
 sg13g2_inv_1 _15378_ (.Y(_08670_),
    .A(_08669_));
 sg13g2_a22oi_1 _15379_ (.Y(_08671_),
    .B1(net625),
    .B2(\cpu.icache.r_tag[1][6] ),
    .A2(net692),
    .A1(\cpu.icache.r_tag[6][6] ));
 sg13g2_nand2_1 _15380_ (.Y(_08672_),
    .A(\cpu.icache.r_tag[4][6] ),
    .B(net693));
 sg13g2_a22oi_1 _15381_ (.Y(_08673_),
    .B1(_08264_),
    .B2(\cpu.icache.r_tag[3][6] ),
    .A2(_08185_),
    .A1(\cpu.icache.r_tag[5][6] ));
 sg13g2_nor2_1 _15382_ (.A(net912),
    .B(_08673_),
    .Y(_08674_));
 sg13g2_a221oi_1 _15383_ (.B2(\cpu.icache.r_tag[7][6] ),
    .C1(_08674_),
    .B1(net623),
    .A1(\cpu.icache.r_tag[2][6] ),
    .Y(_08675_),
    .A2(net559));
 sg13g2_nand4_1 _15384_ (.B(_08671_),
    .C(_08672_),
    .A(net500),
    .Y(_08676_),
    .D(_08675_));
 sg13g2_o21ai_1 _15385_ (.B1(_08676_),
    .Y(_08677_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net449));
 sg13g2_xnor2_1 _15386_ (.Y(_08678_),
    .A(net1046),
    .B(_08677_));
 sg13g2_inv_1 _15387_ (.Y(_08679_),
    .A(\cpu.ex.pc[7] ));
 sg13g2_buf_1 _15388_ (.A(_08679_),
    .X(_08680_));
 sg13g2_a22oi_1 _15389_ (.Y(_08681_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][7] ),
    .A2(net625),
    .A1(\cpu.icache.r_tag[1][7] ));
 sg13g2_a22oi_1 _15390_ (.Y(_08682_),
    .B1(net559),
    .B2(\cpu.icache.r_tag[2][7] ),
    .A2(net693),
    .A1(\cpu.icache.r_tag[4][7] ));
 sg13g2_mux2_1 _15391_ (.A0(\cpu.icache.r_tag[7][7] ),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net1059),
    .X(_08683_));
 sg13g2_a22oi_1 _15392_ (.Y(_08684_),
    .B1(_08683_),
    .B2(net916),
    .A2(net914),
    .A1(\cpu.icache.r_tag[6][7] ));
 sg13g2_nand2b_1 _15393_ (.Y(_08685_),
    .B(net799),
    .A_N(_08684_));
 sg13g2_nand4_1 _15394_ (.B(_08681_),
    .C(_08682_),
    .A(net500),
    .Y(_08686_),
    .D(_08685_));
 sg13g2_o21ai_1 _15395_ (.B1(_08686_),
    .Y(_08687_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(net449));
 sg13g2_xnor2_1 _15396_ (.Y(_08688_),
    .A(net1045),
    .B(_08687_));
 sg13g2_mux4_1 _15397_ (.S0(net798),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net690),
    .X(_08689_));
 sg13g2_mux4_1 _15398_ (.S0(net916),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(_08231_),
    .X(_08690_));
 sg13g2_mux2_1 _15399_ (.A0(_08689_),
    .A1(_08690_),
    .S(_08151_),
    .X(_08691_));
 sg13g2_nand4_1 _15400_ (.B(_08678_),
    .C(_08688_),
    .A(_08668_),
    .Y(_08692_),
    .D(_08691_));
 sg13g2_a22oi_1 _15401_ (.Y(_08693_),
    .B1(net624),
    .B2(\cpu.icache.r_tag[2][8] ),
    .A2(_08181_),
    .A1(\cpu.icache.r_tag[4][8] ));
 sg13g2_a22oi_1 _15402_ (.Y(_08694_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][8] ),
    .A2(net694),
    .A1(\cpu.icache.r_tag[1][8] ));
 sg13g2_mux2_1 _15403_ (.A0(\cpu.icache.r_tag[7][8] ),
    .A1(\cpu.icache.r_tag[3][8] ),
    .S(_08145_),
    .X(_08695_));
 sg13g2_a22oi_1 _15404_ (.Y(_08696_),
    .B1(_08695_),
    .B2(net1058),
    .A2(net914),
    .A1(\cpu.icache.r_tag[6][8] ));
 sg13g2_nand2b_1 _15405_ (.Y(_08697_),
    .B(net797),
    .A_N(_08696_));
 sg13g2_nand4_1 _15406_ (.B(_08693_),
    .C(_08694_),
    .A(net500),
    .Y(_08698_),
    .D(_08697_));
 sg13g2_o21ai_1 _15407_ (.B1(_08698_),
    .Y(_08699_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net449));
 sg13g2_xnor2_1 _15408_ (.Y(_08700_),
    .A(\cpu.ex.pc[8] ),
    .B(_08699_));
 sg13g2_buf_2 _15409_ (.A(\cpu.ex.pc[5] ),
    .X(_08701_));
 sg13g2_a22oi_1 _15410_ (.Y(_08702_),
    .B1(net623),
    .B2(\cpu.icache.r_tag[7][5] ),
    .A2(net694),
    .A1(\cpu.icache.r_tag[1][5] ));
 sg13g2_a22oi_1 _15411_ (.Y(_08703_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][5] ),
    .A2(net624),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_mux2_1 _15412_ (.A0(\cpu.icache.r_tag[4][5] ),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net915),
    .X(_08704_));
 sg13g2_a22oi_1 _15413_ (.Y(_08705_),
    .B1(_08704_),
    .B2(net914),
    .A2(net556),
    .A1(\cpu.icache.r_tag[3][5] ));
 sg13g2_nand4_1 _15414_ (.B(_08702_),
    .C(_08703_),
    .A(net500),
    .Y(_08706_),
    .D(_08705_));
 sg13g2_o21ai_1 _15415_ (.B1(_08706_),
    .Y(_08707_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net449));
 sg13g2_xnor2_1 _15416_ (.Y(_08708_),
    .A(_08701_),
    .B(_08707_));
 sg13g2_nor2_1 _15417_ (.A(_08700_),
    .B(_08708_),
    .Y(_08709_));
 sg13g2_buf_1 _15418_ (.A(\cpu.ex.pc[10] ),
    .X(_08710_));
 sg13g2_a22oi_1 _15419_ (.Y(_08711_),
    .B1(net559),
    .B2(\cpu.icache.r_tag[2][10] ),
    .A2(net693),
    .A1(\cpu.icache.r_tag[4][10] ));
 sg13g2_a22oi_1 _15420_ (.Y(_08712_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][10] ),
    .A2(net625),
    .A1(\cpu.icache.r_tag[1][10] ));
 sg13g2_mux2_1 _15421_ (.A0(\cpu.icache.r_tag[7][10] ),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net917),
    .X(_08713_));
 sg13g2_a22oi_1 _15422_ (.Y(_08714_),
    .B1(_08713_),
    .B2(net916),
    .A2(net914),
    .A1(\cpu.icache.r_tag[6][10] ));
 sg13g2_nand2b_1 _15423_ (.Y(_08715_),
    .B(net799),
    .A_N(_08714_));
 sg13g2_nand4_1 _15424_ (.B(_08711_),
    .C(_08712_),
    .A(net449),
    .Y(_08716_),
    .D(_08715_));
 sg13g2_o21ai_1 _15425_ (.B1(_08716_),
    .Y(_08717_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net449));
 sg13g2_xor2_1 _15426_ (.B(_08717_),
    .A(_08710_),
    .X(_08718_));
 sg13g2_buf_1 _15427_ (.A(\cpu.ex.pc[9] ),
    .X(_08719_));
 sg13g2_inv_1 _15428_ (.Y(_08720_),
    .A(_08719_));
 sg13g2_buf_1 _15429_ (.A(_08720_),
    .X(_08721_));
 sg13g2_mux2_1 _15430_ (.A0(\cpu.icache.r_tag[4][9] ),
    .A1(\cpu.icache.r_tag[6][9] ),
    .S(net797),
    .X(_08722_));
 sg13g2_a22oi_1 _15431_ (.Y(_08723_),
    .B1(_08722_),
    .B2(net914),
    .A2(net556),
    .A1(\cpu.icache.r_tag[3][9] ));
 sg13g2_a22oi_1 _15432_ (.Y(_08724_),
    .B1(net557),
    .B2(\cpu.icache.r_tag[5][9] ),
    .A2(net559),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_a22oi_1 _15433_ (.Y(_08725_),
    .B1(net623),
    .B2(\cpu.icache.r_tag[7][9] ),
    .A2(net625),
    .A1(\cpu.icache.r_tag[1][9] ));
 sg13g2_nand4_1 _15434_ (.B(_08723_),
    .C(_08724_),
    .A(net449),
    .Y(_08726_),
    .D(_08725_));
 sg13g2_o21ai_1 _15435_ (.B1(_08726_),
    .Y(_08727_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net448));
 sg13g2_xnor2_1 _15436_ (.Y(_08728_),
    .A(net903),
    .B(_08727_));
 sg13g2_nand3_1 _15437_ (.B(_08718_),
    .C(_08728_),
    .A(_08709_),
    .Y(_08729_));
 sg13g2_nor3_1 _15438_ (.A(_08657_),
    .B(_08692_),
    .C(_08729_),
    .Y(_08730_));
 sg13g2_nand4_1 _15439_ (.B(_08572_),
    .C(_08637_),
    .A(_08551_),
    .Y(_08731_),
    .D(_08730_));
 sg13g2_or4_2 _15440_ (.A(_08409_),
    .B(_08434_),
    .C(_08530_),
    .D(_08731_),
    .X(_08732_));
 sg13g2_inv_1 _15441_ (.Y(_08733_),
    .A(_00189_));
 sg13g2_buf_8 _15442_ (.A(\cpu.ex.ifetch ),
    .X(_08734_));
 sg13g2_buf_1 _15443_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08735_));
 sg13g2_inv_1 _15444_ (.Y(_08736_),
    .A(_08735_));
 sg13g2_buf_1 _15445_ (.A(_00193_),
    .X(_08737_));
 sg13g2_inv_1 _15446_ (.Y(_08738_),
    .A(_08737_));
 sg13g2_o21ai_1 _15447_ (.B1(_08738_),
    .Y(_08739_),
    .A1(_08734_),
    .A2(_08736_));
 sg13g2_buf_4 _15448_ (.X(_08740_),
    .A(_08739_));
 sg13g2_buf_8 _15449_ (.A(\cpu.addr[12] ),
    .X(_08741_));
 sg13g2_buf_8 _15450_ (.A(\cpu.addr[14] ),
    .X(_08742_));
 sg13g2_buf_8 _15451_ (.A(net1113),
    .X(_08743_));
 sg13g2_buf_8 _15452_ (.A(net1044),
    .X(_08744_));
 sg13g2_mux4_1 _15453_ (.S0(_08741_),
    .A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S1(net902),
    .X(_08745_));
 sg13g2_mux4_1 _15454_ (.S0(_08741_),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(net902),
    .X(_08746_));
 sg13g2_mux4_1 _15455_ (.S0(_08741_),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(net1044),
    .X(_08747_));
 sg13g2_mux4_1 _15456_ (.S0(_08741_),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net1044),
    .X(_08748_));
 sg13g2_buf_2 _15457_ (.A(\cpu.addr[15] ),
    .X(_08749_));
 sg13g2_buf_1 _15458_ (.A(\cpu.addr[13] ),
    .X(_08750_));
 sg13g2_buf_1 _15459_ (.A(_08750_),
    .X(_08751_));
 sg13g2_mux4_1 _15460_ (.S0(net1112),
    .A0(_08745_),
    .A1(_08746_),
    .A2(_08747_),
    .A3(_08748_),
    .S1(net1043),
    .X(_08752_));
 sg13g2_or2_1 _15461_ (.X(_08753_),
    .B(_08752_),
    .A(_08740_));
 sg13g2_buf_8 _15462_ (.A(_08741_),
    .X(_08754_));
 sg13g2_mux4_1 _15463_ (.S0(_08754_),
    .A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[2] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S1(net1043),
    .X(_08755_));
 sg13g2_mux4_1 _15464_ (.S0(_08754_),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(net1043),
    .X(_08756_));
 sg13g2_mux4_1 _15465_ (.S0(_08741_),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(_08750_),
    .X(_08757_));
 sg13g2_mux4_1 _15466_ (.S0(_08741_),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(net1043),
    .X(_08758_));
 sg13g2_mux4_1 _15467_ (.S0(net1112),
    .A0(_08755_),
    .A1(_08756_),
    .A2(_08757_),
    .A3(_08758_),
    .S1(net902),
    .X(_08759_));
 sg13g2_nand2b_1 _15468_ (.Y(_08760_),
    .B(_08740_),
    .A_N(_08759_));
 sg13g2_nand2_1 _15469_ (.Y(_08761_),
    .A(_08753_),
    .B(_08760_));
 sg13g2_buf_2 _15470_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08762_));
 sg13g2_nor2_1 _15471_ (.A(_08762_),
    .B(\cpu.ex.r_wmask[0] ),
    .Y(_08763_));
 sg13g2_buf_2 _15472_ (.A(_08763_),
    .X(_08764_));
 sg13g2_buf_1 _15473_ (.A(\cpu.ex.r_read_stall ),
    .X(_08765_));
 sg13g2_inv_2 _15474_ (.Y(_08766_),
    .A(net1111));
 sg13g2_buf_2 _15475_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08767_));
 sg13g2_buf_1 _15476_ (.A(\cpu.cond[0] ),
    .X(_08768_));
 sg13g2_buf_8 _15477_ (.A(_00198_),
    .X(_08769_));
 sg13g2_a21o_1 _15478_ (.A2(_08768_),
    .A1(_08767_),
    .B1(net1110),
    .X(_08770_));
 sg13g2_buf_2 _15479_ (.A(_08770_),
    .X(_08771_));
 sg13g2_nor2b_2 _15480_ (.A(_08767_),
    .B_N(_08768_),
    .Y(_08772_));
 sg13g2_nand2_1 _15481_ (.Y(_08773_),
    .A(net1115),
    .B(_00197_));
 sg13g2_a221oi_1 _15482_ (.B2(net1110),
    .C1(_08773_),
    .B1(_08772_),
    .A1(_08766_),
    .Y(_08774_),
    .A2(_08771_));
 sg13g2_o21ai_1 _15483_ (.B1(_08774_),
    .Y(_08775_),
    .A1(_08733_),
    .A2(net1111));
 sg13g2_buf_1 _15484_ (.A(\cpu.ex.io_access ),
    .X(_08776_));
 sg13g2_nor2_1 _15485_ (.A(_08513_),
    .B(_08776_),
    .Y(_08777_));
 sg13g2_nor2_1 _15486_ (.A(_08777_),
    .B(_08774_),
    .Y(_08778_));
 sg13g2_a21oi_1 _15487_ (.A1(_08764_),
    .A2(_08775_),
    .Y(_08779_),
    .B1(_08778_));
 sg13g2_nand3_1 _15488_ (.B(_08766_),
    .C(_08764_),
    .A(_00189_),
    .Y(_08780_));
 sg13g2_buf_1 _15489_ (.A(_08780_),
    .X(_08781_));
 sg13g2_buf_8 _15490_ (.A(_08383_),
    .X(_08782_));
 sg13g2_mux4_1 _15491_ (.S0(_08371_),
    .A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S1(_08782_),
    .X(_08783_));
 sg13g2_mux4_1 _15492_ (.S0(_08371_),
    .A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S1(_08782_),
    .X(_08784_));
 sg13g2_mux2_1 _15493_ (.A0(_08783_),
    .A1(_08784_),
    .S(_08360_),
    .X(_08785_));
 sg13g2_nand3b_1 _15494_ (.B(net1115),
    .C(_08734_),
    .Y(_08786_),
    .A_N(net1114));
 sg13g2_nor3_1 _15495_ (.A(_08379_),
    .B(_08785_),
    .C(_08786_),
    .Y(_08787_));
 sg13g2_mux2_1 _15496_ (.A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[12] ),
    .S(net1042),
    .X(_08788_));
 sg13g2_mux2_1 _15497_ (.A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[14] ),
    .S(net1042),
    .X(_08789_));
 sg13g2_mux2_1 _15498_ (.A0(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S(net1042),
    .X(_08790_));
 sg13g2_mux2_1 _15499_ (.A0(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S(net1042),
    .X(_08791_));
 sg13g2_mux4_1 _15500_ (.S0(_08371_),
    .A0(_08788_),
    .A1(_08789_),
    .A2(_08790_),
    .A3(_08791_),
    .S1(_08360_),
    .X(_08792_));
 sg13g2_nor3_1 _15501_ (.A(_08380_),
    .B(_08786_),
    .C(_08792_),
    .Y(_08793_));
 sg13g2_nand3_1 _15502_ (.B(net1115),
    .C(_08734_),
    .A(net1114),
    .Y(_08794_));
 sg13g2_mux4_1 _15503_ (.S0(_08359_),
    .A0(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S1(_08384_),
    .X(_08795_));
 sg13g2_mux4_1 _15504_ (.S0(_08359_),
    .A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S1(_08384_),
    .X(_08796_));
 sg13g2_mux2_1 _15505_ (.A0(_08795_),
    .A1(_08796_),
    .S(_08423_),
    .X(_08797_));
 sg13g2_nor3_1 _15506_ (.A(_08380_),
    .B(_08794_),
    .C(_08797_),
    .Y(_08798_));
 sg13g2_mux2_1 _15507_ (.A0(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S(net1042),
    .X(_08799_));
 sg13g2_mux2_1 _15508_ (.A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[20] ),
    .S(net1042),
    .X(_08800_));
 sg13g2_mux2_1 _15509_ (.A0(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S(net1042),
    .X(_08801_));
 sg13g2_mux2_1 _15510_ (.A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[21] ),
    .S(net1042),
    .X(_08802_));
 sg13g2_mux4_1 _15511_ (.S0(_08423_),
    .A0(_08799_),
    .A1(_08800_),
    .A2(_08801_),
    .A3(_08802_),
    .S1(net1054),
    .X(_08803_));
 sg13g2_nor3_1 _15512_ (.A(_08379_),
    .B(_08794_),
    .C(_08803_),
    .Y(_08804_));
 sg13g2_or4_1 _15513_ (.A(_08787_),
    .B(_08793_),
    .C(_08798_),
    .D(_08804_),
    .X(_08805_));
 sg13g2_buf_1 _15514_ (.A(_08805_),
    .X(_08806_));
 sg13g2_mux2_1 _15515_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .S(_08743_),
    .X(_08807_));
 sg13g2_mux2_1 _15516_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S(_08743_),
    .X(_08808_));
 sg13g2_mux2_1 _15517_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .S(net1113),
    .X(_08809_));
 sg13g2_mux2_1 _15518_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S(_08742_),
    .X(_08810_));
 sg13g2_mux4_1 _15519_ (.S0(_08754_),
    .A0(_08807_),
    .A1(_08808_),
    .A2(_08809_),
    .A3(_08810_),
    .S1(net1043),
    .X(_08811_));
 sg13g2_mux2_1 _15520_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .S(net1044),
    .X(_08812_));
 sg13g2_mux2_1 _15521_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S(net1044),
    .X(_08813_));
 sg13g2_mux2_1 _15522_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .S(net1044),
    .X(_08814_));
 sg13g2_mux2_1 _15523_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S(net1044),
    .X(_08815_));
 sg13g2_mux4_1 _15524_ (.S0(_08754_),
    .A0(_08812_),
    .A1(_08813_),
    .A2(_08814_),
    .A3(_08815_),
    .S1(net1043),
    .X(_08816_));
 sg13g2_mux2_1 _15525_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S(net1113),
    .X(_08817_));
 sg13g2_mux2_1 _15526_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .S(net1113),
    .X(_08818_));
 sg13g2_mux2_1 _15527_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S(net1113),
    .X(_08819_));
 sg13g2_mux2_1 _15528_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .S(_08742_),
    .X(_08820_));
 sg13g2_inv_2 _15529_ (.Y(_08821_),
    .A(_08741_));
 sg13g2_buf_4 _15530_ (.X(_08822_),
    .A(_08821_));
 sg13g2_mux4_1 _15531_ (.S0(_08822_),
    .A0(_08817_),
    .A1(_08818_),
    .A2(_08819_),
    .A3(_08820_),
    .S1(net1043),
    .X(_08823_));
 sg13g2_mux2_1 _15532_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S(net1113),
    .X(_08824_));
 sg13g2_mux2_1 _15533_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .S(net1044),
    .X(_08825_));
 sg13g2_mux2_1 _15534_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S(net1113),
    .X(_08826_));
 sg13g2_mux2_1 _15535_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .S(net1113),
    .X(_08827_));
 sg13g2_mux4_1 _15536_ (.S0(_08822_),
    .A0(_08824_),
    .A1(_08825_),
    .A2(_08826_),
    .A3(_08827_),
    .S1(net1043),
    .X(_08828_));
 sg13g2_inv_2 _15537_ (.Y(_08829_),
    .A(_08734_));
 sg13g2_buf_8 _15538_ (.A(_08829_),
    .X(_08830_));
 sg13g2_a21oi_1 _15539_ (.A1(_08830_),
    .A2(_08735_),
    .Y(_08831_),
    .B1(_08737_));
 sg13g2_buf_1 _15540_ (.A(_08831_),
    .X(_08832_));
 sg13g2_mux4_1 _15541_ (.S0(net683),
    .A0(_08811_),
    .A1(_08816_),
    .A2(_08823_),
    .A3(_08828_),
    .S1(net1112),
    .X(_08833_));
 sg13g2_nor4_1 _15542_ (.A(_08513_),
    .B(_08776_),
    .C(_08833_),
    .D(_08764_),
    .Y(_08834_));
 sg13g2_a221oi_1 _15543_ (.B2(_08806_),
    .C1(_08834_),
    .B1(_08781_),
    .A1(_08761_),
    .Y(_08835_),
    .A2(_08779_));
 sg13g2_buf_1 _15544_ (.A(_08835_),
    .X(_08836_));
 sg13g2_buf_8 _15545_ (.A(_08836_),
    .X(_08837_));
 sg13g2_buf_1 _15546_ (.A(_08837_),
    .X(_08838_));
 sg13g2_nand3b_1 _15547_ (.B(_08733_),
    .C(_08838_),
    .Y(_08839_),
    .A_N(_08732_));
 sg13g2_buf_2 _15548_ (.A(_08839_),
    .X(_08840_));
 sg13g2_buf_1 _15549_ (.A(_08840_),
    .X(_08841_));
 sg13g2_mux2_1 _15550_ (.A0(_08356_),
    .A1(_08358_),
    .S(net111),
    .X(_00016_));
 sg13g2_buf_1 _15551_ (.A(\cpu.dec.r_op[6] ),
    .X(_08842_));
 sg13g2_buf_1 _15552_ (.A(_08842_),
    .X(_08843_));
 sg13g2_buf_1 _15553_ (.A(_08843_),
    .X(_08844_));
 sg13g2_buf_1 _15554_ (.A(_08840_),
    .X(_08845_));
 sg13g2_nor2_1 _15555_ (.A(_00212_),
    .B(net500),
    .Y(_08846_));
 sg13g2_mux2_1 _15556_ (.A0(\cpu.icache.r_data[4][22] ),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(net915),
    .X(_08847_));
 sg13g2_a22oi_1 _15557_ (.Y(_08848_),
    .B1(_08847_),
    .B2(net912),
    .A2(_08285_),
    .A1(\cpu.icache.r_data[5][22] ));
 sg13g2_nor2_1 _15558_ (.A(_08225_),
    .B(_08848_),
    .Y(_08849_));
 sg13g2_a22oi_1 _15559_ (.Y(_08850_),
    .B1(net694),
    .B2(\cpu.icache.r_data[1][22] ),
    .A2(net624),
    .A1(\cpu.icache.r_data[2][22] ));
 sg13g2_a22oi_1 _15560_ (.Y(_08851_),
    .B1(_08176_),
    .B2(\cpu.icache.r_data[7][22] ),
    .A2(_08199_),
    .A1(\cpu.icache.r_data[3][22] ));
 sg13g2_nand2_1 _15561_ (.Y(_08852_),
    .A(_08850_),
    .B(_08851_));
 sg13g2_nor3_1 _15562_ (.A(_08846_),
    .B(_08849_),
    .C(_08852_),
    .Y(_08853_));
 sg13g2_nand2_1 _15563_ (.Y(_08854_),
    .A(_00211_),
    .B(net506));
 sg13g2_a22oi_1 _15564_ (.Y(_08855_),
    .B1(net694),
    .B2(\cpu.icache.r_data[1][6] ),
    .A2(net624),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_a22oi_1 _15565_ (.Y(_08856_),
    .B1(net623),
    .B2(\cpu.icache.r_data[7][6] ),
    .A2(_08198_),
    .A1(\cpu.icache.r_data[3][6] ));
 sg13g2_mux2_1 _15566_ (.A0(\cpu.icache.r_data[4][6] ),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(net1057),
    .X(_08857_));
 sg13g2_a22oi_1 _15567_ (.Y(_08858_),
    .B1(_08857_),
    .B2(_08159_),
    .A2(_08285_),
    .A1(\cpu.icache.r_data[5][6] ));
 sg13g2_or2_1 _15568_ (.X(_08859_),
    .B(_08858_),
    .A(net917));
 sg13g2_nand4_1 _15569_ (.B(_08855_),
    .C(_08856_),
    .A(_08207_),
    .Y(_08860_),
    .D(_08859_));
 sg13g2_a21oi_1 _15570_ (.A1(_08854_),
    .A2(_08860_),
    .Y(_08861_),
    .B1(net1117));
 sg13g2_a21oi_1 _15571_ (.A1(net1060),
    .A2(_08853_),
    .Y(_08862_),
    .B1(_08861_));
 sg13g2_buf_1 _15572_ (.A(_08862_),
    .X(_08863_));
 sg13g2_nor2_1 _15573_ (.A(_00210_),
    .B(net555),
    .Y(_08864_));
 sg13g2_mux2_1 _15574_ (.A0(\cpu.icache.r_data[4][21] ),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_08228_),
    .X(_08865_));
 sg13g2_a22oi_1 _15575_ (.Y(_08866_),
    .B1(_08865_),
    .B2(net912),
    .A2(_08285_),
    .A1(\cpu.icache.r_data[5][21] ));
 sg13g2_nor2_1 _15576_ (.A(net917),
    .B(_08866_),
    .Y(_08867_));
 sg13g2_a22oi_1 _15577_ (.Y(_08868_),
    .B1(net694),
    .B2(\cpu.icache.r_data[1][21] ),
    .A2(net624),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_a22oi_1 _15578_ (.Y(_08869_),
    .B1(_08175_),
    .B2(\cpu.icache.r_data[7][21] ),
    .A2(_08198_),
    .A1(\cpu.icache.r_data[3][21] ));
 sg13g2_nand2_1 _15579_ (.Y(_08870_),
    .A(_08868_),
    .B(_08869_));
 sg13g2_nor3_1 _15580_ (.A(_08864_),
    .B(_08867_),
    .C(_08870_),
    .Y(_08871_));
 sg13g2_nand2_1 _15581_ (.Y(_08872_),
    .A(_00209_),
    .B(_08157_));
 sg13g2_and2_1 _15582_ (.A(\cpu.icache.r_data[4][5] ),
    .B(_08181_),
    .X(_08873_));
 sg13g2_a221oi_1 _15583_ (.B2(\cpu.icache.r_data[7][5] ),
    .C1(_08873_),
    .B1(_08175_),
    .A1(\cpu.icache.r_data[2][5] ),
    .Y(_08874_),
    .A2(_08169_));
 sg13g2_a22oi_1 _15584_ (.Y(_08875_),
    .B1(_08187_),
    .B2(\cpu.icache.r_data[5][5] ),
    .A2(_08198_),
    .A1(\cpu.icache.r_data[3][5] ));
 sg13g2_a22oi_1 _15585_ (.Y(_08876_),
    .B1(_08163_),
    .B2(\cpu.icache.r_data[1][5] ),
    .A2(_08193_),
    .A1(\cpu.icache.r_data[6][5] ));
 sg13g2_nand4_1 _15586_ (.B(_08874_),
    .C(_08875_),
    .A(_08206_),
    .Y(_08877_),
    .D(_08876_));
 sg13g2_a21oi_1 _15587_ (.A1(_08872_),
    .A2(_08877_),
    .Y(_08878_),
    .B1(net1117));
 sg13g2_a21o_1 _15588_ (.A2(_08871_),
    .A1(net1060),
    .B1(_08878_),
    .X(_08879_));
 sg13g2_buf_2 _15589_ (.A(_08879_),
    .X(_08880_));
 sg13g2_nand2b_1 _15590_ (.Y(_08881_),
    .B(_08880_),
    .A_N(_08863_));
 sg13g2_inv_1 _15591_ (.Y(_08882_),
    .A(_08271_));
 sg13g2_nand2_1 _15592_ (.Y(_08883_),
    .A(_08293_),
    .B(_08307_));
 sg13g2_buf_2 _15593_ (.A(_08883_),
    .X(_08884_));
 sg13g2_nor2_1 _15594_ (.A(_08882_),
    .B(_08884_),
    .Y(_08885_));
 sg13g2_buf_2 _15595_ (.A(_08885_),
    .X(_08886_));
 sg13g2_inv_1 _15596_ (.Y(_08887_),
    .A(_08354_));
 sg13g2_nor2_2 _15597_ (.A(_08335_),
    .B(_08887_),
    .Y(_08888_));
 sg13g2_nand2_1 _15598_ (.Y(_08889_),
    .A(_08886_),
    .B(_08888_));
 sg13g2_nor4_1 _15599_ (.A(_08840_),
    .B(net125),
    .C(_08881_),
    .D(_08889_),
    .Y(_08890_));
 sg13g2_a21o_1 _15600_ (.A2(net110),
    .A1(net901),
    .B1(_08890_),
    .X(_00017_));
 sg13g2_buf_1 _15601_ (.A(\cpu.dec.r_op[4] ),
    .X(_08891_));
 sg13g2_buf_1 _15602_ (.A(net1109),
    .X(_08892_));
 sg13g2_buf_1 _15603_ (.A(_08840_),
    .X(_08893_));
 sg13g2_buf_1 _15604_ (.A(net622),
    .X(_08894_));
 sg13g2_nand2_1 _15605_ (.Y(_08895_),
    .A(\cpu.icache.r_data[4][12] ),
    .B(net554));
 sg13g2_a22oi_1 _15606_ (.Y(_08896_),
    .B1(net503),
    .B2(\cpu.icache.r_data[7][12] ),
    .A2(net451),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15607_ (.Y(_08897_),
    .B1(_08264_),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(_08185_),
    .A1(\cpu.icache.r_data[5][12] ));
 sg13g2_nand2b_1 _15608_ (.Y(_08898_),
    .B(_08233_),
    .A_N(_08897_));
 sg13g2_buf_1 _15609_ (.A(net621),
    .X(_08899_));
 sg13g2_a22oi_1 _15610_ (.Y(_08900_),
    .B1(net505),
    .B2(\cpu.icache.r_data[1][12] ),
    .A2(net553),
    .A1(\cpu.icache.r_data[6][12] ));
 sg13g2_nand4_1 _15611_ (.B(_08896_),
    .C(_08898_),
    .A(_08895_),
    .Y(_08901_),
    .D(_08900_));
 sg13g2_nand2_1 _15612_ (.Y(_08902_),
    .A(_00213_),
    .B(net452));
 sg13g2_o21ai_1 _15613_ (.B1(_08902_),
    .Y(_08903_),
    .A1(net452),
    .A2(_08901_));
 sg13g2_nor2_1 _15614_ (.A(_00214_),
    .B(net349),
    .Y(_08904_));
 sg13g2_mux2_1 _15615_ (.A0(\cpu.icache.r_data[4][28] ),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_08231_),
    .X(_08905_));
 sg13g2_a22oi_1 _15616_ (.Y(_08906_),
    .B1(_08905_),
    .B2(net796),
    .A2(_08316_),
    .A1(\cpu.icache.r_data[5][28] ));
 sg13g2_nor2_1 _15617_ (.A(net691),
    .B(_08906_),
    .Y(_08907_));
 sg13g2_buf_1 _15618_ (.A(net451),
    .X(_08908_));
 sg13g2_buf_1 _15619_ (.A(net505),
    .X(_08909_));
 sg13g2_a22oi_1 _15620_ (.Y(_08910_),
    .B1(net441),
    .B2(\cpu.icache.r_data[1][28] ),
    .A2(net378),
    .A1(\cpu.icache.r_data[2][28] ));
 sg13g2_buf_1 _15621_ (.A(net503),
    .X(_08911_));
 sg13g2_a22oi_1 _15622_ (.Y(_08912_),
    .B1(net440),
    .B2(\cpu.icache.r_data[7][28] ),
    .A2(net386),
    .A1(\cpu.icache.r_data[3][28] ));
 sg13g2_nand2_1 _15623_ (.Y(_08913_),
    .A(_08910_),
    .B(_08912_));
 sg13g2_nor4_1 _15624_ (.A(net913),
    .B(_08904_),
    .C(_08907_),
    .D(_08913_),
    .Y(_08914_));
 sg13g2_a21oi_1 _15625_ (.A1(net913),
    .A2(_08903_),
    .Y(_08915_),
    .B1(_08914_));
 sg13g2_buf_1 _15626_ (.A(_08915_),
    .X(_08916_));
 sg13g2_inv_2 _15627_ (.Y(_08917_),
    .A(net190));
 sg13g2_a21oi_1 _15628_ (.A1(net919),
    .A2(_08871_),
    .Y(_08918_),
    .B1(_08878_));
 sg13g2_buf_2 _15629_ (.A(_08918_),
    .X(_08919_));
 sg13g2_nor2_1 _15630_ (.A(_08863_),
    .B(_08919_),
    .Y(_08920_));
 sg13g2_a21o_1 _15631_ (.A2(_08239_),
    .A1(_08143_),
    .B1(_08246_),
    .X(_08921_));
 sg13g2_buf_2 _15632_ (.A(_08921_),
    .X(_08922_));
 sg13g2_nand2_1 _15633_ (.Y(_08923_),
    .A(_08223_),
    .B(_08922_));
 sg13g2_buf_2 _15634_ (.A(_08923_),
    .X(_08924_));
 sg13g2_nor2_1 _15635_ (.A(_08889_),
    .B(_08924_),
    .Y(_08925_));
 sg13g2_nand2_1 _15636_ (.Y(_08926_),
    .A(_08920_),
    .B(_08925_));
 sg13g2_nor3_1 _15637_ (.A(net109),
    .B(_08917_),
    .C(_08926_),
    .Y(_08927_));
 sg13g2_a21o_1 _15638_ (.A2(net110),
    .A1(_08892_),
    .B1(_08927_),
    .X(_00015_));
 sg13g2_buf_1 _15639_ (.A(_08893_),
    .X(_08928_));
 sg13g2_nand2_1 _15640_ (.Y(_08929_),
    .A(\cpu.icache.r_data[4][4] ),
    .B(_08182_));
 sg13g2_a22oi_1 _15641_ (.Y(_08930_),
    .B1(net623),
    .B2(\cpu.icache.r_data[7][4] ),
    .A2(net559),
    .A1(\cpu.icache.r_data[2][4] ));
 sg13g2_a22oi_1 _15642_ (.Y(_08931_),
    .B1(_08264_),
    .B2(\cpu.icache.r_data[3][4] ),
    .A2(_08185_),
    .A1(\cpu.icache.r_data[5][4] ));
 sg13g2_nand2b_1 _15643_ (.Y(_08932_),
    .B(_08227_),
    .A_N(_08931_));
 sg13g2_a22oi_1 _15644_ (.Y(_08933_),
    .B1(_08164_),
    .B2(\cpu.icache.r_data[1][4] ),
    .A2(_08194_),
    .A1(\cpu.icache.r_data[6][4] ));
 sg13g2_nand4_1 _15645_ (.B(_08930_),
    .C(_08932_),
    .A(_08929_),
    .Y(_08934_),
    .D(_08933_));
 sg13g2_nand2_1 _15646_ (.Y(_08935_),
    .A(_00219_),
    .B(net506));
 sg13g2_o21ai_1 _15647_ (.B1(_08935_),
    .Y(_08936_),
    .A1(net506),
    .A2(_08934_));
 sg13g2_nor2_1 _15648_ (.A(_00220_),
    .B(_08208_),
    .Y(_08937_));
 sg13g2_mux2_1 _15649_ (.A0(\cpu.icache.r_data[4][20] ),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_08317_),
    .X(_08938_));
 sg13g2_a22oi_1 _15650_ (.Y(_08939_),
    .B1(_08938_),
    .B2(net912),
    .A2(net689),
    .A1(\cpu.icache.r_data[5][20] ));
 sg13g2_nor2_1 _15651_ (.A(net800),
    .B(_08939_),
    .Y(_08940_));
 sg13g2_a22oi_1 _15652_ (.Y(_08941_),
    .B1(_08164_),
    .B2(\cpu.icache.r_data[1][20] ),
    .A2(_08171_),
    .A1(\cpu.icache.r_data[2][20] ));
 sg13g2_a22oi_1 _15653_ (.Y(_08942_),
    .B1(_08176_),
    .B2(\cpu.icache.r_data[7][20] ),
    .A2(_08199_),
    .A1(\cpu.icache.r_data[3][20] ));
 sg13g2_nand2_1 _15654_ (.Y(_08943_),
    .A(_08941_),
    .B(_08942_));
 sg13g2_nor4_1 _15655_ (.A(_08253_),
    .B(_08937_),
    .C(_08940_),
    .D(_08943_),
    .Y(_08944_));
 sg13g2_a21oi_1 _15656_ (.A1(_08253_),
    .A2(_08936_),
    .Y(_08945_),
    .B1(_08944_));
 sg13g2_buf_1 _15657_ (.A(_08945_),
    .X(_08946_));
 sg13g2_nor2_1 _15658_ (.A(_08880_),
    .B(_08946_),
    .Y(_08947_));
 sg13g2_nand3b_1 _15659_ (.B(_08915_),
    .C(_08947_),
    .Y(_08948_),
    .A_N(_08863_));
 sg13g2_buf_1 _15660_ (.A(_08948_),
    .X(_08949_));
 sg13g2_inv_1 _15661_ (.Y(_08950_),
    .A(_08949_));
 sg13g2_nand2_1 _15662_ (.Y(_08951_),
    .A(_08925_),
    .B(_08950_));
 sg13g2_nor2_1 _15663_ (.A(_00218_),
    .B(net555),
    .Y(_08952_));
 sg13g2_mux2_1 _15664_ (.A0(\cpu.icache.r_data[4][19] ),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(net1057),
    .X(_08953_));
 sg13g2_a22oi_1 _15665_ (.Y(_08954_),
    .B1(_08953_),
    .B2(_08319_),
    .A2(_08285_),
    .A1(\cpu.icache.r_data[5][19] ));
 sg13g2_nor2_1 _15666_ (.A(_08224_),
    .B(_08954_),
    .Y(_08955_));
 sg13g2_a22oi_1 _15667_ (.Y(_08956_),
    .B1(_08162_),
    .B2(\cpu.icache.r_data[1][19] ),
    .A2(_08169_),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_a22oi_1 _15668_ (.Y(_08957_),
    .B1(_08175_),
    .B2(\cpu.icache.r_data[7][19] ),
    .A2(_08198_),
    .A1(\cpu.icache.r_data[3][19] ));
 sg13g2_nand2_1 _15669_ (.Y(_08958_),
    .A(_08956_),
    .B(_08957_));
 sg13g2_nor3_1 _15670_ (.A(_08952_),
    .B(_08955_),
    .C(_08958_),
    .Y(_08959_));
 sg13g2_nand2_1 _15671_ (.Y(_08960_),
    .A(_00217_),
    .B(_08156_));
 sg13g2_a22oi_1 _15672_ (.Y(_08961_),
    .B1(_08187_),
    .B2(\cpu.icache.r_data[5][3] ),
    .A2(_08162_),
    .A1(\cpu.icache.r_data[1][3] ));
 sg13g2_a22oi_1 _15673_ (.Y(_08962_),
    .B1(_08169_),
    .B2(\cpu.icache.r_data[2][3] ),
    .A2(_08181_),
    .A1(\cpu.icache.r_data[4][3] ));
 sg13g2_mux2_1 _15674_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_08144_),
    .X(_08963_));
 sg13g2_a22oi_1 _15675_ (.Y(_08964_),
    .B1(_08963_),
    .B2(net1058),
    .A2(_08191_),
    .A1(\cpu.icache.r_data[6][3] ));
 sg13g2_nand2b_1 _15676_ (.Y(_08965_),
    .B(net915),
    .A_N(_08964_));
 sg13g2_nand4_1 _15677_ (.B(_08961_),
    .C(_08962_),
    .A(net555),
    .Y(_08966_),
    .D(_08965_));
 sg13g2_a21oi_1 _15678_ (.A1(_08960_),
    .A2(_08966_),
    .Y(_08967_),
    .B1(net1117));
 sg13g2_a21oi_1 _15679_ (.A1(_08141_),
    .A2(_08959_),
    .Y(_08968_),
    .B1(_08967_));
 sg13g2_buf_1 _15680_ (.A(_08968_),
    .X(_08969_));
 sg13g2_nor2_1 _15681_ (.A(_00216_),
    .B(net555),
    .Y(_08970_));
 sg13g2_mux2_1 _15682_ (.A0(\cpu.icache.r_data[4][18] ),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(net915),
    .X(_08971_));
 sg13g2_a22oi_1 _15683_ (.Y(_08972_),
    .B1(_08971_),
    .B2(_08319_),
    .A2(_08285_),
    .A1(\cpu.icache.r_data[5][18] ));
 sg13g2_nor2_1 _15684_ (.A(_08224_),
    .B(_08972_),
    .Y(_08973_));
 sg13g2_a22oi_1 _15685_ (.Y(_08974_),
    .B1(net694),
    .B2(\cpu.icache.r_data[1][18] ),
    .A2(_08170_),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_a22oi_1 _15686_ (.Y(_08975_),
    .B1(_08175_),
    .B2(\cpu.icache.r_data[7][18] ),
    .A2(_08198_),
    .A1(\cpu.icache.r_data[3][18] ));
 sg13g2_nand2_1 _15687_ (.Y(_08976_),
    .A(_08974_),
    .B(_08975_));
 sg13g2_nor3_1 _15688_ (.A(_08970_),
    .B(_08973_),
    .C(_08976_),
    .Y(_08977_));
 sg13g2_nand2_1 _15689_ (.Y(_08978_),
    .A(_00215_),
    .B(_08156_));
 sg13g2_a22oi_1 _15690_ (.Y(_08979_),
    .B1(_08187_),
    .B2(\cpu.icache.r_data[5][2] ),
    .A2(_08162_),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_a22oi_1 _15691_ (.Y(_08980_),
    .B1(_08170_),
    .B2(\cpu.icache.r_data[2][2] ),
    .A2(_08181_),
    .A1(\cpu.icache.r_data[4][2] ));
 sg13g2_mux2_1 _15692_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(net1059),
    .X(_08981_));
 sg13g2_a22oi_1 _15693_ (.Y(_08982_),
    .B1(_08981_),
    .B2(net1058),
    .A2(_08273_),
    .A1(\cpu.icache.r_data[6][2] ));
 sg13g2_nand2b_1 _15694_ (.Y(_08983_),
    .B(_08317_),
    .A_N(_08982_));
 sg13g2_nand4_1 _15695_ (.B(_08979_),
    .C(_08980_),
    .A(net555),
    .Y(_08984_),
    .D(_08983_));
 sg13g2_a21oi_1 _15696_ (.A1(_08978_),
    .A2(_08984_),
    .Y(_08985_),
    .B1(_08141_));
 sg13g2_a21oi_1 _15697_ (.A1(net1060),
    .A2(_08977_),
    .Y(_08986_),
    .B1(_08985_));
 sg13g2_nand2_1 _15698_ (.Y(_08987_),
    .A(_08969_),
    .B(_08986_));
 sg13g2_nor2_1 _15699_ (.A(_08951_),
    .B(_08987_),
    .Y(_08988_));
 sg13g2_nor2_1 _15700_ (.A(net125),
    .B(_08311_),
    .Y(_08989_));
 sg13g2_buf_1 _15701_ (.A(_08863_),
    .X(_08990_));
 sg13g2_buf_1 _15702_ (.A(net190),
    .X(_08991_));
 sg13g2_nor2_1 _15703_ (.A(net249),
    .B(net165),
    .Y(_08992_));
 sg13g2_nand4_1 _15704_ (.B(_08919_),
    .C(_08888_),
    .A(_08989_),
    .Y(_08993_),
    .D(_08992_));
 sg13g2_nor2b_1 _15705_ (.A(_08988_),
    .B_N(_08993_),
    .Y(_08994_));
 sg13g2_buf_1 _15706_ (.A(\cpu.dec.r_op[3] ),
    .X(_08995_));
 sg13g2_buf_1 _15707_ (.A(net1108),
    .X(_08996_));
 sg13g2_buf_1 _15708_ (.A(_08840_),
    .X(_08997_));
 sg13g2_nand2_1 _15709_ (.Y(_08998_),
    .A(_08996_),
    .B(net108));
 sg13g2_o21ai_1 _15710_ (.B1(_08998_),
    .Y(_00014_),
    .A1(net92),
    .A2(_08994_));
 sg13g2_buf_1 _15711_ (.A(\cpu.spi.r_count[7] ),
    .X(_08999_));
 sg13g2_buf_1 _15712_ (.A(\cpu.spi.r_count[3] ),
    .X(_09000_));
 sg13g2_buf_1 _15713_ (.A(\cpu.spi.r_count[0] ),
    .X(_09001_));
 sg13g2_nor2_1 _15714_ (.A(_09001_),
    .B(\cpu.spi.r_count[1] ),
    .Y(_09002_));
 sg13g2_nand2b_1 _15715_ (.Y(_09003_),
    .B(_09002_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_nor3_1 _15716_ (.A(_09000_),
    .B(\cpu.spi.r_count[4] ),
    .C(_09003_),
    .Y(_09004_));
 sg13g2_nor2b_1 _15717_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09004_),
    .Y(_09005_));
 sg13g2_nor2b_1 _15718_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09005_),
    .Y(_09006_));
 sg13g2_buf_1 _15719_ (.A(_09006_),
    .X(_09007_));
 sg13g2_nand2b_1 _15720_ (.Y(_09008_),
    .B(_09007_),
    .A_N(_08999_));
 sg13g2_buf_2 _15721_ (.A(_09008_),
    .X(_09009_));
 sg13g2_buf_2 _15722_ (.A(\cpu.addr[6] ),
    .X(_09010_));
 sg13g2_buf_1 _15723_ (.A(\cpu.addr[8] ),
    .X(_09011_));
 sg13g2_buf_1 _15724_ (.A(_09011_),
    .X(_09012_));
 sg13g2_buf_2 _15725_ (.A(\cpu.addr[7] ),
    .X(_09013_));
 sg13g2_buf_2 _15726_ (.A(_09013_),
    .X(_09014_));
 sg13g2_nor2b_1 _15727_ (.A(net1038),
    .B_N(net1037),
    .Y(_09015_));
 sg13g2_buf_1 _15728_ (.A(_09015_),
    .X(_09016_));
 sg13g2_nand2_2 _15729_ (.Y(_09017_),
    .A(_09010_),
    .B(_09016_));
 sg13g2_buf_1 _15730_ (.A(\cpu.dec.r_trap ),
    .X(_09018_));
 sg13g2_buf_1 _15731_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_09019_));
 sg13g2_or2_1 _15732_ (.X(_09020_),
    .B(net1107),
    .A(_08762_));
 sg13g2_buf_1 _15733_ (.A(_09020_),
    .X(_09021_));
 sg13g2_nand3b_1 _15734_ (.B(_09021_),
    .C(_08777_),
    .Y(_09022_),
    .A_N(_08833_));
 sg13g2_buf_1 _15735_ (.A(_09022_),
    .X(_09023_));
 sg13g2_buf_1 _15736_ (.A(_08806_),
    .X(_09024_));
 sg13g2_a221oi_1 _15737_ (.B2(_08764_),
    .C1(_08778_),
    .B1(_08775_),
    .A1(_08753_),
    .Y(_09025_),
    .A2(_08760_));
 sg13g2_a21oi_1 _15738_ (.A1(_08781_),
    .A2(_09024_),
    .Y(_09026_),
    .B1(_09025_));
 sg13g2_nand2_1 _15739_ (.Y(_09027_),
    .A(_09023_),
    .B(_09026_));
 sg13g2_buf_1 _15740_ (.A(_09027_),
    .X(_09028_));
 sg13g2_nor2_1 _15741_ (.A(_09018_),
    .B(_09028_),
    .Y(_09029_));
 sg13g2_buf_1 _15742_ (.A(\cpu.intr.r_timer ),
    .X(_09030_));
 sg13g2_buf_1 _15743_ (.A(\cpu.intr.r_swi ),
    .X(_09031_));
 sg13g2_a22oi_1 _15744_ (.Y(_09032_),
    .B1(\cpu.intr.r_enable[3] ),
    .B2(_09031_),
    .A2(\cpu.intr.r_enable[2] ),
    .A1(_09030_));
 sg13g2_buf_2 _15745_ (.A(\cpu.uart.r_x_int ),
    .X(_09033_));
 sg13g2_buf_1 _15746_ (.A(\cpu.uart.r_r_int ),
    .X(_09034_));
 sg13g2_o21ai_1 _15747_ (.B1(\cpu.intr.r_enable[0] ),
    .Y(_09035_),
    .A1(_09033_),
    .A2(_09034_));
 sg13g2_buf_1 _15748_ (.A(\cpu.intr.r_clock ),
    .X(_09036_));
 sg13g2_buf_1 _15749_ (.A(\cpu.intr.r_enable[1] ),
    .X(_09037_));
 sg13g2_buf_2 _15750_ (.A(\cpu.intr.spi_intr ),
    .X(_09038_));
 sg13g2_a22oi_1 _15751_ (.Y(_09039_),
    .B1(_09038_),
    .B2(\cpu.intr.r_enable[5] ),
    .A2(_09037_),
    .A1(_09036_));
 sg13g2_nand3_1 _15752_ (.B(_09035_),
    .C(_09039_),
    .A(_09032_),
    .Y(_09040_));
 sg13g2_inv_1 _15753_ (.Y(_09041_),
    .A(_09040_));
 sg13g2_buf_1 _15754_ (.A(\cpu.gpio.r_enable_in[1] ),
    .X(_09042_));
 sg13g2_buf_2 _15755_ (.A(ui_in[1]),
    .X(_09043_));
 sg13g2_buf_1 _15756_ (.A(\cpu.gpio.r_enable_in[2] ),
    .X(_09044_));
 sg13g2_buf_2 _15757_ (.A(ui_in[2]),
    .X(_09045_));
 sg13g2_a22oi_1 _15758_ (.Y(_09046_),
    .B1(_09044_),
    .B2(_09045_),
    .A2(_09043_),
    .A1(_09042_));
 sg13g2_buf_2 _15759_ (.A(uio_in[6]),
    .X(_09047_));
 sg13g2_buf_1 _15760_ (.A(uio_in[7]),
    .X(_09048_));
 sg13g2_a22oi_1 _15761_ (.Y(_09049_),
    .B1(\cpu.gpio.r_enable_io[7] ),
    .B2(_09048_),
    .A2(_09047_),
    .A1(\cpu.gpio.r_enable_io[6] ));
 sg13g2_buf_1 _15762_ (.A(\cpu.gpio.r_enable_in[0] ),
    .X(_09050_));
 sg13g2_buf_2 _15763_ (.A(ui_in[0]),
    .X(_09051_));
 sg13g2_buf_1 _15764_ (.A(uio_in[4]),
    .X(_09052_));
 sg13g2_a22oi_1 _15765_ (.Y(_09053_),
    .B1(\cpu.gpio.r_enable_io[4] ),
    .B2(_09052_),
    .A2(_09051_),
    .A1(_09050_));
 sg13g2_buf_1 _15766_ (.A(\cpu.gpio.r_enable_in[3] ),
    .X(_09054_));
 sg13g2_buf_2 _15767_ (.A(ui_in[3]),
    .X(_09055_));
 sg13g2_buf_1 _15768_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_09056_));
 sg13g2_buf_2 _15769_ (.A(uio_in[5]),
    .X(_09057_));
 sg13g2_a22oi_1 _15770_ (.Y(_09058_),
    .B1(_09056_),
    .B2(_09057_),
    .A2(_09055_),
    .A1(_09054_));
 sg13g2_nand4_1 _15771_ (.B(_09049_),
    .C(_09053_),
    .A(_09046_),
    .Y(_09059_),
    .D(_09058_));
 sg13g2_buf_1 _15772_ (.A(_09059_),
    .X(_09060_));
 sg13g2_buf_2 _15773_ (.A(ui_in[5]),
    .X(_09061_));
 sg13g2_nand2_1 _15774_ (.Y(_09062_),
    .A(\cpu.gpio.r_enable_in[5] ),
    .B(_09061_));
 sg13g2_buf_2 _15775_ (.A(ui_in[7]),
    .X(_09063_));
 sg13g2_nand2_1 _15776_ (.Y(_09064_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_09063_));
 sg13g2_buf_2 _15777_ (.A(ui_in[4]),
    .X(_09065_));
 sg13g2_nand2_1 _15778_ (.Y(_09066_),
    .A(\cpu.gpio.r_enable_in[4] ),
    .B(_09065_));
 sg13g2_buf_2 _15779_ (.A(ui_in[6]),
    .X(_09067_));
 sg13g2_nand2_1 _15780_ (.Y(_09068_),
    .A(\cpu.gpio.r_enable_in[6] ),
    .B(_09067_));
 sg13g2_nand4_1 _15781_ (.B(_09064_),
    .C(_09066_),
    .A(_09062_),
    .Y(_09069_),
    .D(_09068_));
 sg13g2_buf_1 _15782_ (.A(_09069_),
    .X(_09070_));
 sg13g2_buf_1 _15783_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09071_));
 sg13g2_o21ai_1 _15784_ (.B1(_09071_),
    .Y(_09072_),
    .A1(_09060_),
    .A2(_09070_));
 sg13g2_buf_2 _15785_ (.A(\cpu.ex.r_ie ),
    .X(_09073_));
 sg13g2_inv_1 _15786_ (.Y(_09074_),
    .A(_09073_));
 sg13g2_a21oi_2 _15787_ (.B1(_09074_),
    .Y(_09075_),
    .A2(_09072_),
    .A1(_09041_));
 sg13g2_nand2_1 _15788_ (.Y(_09076_),
    .A(net1114),
    .B(_09075_));
 sg13g2_and2_1 _15789_ (.A(_09029_),
    .B(_09076_),
    .X(_09077_));
 sg13g2_buf_1 _15790_ (.A(_09077_),
    .X(_09078_));
 sg13g2_buf_1 _15791_ (.A(\cpu.addr[1] ),
    .X(_09079_));
 sg13g2_buf_1 _15792_ (.A(net1106),
    .X(_09080_));
 sg13g2_buf_2 _15793_ (.A(\cpu.addr[2] ),
    .X(_09081_));
 sg13g2_buf_1 _15794_ (.A(_09081_),
    .X(_09082_));
 sg13g2_buf_2 _15795_ (.A(_09082_),
    .X(_09083_));
 sg13g2_buf_2 _15796_ (.A(net900),
    .X(_09084_));
 sg13g2_buf_1 _15797_ (.A(net784),
    .X(_09085_));
 sg13g2_buf_1 _15798_ (.A(net682),
    .X(_09086_));
 sg13g2_buf_1 _15799_ (.A(\cpu.addr[3] ),
    .X(_09087_));
 sg13g2_buf_8 _15800_ (.A(_09087_),
    .X(_09088_));
 sg13g2_buf_1 _15801_ (.A(net1034),
    .X(_09089_));
 sg13g2_buf_2 _15802_ (.A(_09089_),
    .X(_09090_));
 sg13g2_buf_1 _15803_ (.A(net783),
    .X(_09091_));
 sg13g2_buf_1 _15804_ (.A(net681),
    .X(_09092_));
 sg13g2_buf_1 _15805_ (.A(net619),
    .X(_09093_));
 sg13g2_buf_1 _15806_ (.A(net552),
    .X(_09094_));
 sg13g2_nor3_2 _15807_ (.A(net1036),
    .B(net620),
    .C(net496),
    .Y(_09095_));
 sg13g2_nand3b_1 _15808_ (.B(_09078_),
    .C(_09095_),
    .Y(_09096_),
    .A_N(_00197_));
 sg13g2_inv_1 _15809_ (.Y(_09097_),
    .A(_08768_));
 sg13g2_buf_1 _15810_ (.A(_08767_),
    .X(_09098_));
 sg13g2_nand2_1 _15811_ (.Y(_09099_),
    .A(net1032),
    .B(_08765_));
 sg13g2_o21ai_1 _15812_ (.B1(_09099_),
    .Y(_09100_),
    .A1(net1032),
    .A2(net1110));
 sg13g2_nand2_1 _15813_ (.Y(_09101_),
    .A(net1110),
    .B(_08766_));
 sg13g2_o21ai_1 _15814_ (.B1(_09101_),
    .Y(_09102_),
    .A1(net1033),
    .A2(_09100_));
 sg13g2_buf_1 _15815_ (.A(_09102_),
    .X(_09103_));
 sg13g2_nor3_2 _15816_ (.A(_09017_),
    .B(_09096_),
    .C(_09103_),
    .Y(_09104_));
 sg13g2_buf_2 _15817_ (.A(\cpu.spi.r_state[1] ),
    .X(_09105_));
 sg13g2_inv_2 _15818_ (.Y(_09106_),
    .A(_09105_));
 sg13g2_buf_1 _15819_ (.A(_08776_),
    .X(_09107_));
 sg13g2_nand3_1 _15820_ (.B(_09021_),
    .C(_09078_),
    .A(net1031),
    .Y(_09108_));
 sg13g2_buf_2 _15821_ (.A(_09108_),
    .X(_09109_));
 sg13g2_or2_1 _15822_ (.X(_09110_),
    .B(_09109_),
    .A(_09017_));
 sg13g2_buf_1 _15823_ (.A(_09110_),
    .X(_09111_));
 sg13g2_nor2_1 _15824_ (.A(net496),
    .B(_09111_),
    .Y(_09112_));
 sg13g2_buf_1 _15825_ (.A(_09112_),
    .X(_09113_));
 sg13g2_nor2_1 _15826_ (.A(_09106_),
    .B(_09113_),
    .Y(_09114_));
 sg13g2_a21oi_1 _15827_ (.A1(_09104_),
    .A2(_09114_),
    .Y(_09115_),
    .B1(\cpu.spi.r_state[3] ));
 sg13g2_buf_2 _15828_ (.A(\cpu.spi.r_state[0] ),
    .X(_09116_));
 sg13g2_buf_1 _15829_ (.A(net1036),
    .X(_09117_));
 sg13g2_buf_1 _15830_ (.A(net898),
    .X(_09118_));
 sg13g2_buf_2 _15831_ (.A(net620),
    .X(_09119_));
 sg13g2_nor2_1 _15832_ (.A(net782),
    .B(net551),
    .Y(_09120_));
 sg13g2_nand2_2 _15833_ (.Y(_09121_),
    .A(_09120_),
    .B(_09113_));
 sg13g2_nand2b_1 _15834_ (.Y(_09122_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _15835_ (.A(_09122_),
    .X(_09123_));
 sg13g2_a21oi_2 _15836_ (.B1(net1030),
    .Y(_09124_),
    .A2(_09121_),
    .A1(_09116_));
 sg13g2_o21ai_1 _15837_ (.B1(_09124_),
    .Y(_00029_),
    .A1(_09009_),
    .A2(_09115_));
 sg13g2_nor2b_1 _15838_ (.A(r_reset),
    .B_N(net1),
    .Y(_09125_));
 sg13g2_buf_1 _15839_ (.A(_09125_),
    .X(_09126_));
 sg13g2_buf_1 _15840_ (.A(_09126_),
    .X(_09127_));
 sg13g2_buf_1 _15841_ (.A(_09127_),
    .X(_09128_));
 sg13g2_buf_1 _15842_ (.A(net781),
    .X(_09129_));
 sg13g2_inv_2 _15843_ (.Y(_09130_),
    .A(net1034));
 sg13g2_buf_1 _15844_ (.A(_09130_),
    .X(_09131_));
 sg13g2_nor2_1 _15845_ (.A(_09017_),
    .B(_09109_),
    .Y(_09132_));
 sg13g2_buf_1 _15846_ (.A(_09132_),
    .X(_09133_));
 sg13g2_nand2_2 _15847_ (.Y(_09134_),
    .A(net780),
    .B(_09133_));
 sg13g2_nand2_1 _15848_ (.Y(_09135_),
    .A(_09105_),
    .B(_09134_));
 sg13g2_buf_1 _15849_ (.A(\cpu.spi.r_state[6] ),
    .X(_09136_));
 sg13g2_buf_1 _15850_ (.A(_09136_),
    .X(_09137_));
 sg13g2_nor2b_1 _15851_ (.A(_08999_),
    .B_N(_09007_),
    .Y(_09138_));
 sg13g2_buf_1 _15852_ (.A(_09138_),
    .X(_09139_));
 sg13g2_buf_1 _15853_ (.A(_09139_),
    .X(_09140_));
 sg13g2_buf_1 _15854_ (.A(net377),
    .X(_09141_));
 sg13g2_buf_1 _15855_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09142_));
 sg13g2_buf_1 _15856_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09143_));
 sg13g2_nor3_1 _15857_ (.A(_09142_),
    .B(_09143_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09144_));
 sg13g2_buf_1 _15858_ (.A(\cpu.spi.r_timeout_count[7] ),
    .X(_09145_));
 sg13g2_buf_1 _15859_ (.A(\cpu.spi.r_timeout_count[0] ),
    .X(_09146_));
 sg13g2_buf_1 _15860_ (.A(\cpu.spi.r_timeout_count[1] ),
    .X(_09147_));
 sg13g2_or3_1 _15861_ (.A(_09146_),
    .B(_09147_),
    .C(\cpu.spi.r_timeout_count[2] ),
    .X(_09148_));
 sg13g2_buf_1 _15862_ (.A(_09148_),
    .X(_09149_));
 sg13g2_or2_1 _15863_ (.X(_09150_),
    .B(_09149_),
    .A(\cpu.spi.r_timeout_count[3] ));
 sg13g2_buf_1 _15864_ (.A(_09150_),
    .X(_09151_));
 sg13g2_or2_1 _15865_ (.X(_09152_),
    .B(_09151_),
    .A(\cpu.spi.r_timeout_count[4] ));
 sg13g2_buf_1 _15866_ (.A(_09152_),
    .X(_09153_));
 sg13g2_or2_1 _15867_ (.X(_09154_),
    .B(_09153_),
    .A(\cpu.spi.r_timeout_count[5] ));
 sg13g2_buf_1 _15868_ (.A(_09154_),
    .X(_09155_));
 sg13g2_or2_1 _15869_ (.X(_09156_),
    .B(_09155_),
    .A(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _15870_ (.A(_09156_),
    .X(_09157_));
 sg13g2_o21ai_1 _15871_ (.B1(\cpu.spi.r_searching ),
    .Y(_09158_),
    .A1(_09145_),
    .A2(_09157_));
 sg13g2_nand2_1 _15872_ (.Y(_09159_),
    .A(_09144_),
    .B(_09158_));
 sg13g2_buf_1 _15873_ (.A(\cpu.spi.r_in[3] ),
    .X(_09160_));
 sg13g2_buf_1 _15874_ (.A(\cpu.spi.r_in[6] ),
    .X(_09161_));
 sg13g2_buf_1 _15875_ (.A(\cpu.spi.r_in[1] ),
    .X(_09162_));
 sg13g2_buf_1 _15876_ (.A(\cpu.spi.r_in[0] ),
    .X(_09163_));
 sg13g2_nand2_1 _15877_ (.Y(_09164_),
    .A(_09162_),
    .B(_09163_));
 sg13g2_nand3_1 _15878_ (.B(_09161_),
    .C(_09164_),
    .A(_09160_),
    .Y(_09165_));
 sg13g2_buf_1 _15879_ (.A(\cpu.spi.r_in[2] ),
    .X(_09166_));
 sg13g2_buf_1 _15880_ (.A(\cpu.spi.r_in[5] ),
    .X(_09167_));
 sg13g2_buf_1 _15881_ (.A(\cpu.spi.r_in[4] ),
    .X(_09168_));
 sg13g2_nand4_1 _15882_ (.B(_09167_),
    .C(_09168_),
    .A(_09166_),
    .Y(_09169_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _15883_ (.A(_09165_),
    .B(_09169_),
    .Y(_09170_));
 sg13g2_o21ai_1 _15884_ (.B1(\cpu.spi.r_searching ),
    .Y(_09171_),
    .A1(_00222_),
    .A2(_09170_));
 sg13g2_nand2_1 _15885_ (.Y(_09172_),
    .A(_09159_),
    .B(_09171_));
 sg13g2_nand3_1 _15886_ (.B(net345),
    .C(_09172_),
    .A(net1029),
    .Y(_09173_));
 sg13g2_o21ai_1 _15887_ (.B1(_09173_),
    .Y(_09174_),
    .A1(_09104_),
    .A2(_09135_));
 sg13g2_and2_1 _15888_ (.A(net680),
    .B(_09174_),
    .X(_00030_));
 sg13g2_nand4_1 _15889_ (.B(net377),
    .C(_09159_),
    .A(net1029),
    .Y(_09175_),
    .D(_09171_));
 sg13g2_buf_1 _15890_ (.A(\cpu.spi.r_state[2] ),
    .X(_09176_));
 sg13g2_buf_1 _15891_ (.A(\cpu.spi.r_state[4] ),
    .X(_09177_));
 sg13g2_nor3_1 _15892_ (.A(\cpu.spi.r_state[5] ),
    .B(net1104),
    .C(_09009_),
    .Y(_09178_));
 sg13g2_o21ai_1 _15893_ (.B1(_09178_),
    .Y(_09179_),
    .A1(_09106_),
    .A2(_09134_));
 sg13g2_o21ai_1 _15894_ (.B1(_09179_),
    .Y(_09180_),
    .A1(net1105),
    .A2(net345));
 sg13g2_buf_2 _15895_ (.A(net1030),
    .X(_09181_));
 sg13g2_buf_1 _15896_ (.A(net896),
    .X(_09182_));
 sg13g2_buf_2 _15897_ (.A(net779),
    .X(_09183_));
 sg13g2_buf_1 _15898_ (.A(_09183_),
    .X(_09184_));
 sg13g2_a21oi_1 _15899_ (.A1(_09175_),
    .A2(_09180_),
    .Y(_00031_),
    .B1(net618));
 sg13g2_buf_1 _15900_ (.A(net779),
    .X(_09185_));
 sg13g2_nor3_1 _15901_ (.A(net679),
    .B(net345),
    .C(_09115_),
    .Y(_00032_));
 sg13g2_buf_1 _15902_ (.A(net779),
    .X(_09186_));
 sg13g2_buf_1 _15903_ (.A(_09186_),
    .X(_09187_));
 sg13g2_inv_1 _15904_ (.Y(_09188_),
    .A(_09121_));
 sg13g2_a22oi_1 _15905_ (.Y(_09189_),
    .B1(_09009_),
    .B2(net1104),
    .A2(_09188_),
    .A1(_09116_));
 sg13g2_nor2_1 _15906_ (.A(net617),
    .B(_09189_),
    .Y(_00033_));
 sg13g2_buf_1 _15907_ (.A(_09105_),
    .X(_09190_));
 sg13g2_buf_1 _15908_ (.A(_09113_),
    .X(_09191_));
 sg13g2_buf_1 _15909_ (.A(net80),
    .X(_09192_));
 sg13g2_a21oi_1 _15910_ (.A1(_09190_),
    .A2(net70),
    .Y(_09193_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_nor3_1 _15911_ (.A(net679),
    .B(_09141_),
    .C(_09193_),
    .Y(_00034_));
 sg13g2_and2_1 _15912_ (.A(_09136_),
    .B(_09009_),
    .X(_09194_));
 sg13g2_a21oi_1 _15913_ (.A1(net1105),
    .A2(_09141_),
    .Y(_09195_),
    .B1(_09194_));
 sg13g2_nor2_1 _15914_ (.A(net617),
    .B(_09195_),
    .Y(_00035_));
 sg13g2_buf_1 _15915_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09196_));
 sg13g2_buf_1 _15916_ (.A(\cpu.dec.mult ),
    .X(_09197_));
 sg13g2_inv_1 _15917_ (.Y(_09198_),
    .A(_09197_));
 sg13g2_nand3b_1 _15918_ (.B(\cpu.dec.iready ),
    .C(_00199_),
    .Y(_09199_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_1 _15919_ (.A(_09199_),
    .X(_09200_));
 sg13g2_nor3_2 _15920_ (.A(_09198_),
    .B(net1030),
    .C(net1027),
    .Y(_09201_));
 sg13g2_buf_1 _15921_ (.A(\cpu.dec.div ),
    .X(_09202_));
 sg13g2_inv_1 _15922_ (.Y(_09203_),
    .A(_09202_));
 sg13g2_nor3_1 _15923_ (.A(_09203_),
    .B(net1030),
    .C(net1027),
    .Y(_09204_));
 sg13g2_buf_2 _15924_ (.A(_09204_),
    .X(_09205_));
 sg13g2_nor2_1 _15925_ (.A(_09201_),
    .B(_09205_),
    .Y(_09206_));
 sg13g2_buf_2 _15926_ (.A(_09206_),
    .X(_09207_));
 sg13g2_nand2_1 _15927_ (.Y(_09208_),
    .A(_09196_),
    .B(_09207_));
 sg13g2_buf_1 _15928_ (.A(_09208_),
    .X(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _15929_ (.A(\cpu.ex.r_div_running ),
    .X(_09209_));
 sg13g2_buf_1 _15930_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09210_));
 sg13g2_nor4_2 _15931_ (.A(_09210_),
    .B(\cpu.ex.r_mult_off[2] ),
    .C(\cpu.ex.r_mult_off[3] ),
    .Y(_09211_),
    .D(net495));
 sg13g2_buf_1 _15932_ (.A(_09205_),
    .X(_09212_));
 sg13g2_buf_1 _15933_ (.A(_09212_),
    .X(_09213_));
 sg13g2_o21ai_1 _15934_ (.B1(_09126_),
    .Y(_09214_),
    .A1(_09209_),
    .A2(net616));
 sg13g2_a21oi_1 _15935_ (.A1(_09209_),
    .A2(_09211_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09214_));
 sg13g2_buf_1 _15936_ (.A(\cpu.ex.r_mult_running ),
    .X(_09215_));
 sg13g2_inv_1 _15937_ (.Y(_09216_),
    .A(net1103));
 sg13g2_nor2_1 _15938_ (.A(net1030),
    .B(net1027),
    .Y(_09217_));
 sg13g2_nand2_1 _15939_ (.Y(_09218_),
    .A(_09197_),
    .B(_09217_));
 sg13g2_buf_1 _15940_ (.A(_09218_),
    .X(_09219_));
 sg13g2_nand2_1 _15941_ (.Y(_09220_),
    .A(_09216_),
    .B(net677));
 sg13g2_buf_2 _15942_ (.A(_09220_),
    .X(_09221_));
 sg13g2_nand2_1 _15943_ (.Y(_09222_),
    .A(_09126_),
    .B(_09221_));
 sg13g2_a21oi_1 _15944_ (.A1(net1103),
    .A2(_09211_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09222_));
 sg13g2_buf_2 _15945_ (.A(\cpu.dcache.flush_write ),
    .X(_09223_));
 sg13g2_buf_4 _15946_ (.X(_09224_),
    .A(_08754_));
 sg13g2_buf_2 _15947_ (.A(_09224_),
    .X(_09225_));
 sg13g2_buf_2 _15948_ (.A(_08751_),
    .X(_09226_));
 sg13g2_buf_1 _15949_ (.A(_09226_),
    .X(_09227_));
 sg13g2_buf_1 _15950_ (.A(net777),
    .X(_09228_));
 sg13g2_mux4_1 _15951_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net676),
    .X(_09229_));
 sg13g2_buf_8 _15952_ (.A(_09224_),
    .X(_09230_));
 sg13g2_buf_2 _15953_ (.A(net776),
    .X(_09231_));
 sg13g2_mux4_1 _15954_ (.S0(net675),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net676),
    .X(_09232_));
 sg13g2_buf_1 _15955_ (.A(_08751_),
    .X(_09233_));
 sg13g2_buf_2 _15956_ (.A(net895),
    .X(_09234_));
 sg13g2_mux4_1 _15957_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net775),
    .X(_09235_));
 sg13g2_mux4_1 _15958_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(net775),
    .X(_09236_));
 sg13g2_buf_2 _15959_ (.A(net902),
    .X(_09237_));
 sg13g2_buf_1 _15960_ (.A(net1112),
    .X(_09238_));
 sg13g2_mux4_1 _15961_ (.S0(net774),
    .A0(_09229_),
    .A1(_09232_),
    .A2(_09235_),
    .A3(_09236_),
    .S1(net1026),
    .X(_09239_));
 sg13g2_mux4_1 _15962_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(net676),
    .X(_09240_));
 sg13g2_mux4_1 _15963_ (.S0(_09225_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net676),
    .X(_09241_));
 sg13g2_mux4_1 _15964_ (.S0(_09225_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(_09234_),
    .X(_09242_));
 sg13g2_mux4_1 _15965_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(_09234_),
    .X(_09243_));
 sg13g2_mux4_1 _15966_ (.S0(_09237_),
    .A0(_09240_),
    .A1(_09241_),
    .A2(_09242_),
    .A3(_09243_),
    .S1(net1026),
    .X(_09244_));
 sg13g2_buf_1 _15967_ (.A(_08740_),
    .X(_09245_));
 sg13g2_mux2_1 _15968_ (.A0(_09239_),
    .A1(_09244_),
    .S(net674),
    .X(_09246_));
 sg13g2_nand2_1 _15969_ (.Y(_09247_),
    .A(net1053),
    .B(_09246_));
 sg13g2_o21ai_1 _15970_ (.B1(_09247_),
    .Y(_09248_),
    .A1(_08365_),
    .A2(_08822_));
 sg13g2_buf_1 _15971_ (.A(_09248_),
    .X(_09249_));
 sg13g2_buf_2 _15972_ (.A(_00227_),
    .X(_09250_));
 sg13g2_buf_1 _15973_ (.A(_09250_),
    .X(_09251_));
 sg13g2_inv_2 _15974_ (.Y(_09252_),
    .A(_09081_));
 sg13g2_nand2_1 _15975_ (.Y(_09253_),
    .A(_09252_),
    .B(_09130_));
 sg13g2_buf_1 _15976_ (.A(\cpu.addr[4] ),
    .X(_09254_));
 sg13g2_buf_1 _15977_ (.A(_09254_),
    .X(_09255_));
 sg13g2_a21oi_1 _15978_ (.A1(net1025),
    .A2(_09253_),
    .Y(_09256_),
    .B1(net1024));
 sg13g2_buf_1 _15979_ (.A(_09256_),
    .X(_09257_));
 sg13g2_buf_1 _15980_ (.A(net615),
    .X(_09258_));
 sg13g2_a21o_1 _15981_ (.A2(_09253_),
    .A1(_09250_),
    .B1(net1024),
    .X(_09259_));
 sg13g2_buf_2 _15982_ (.A(_09259_),
    .X(_09260_));
 sg13g2_buf_1 _15983_ (.A(_09260_),
    .X(_09261_));
 sg13g2_buf_1 _15984_ (.A(net549),
    .X(_09262_));
 sg13g2_nor2b_1 _15985_ (.A(_09081_),
    .B_N(_09087_),
    .Y(_09263_));
 sg13g2_buf_1 _15986_ (.A(_09263_),
    .X(_09264_));
 sg13g2_and2_1 _15987_ (.A(_09250_),
    .B(_09264_),
    .X(_09265_));
 sg13g2_buf_1 _15988_ (.A(_09265_),
    .X(_09266_));
 sg13g2_buf_1 _15989_ (.A(_09266_),
    .X(_09267_));
 sg13g2_buf_1 _15990_ (.A(net614),
    .X(_09268_));
 sg13g2_nor2b_1 _15991_ (.A(net1034),
    .B_N(_09081_),
    .Y(_09269_));
 sg13g2_buf_1 _15992_ (.A(_09269_),
    .X(_09270_));
 sg13g2_and2_1 _15993_ (.A(_09250_),
    .B(_09270_),
    .X(_09271_));
 sg13g2_buf_2 _15994_ (.A(_09271_),
    .X(_09272_));
 sg13g2_buf_1 _15995_ (.A(_09272_),
    .X(_09273_));
 sg13g2_buf_1 _15996_ (.A(net547),
    .X(_09274_));
 sg13g2_a22oi_1 _15997_ (.Y(_09275_),
    .B1(net493),
    .B2(\cpu.dcache.r_tag[1][12] ),
    .A2(net548),
    .A1(\cpu.dcache.r_tag[2][12] ));
 sg13g2_and2_1 _15998_ (.A(_09081_),
    .B(_09087_),
    .X(_09276_));
 sg13g2_buf_1 _15999_ (.A(_09276_),
    .X(_09277_));
 sg13g2_and2_1 _16000_ (.A(_09250_),
    .B(_09277_),
    .X(_09278_));
 sg13g2_buf_1 _16001_ (.A(_09278_),
    .X(_09279_));
 sg13g2_buf_1 _16002_ (.A(_09279_),
    .X(_09280_));
 sg13g2_buf_1 _16003_ (.A(net613),
    .X(_09281_));
 sg13g2_nor2b_1 _16004_ (.A(_09081_),
    .B_N(_09254_),
    .Y(_09282_));
 sg13g2_buf_1 _16005_ (.A(_09282_),
    .X(_09283_));
 sg13g2_and2_1 _16006_ (.A(net1034),
    .B(_09283_),
    .X(_09284_));
 sg13g2_buf_2 _16007_ (.A(_09284_),
    .X(_09285_));
 sg13g2_buf_1 _16008_ (.A(_09285_),
    .X(_09286_));
 sg13g2_a22oi_1 _16009_ (.Y(_09287_),
    .B1(net612),
    .B2(\cpu.dcache.r_tag[6][12] ),
    .A2(net546),
    .A1(\cpu.dcache.r_tag[3][12] ));
 sg13g2_nor2_1 _16010_ (.A(_09081_),
    .B(net1034),
    .Y(_09288_));
 sg13g2_buf_1 _16011_ (.A(_09288_),
    .X(_09289_));
 sg13g2_buf_1 _16012_ (.A(_09289_),
    .X(_09290_));
 sg13g2_mux2_1 _16013_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(\cpu.dcache.r_tag[7][12] ),
    .S(net783),
    .X(_09291_));
 sg13g2_a22oi_1 _16014_ (.Y(_09292_),
    .B1(_09291_),
    .B2(_09084_),
    .A2(net673),
    .A1(\cpu.dcache.r_tag[4][12] ));
 sg13g2_buf_1 _16015_ (.A(net1024),
    .X(_09293_));
 sg13g2_buf_1 _16016_ (.A(net893),
    .X(_09294_));
 sg13g2_nand2b_1 _16017_ (.Y(_09295_),
    .B(_09294_),
    .A_N(_09292_));
 sg13g2_and4_1 _16018_ (.A(net494),
    .B(_09275_),
    .C(_09287_),
    .D(_09295_),
    .X(_09296_));
 sg13g2_a21oi_1 _16019_ (.A1(_00243_),
    .A2(_09258_),
    .Y(_09297_),
    .B1(_09296_));
 sg13g2_xnor2_1 _16020_ (.Y(_09298_),
    .A(net344),
    .B(_09297_));
 sg13g2_mux4_1 _16021_ (.S0(net675),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(_09228_),
    .X(_09299_));
 sg13g2_mux4_1 _16022_ (.S0(net675),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(_09228_),
    .X(_09300_));
 sg13g2_mux4_1 _16023_ (.S0(net675),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(net676),
    .X(_09301_));
 sg13g2_mux4_1 _16024_ (.S0(_09231_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(net676),
    .X(_09302_));
 sg13g2_mux4_1 _16025_ (.S0(net774),
    .A0(_09299_),
    .A1(_09300_),
    .A2(_09301_),
    .A3(_09302_),
    .S1(net1026),
    .X(_09303_));
 sg13g2_mux4_1 _16026_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net775),
    .X(_09304_));
 sg13g2_mux4_1 _16027_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(net775),
    .X(_09305_));
 sg13g2_buf_2 _16028_ (.A(_09224_),
    .X(_09306_));
 sg13g2_buf_2 _16029_ (.A(_09226_),
    .X(_09307_));
 sg13g2_mux4_1 _16030_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net770),
    .X(_09308_));
 sg13g2_mux4_1 _16031_ (.S0(_09306_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net770),
    .X(_09309_));
 sg13g2_mux4_1 _16032_ (.S0(_09237_),
    .A0(_09304_),
    .A1(_09305_),
    .A2(_09308_),
    .A3(_09309_),
    .S1(net1026),
    .X(_09310_));
 sg13g2_and2_1 _16033_ (.A(net683),
    .B(_09310_),
    .X(_09311_));
 sg13g2_a21oi_1 _16034_ (.A1(net674),
    .A2(_09303_),
    .Y(_09312_),
    .B1(_09311_));
 sg13g2_buf_1 _16035_ (.A(net676),
    .X(_09313_));
 sg13g2_nor2_1 _16036_ (.A(net1115),
    .B(net611),
    .Y(_09314_));
 sg13g2_a21oi_1 _16037_ (.A1(_08365_),
    .A2(_09312_),
    .Y(_09315_),
    .B1(_09314_));
 sg13g2_buf_1 _16038_ (.A(_09315_),
    .X(_09316_));
 sg13g2_a22oi_1 _16039_ (.Y(_09317_),
    .B1(net493),
    .B2(\cpu.dcache.r_tag[1][13] ),
    .A2(net548),
    .A1(\cpu.dcache.r_tag[2][13] ));
 sg13g2_a22oi_1 _16040_ (.Y(_09318_),
    .B1(_09286_),
    .B2(\cpu.dcache.r_tag[6][13] ),
    .A2(net546),
    .A1(\cpu.dcache.r_tag[3][13] ));
 sg13g2_mux2_1 _16041_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(\cpu.dcache.r_tag[7][13] ),
    .S(net783),
    .X(_09319_));
 sg13g2_a22oi_1 _16042_ (.Y(_09320_),
    .B1(_09319_),
    .B2(net900),
    .A2(net673),
    .A1(\cpu.dcache.r_tag[4][13] ));
 sg13g2_nand2b_1 _16043_ (.Y(_09321_),
    .B(net772),
    .A_N(_09320_));
 sg13g2_and4_1 _16044_ (.A(net494),
    .B(_09317_),
    .C(_09318_),
    .D(_09321_),
    .X(_09322_));
 sg13g2_a21oi_1 _16045_ (.A1(_00244_),
    .A2(_09258_),
    .Y(_09323_),
    .B1(_09322_));
 sg13g2_xnor2_1 _16046_ (.Y(_09324_),
    .A(net376),
    .B(_09323_));
 sg13g2_buf_2 _16047_ (.A(_09224_),
    .X(_09325_));
 sg13g2_mux4_1 _16048_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net770),
    .X(_09326_));
 sg13g2_mux4_1 _16049_ (.S0(_09306_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net770),
    .X(_09327_));
 sg13g2_buf_2 _16050_ (.A(_09226_),
    .X(_09328_));
 sg13g2_mux4_1 _16051_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net768),
    .X(_09329_));
 sg13g2_mux4_1 _16052_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net768),
    .X(_09330_));
 sg13g2_buf_2 _16053_ (.A(net902),
    .X(_09331_));
 sg13g2_mux4_1 _16054_ (.S0(net767),
    .A0(_09326_),
    .A1(_09327_),
    .A2(_09329_),
    .A3(_09330_),
    .S1(_09238_),
    .X(_09332_));
 sg13g2_nand2_1 _16055_ (.Y(_09333_),
    .A(_08832_),
    .B(_09332_));
 sg13g2_mux4_1 _16056_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(_09307_),
    .X(_09334_));
 sg13g2_mux4_1 _16057_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(_09307_),
    .X(_09335_));
 sg13g2_buf_2 _16058_ (.A(_09224_),
    .X(_09336_));
 sg13g2_mux4_1 _16059_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net768),
    .X(_09337_));
 sg13g2_mux4_1 _16060_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(_09328_),
    .X(_09338_));
 sg13g2_mux4_1 _16061_ (.S0(net767),
    .A0(_09334_),
    .A1(_09335_),
    .A2(_09337_),
    .A3(_09338_),
    .S1(_09238_),
    .X(_09339_));
 sg13g2_nand2_1 _16062_ (.Y(_09340_),
    .A(net674),
    .B(_09339_));
 sg13g2_a21oi_2 _16063_ (.B1(_08436_),
    .Y(_09341_),
    .A2(_09340_),
    .A1(_09333_));
 sg13g2_buf_1 _16064_ (.A(_09341_),
    .X(_09342_));
 sg13g2_inv_1 _16065_ (.Y(_09343_),
    .A(_00249_));
 sg13g2_and2_1 _16066_ (.A(_09254_),
    .B(net773),
    .X(_09344_));
 sg13g2_buf_2 _16067_ (.A(_09344_),
    .X(_09345_));
 sg13g2_buf_1 _16068_ (.A(_09345_),
    .X(_09346_));
 sg13g2_a22oi_1 _16069_ (.Y(_09347_),
    .B1(net545),
    .B2(\cpu.dcache.r_tag[5][18] ),
    .A2(net493),
    .A1(\cpu.dcache.r_tag[1][18] ));
 sg13g2_a22oi_1 _16070_ (.Y(_09348_),
    .B1(net546),
    .B2(\cpu.dcache.r_tag[3][18] ),
    .A2(net548),
    .A1(\cpu.dcache.r_tag[2][18] ));
 sg13g2_buf_1 _16071_ (.A(_09277_),
    .X(_09349_));
 sg13g2_mux2_1 _16072_ (.A0(\cpu.dcache.r_tag[4][18] ),
    .A1(\cpu.dcache.r_tag[6][18] ),
    .S(net899),
    .X(_09350_));
 sg13g2_buf_1 _16073_ (.A(_09252_),
    .X(_09351_));
 sg13g2_a22oi_1 _16074_ (.Y(_09352_),
    .B1(_09350_),
    .B2(net892),
    .A2(net765),
    .A1(\cpu.dcache.r_tag[7][18] ));
 sg13g2_nand2b_1 _16075_ (.Y(_09353_),
    .B(net893),
    .A_N(_09352_));
 sg13g2_nand4_1 _16076_ (.B(_09347_),
    .C(_09348_),
    .A(_09262_),
    .Y(_09354_),
    .D(_09353_));
 sg13g2_o21ai_1 _16077_ (.B1(_09354_),
    .Y(_09355_),
    .A1(_09343_),
    .A2(net494));
 sg13g2_xnor2_1 _16078_ (.Y(_09356_),
    .A(net439),
    .B(_09355_));
 sg13g2_inv_1 _16079_ (.Y(_09357_),
    .A(_00237_));
 sg13g2_inv_1 _16080_ (.Y(_09358_),
    .A(_09254_));
 sg13g2_buf_1 _16081_ (.A(_09358_),
    .X(_09359_));
 sg13g2_mux2_1 _16082_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(\cpu.dcache.r_tag[7][9] ),
    .S(net783),
    .X(_09360_));
 sg13g2_a22oi_1 _16083_ (.Y(_09361_),
    .B1(_09360_),
    .B2(net900),
    .A2(net673),
    .A1(\cpu.dcache.r_tag[4][9] ));
 sg13g2_a22oi_1 _16084_ (.Y(_09362_),
    .B1(\cpu.dcache.r_tag[2][9] ),
    .B2(net1025),
    .A2(\cpu.dcache.r_tag[6][9] ),
    .A1(_09255_));
 sg13g2_nand3_1 _16085_ (.B(net1025),
    .C(\cpu.dcache.r_tag[3][9] ),
    .A(net1035),
    .Y(_09363_));
 sg13g2_o21ai_1 _16086_ (.B1(_09363_),
    .Y(_09364_),
    .A1(net900),
    .A2(_09362_));
 sg13g2_a22oi_1 _16087_ (.Y(_09365_),
    .B1(_09364_),
    .B2(net783),
    .A2(net547),
    .A1(\cpu.dcache.r_tag[1][9] ));
 sg13g2_o21ai_1 _16088_ (.B1(_09365_),
    .Y(_09366_),
    .A1(net891),
    .A2(_09361_));
 sg13g2_nand2b_1 _16089_ (.Y(_09367_),
    .B(net615),
    .A_N(_00238_));
 sg13g2_nand2b_1 _16090_ (.Y(_09368_),
    .B(_09367_),
    .A_N(_09366_));
 sg13g2_xnor2_1 _16091_ (.Y(_09369_),
    .A(_09357_),
    .B(_09368_));
 sg13g2_mux2_1 _16092_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(\cpu.dcache.r_tag[7][8] ),
    .S(_09090_),
    .X(_09370_));
 sg13g2_a22oi_1 _16093_ (.Y(_09371_),
    .B1(_09370_),
    .B2(net900),
    .A2(net673),
    .A1(\cpu.dcache.r_tag[4][8] ));
 sg13g2_inv_1 _16094_ (.Y(_09372_),
    .A(_00236_));
 sg13g2_a22oi_1 _16095_ (.Y(_09373_),
    .B1(\cpu.dcache.r_tag[2][8] ),
    .B2(_09250_),
    .A2(\cpu.dcache.r_tag[6][8] ),
    .A1(net1024));
 sg13g2_nand3_1 _16096_ (.B(_09250_),
    .C(\cpu.dcache.r_tag[3][8] ),
    .A(net1035),
    .Y(_09374_));
 sg13g2_o21ai_1 _16097_ (.B1(_09374_),
    .Y(_09375_),
    .A1(net1035),
    .A2(_09373_));
 sg13g2_and2_1 _16098_ (.A(net783),
    .B(_09375_),
    .X(_09376_));
 sg13g2_a221oi_1 _16099_ (.B2(\cpu.dcache.r_tag[1][8] ),
    .C1(_09376_),
    .B1(net493),
    .A1(_09372_),
    .Y(_09377_),
    .A2(_09256_));
 sg13g2_o21ai_1 _16100_ (.B1(_09377_),
    .Y(_09378_),
    .A1(net891),
    .A2(_09371_));
 sg13g2_xor2_1 _16101_ (.B(_09378_),
    .A(_00235_),
    .X(_09379_));
 sg13g2_a22oi_1 _16102_ (.Y(_09380_),
    .B1(net547),
    .B2(\cpu.dcache.r_tag[1][7] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][7] ));
 sg13g2_a22oi_1 _16103_ (.Y(_09381_),
    .B1(_09285_),
    .B2(\cpu.dcache.r_tag[6][7] ),
    .A2(net613),
    .A1(\cpu.dcache.r_tag[3][7] ));
 sg13g2_mux2_1 _16104_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(\cpu.dcache.r_tag[7][7] ),
    .S(net1034),
    .X(_09382_));
 sg13g2_a22oi_1 _16105_ (.Y(_09383_),
    .B1(_09382_),
    .B2(net1035),
    .A2(_09289_),
    .A1(\cpu.dcache.r_tag[4][7] ));
 sg13g2_nand2b_1 _16106_ (.Y(_09384_),
    .B(net1024),
    .A_N(_09383_));
 sg13g2_and4_1 _16107_ (.A(_09260_),
    .B(_09380_),
    .C(_09381_),
    .D(_09384_),
    .X(_09385_));
 sg13g2_a21oi_1 _16108_ (.A1(_00234_),
    .A2(net615),
    .Y(_09386_),
    .B1(_09385_));
 sg13g2_xor2_1 _16109_ (.B(_09386_),
    .A(_00233_),
    .X(_09387_));
 sg13g2_nand3_1 _16110_ (.B(_09379_),
    .C(_09387_),
    .A(_09369_),
    .Y(_09388_));
 sg13g2_buf_2 _16111_ (.A(_00229_),
    .X(_09389_));
 sg13g2_and2_1 _16112_ (.A(net1024),
    .B(net765),
    .X(_09390_));
 sg13g2_buf_1 _16113_ (.A(_09390_),
    .X(_09391_));
 sg13g2_a22oi_1 _16114_ (.Y(_09392_),
    .B1(_09391_),
    .B2(\cpu.dcache.r_tag[7][5] ),
    .A2(_09285_),
    .A1(\cpu.dcache.r_tag[6][5] ));
 sg13g2_and2_1 _16115_ (.A(_09130_),
    .B(_09283_),
    .X(_09393_));
 sg13g2_buf_2 _16116_ (.A(_09393_),
    .X(_09394_));
 sg13g2_a22oi_1 _16117_ (.Y(_09395_),
    .B1(_09345_),
    .B2(\cpu.dcache.r_tag[5][5] ),
    .A2(_09394_),
    .A1(\cpu.dcache.r_tag[4][5] ));
 sg13g2_mux2_1 _16118_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(\cpu.dcache.r_tag[3][5] ),
    .S(_09088_),
    .X(_09396_));
 sg13g2_a22oi_1 _16119_ (.Y(_09397_),
    .B1(_09396_),
    .B2(net1035),
    .A2(net894),
    .A1(\cpu.dcache.r_tag[2][5] ));
 sg13g2_nand2b_1 _16120_ (.Y(_09398_),
    .B(_09251_),
    .A_N(_09397_));
 sg13g2_and4_1 _16121_ (.A(_09260_),
    .B(_09392_),
    .C(_09395_),
    .D(_09398_),
    .X(_09399_));
 sg13g2_a21oi_1 _16122_ (.A1(_00230_),
    .A2(net615),
    .Y(_09400_),
    .B1(_09399_));
 sg13g2_xnor2_1 _16123_ (.Y(_09401_),
    .A(_09389_),
    .B(_09400_));
 sg13g2_a22oi_1 _16124_ (.Y(_09402_),
    .B1(_09272_),
    .B2(\cpu.dcache.r_tag[1][10] ),
    .A2(_09266_),
    .A1(\cpu.dcache.r_tag[2][10] ));
 sg13g2_a22oi_1 _16125_ (.Y(_09403_),
    .B1(_09285_),
    .B2(\cpu.dcache.r_tag[6][10] ),
    .A2(_09279_),
    .A1(\cpu.dcache.r_tag[3][10] ));
 sg13g2_mux2_1 _16126_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(\cpu.dcache.r_tag[7][10] ),
    .S(net1034),
    .X(_09404_));
 sg13g2_a22oi_1 _16127_ (.Y(_09405_),
    .B1(_09404_),
    .B2(net1035),
    .A2(_09289_),
    .A1(\cpu.dcache.r_tag[4][10] ));
 sg13g2_nand2b_1 _16128_ (.Y(_09406_),
    .B(net1024),
    .A_N(_09405_));
 sg13g2_and4_1 _16129_ (.A(_09260_),
    .B(_09402_),
    .C(_09403_),
    .D(_09406_),
    .X(_09407_));
 sg13g2_a21oi_1 _16130_ (.A1(_00240_),
    .A2(net615),
    .Y(_09408_),
    .B1(_09407_));
 sg13g2_xnor2_1 _16131_ (.Y(_09409_),
    .A(_00239_),
    .B(_09408_));
 sg13g2_a22oi_1 _16132_ (.Y(_09410_),
    .B1(_09272_),
    .B2(\cpu.dcache.r_tag[1][6] ),
    .A2(_09266_),
    .A1(\cpu.dcache.r_tag[2][6] ));
 sg13g2_a22oi_1 _16133_ (.Y(_09411_),
    .B1(_09285_),
    .B2(\cpu.dcache.r_tag[6][6] ),
    .A2(_09279_),
    .A1(\cpu.dcache.r_tag[3][6] ));
 sg13g2_mux2_1 _16134_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(\cpu.dcache.r_tag[7][6] ),
    .S(_09088_),
    .X(_09412_));
 sg13g2_a22oi_1 _16135_ (.Y(_09413_),
    .B1(_09412_),
    .B2(net1035),
    .A2(_09289_),
    .A1(\cpu.dcache.r_tag[4][6] ));
 sg13g2_nand2b_1 _16136_ (.Y(_09414_),
    .B(net1024),
    .A_N(_09413_));
 sg13g2_and4_1 _16137_ (.A(_09260_),
    .B(_09410_),
    .C(_09411_),
    .D(_09414_),
    .X(_09415_));
 sg13g2_a21oi_1 _16138_ (.A1(_00232_),
    .A2(net615),
    .Y(_09416_),
    .B1(_09415_));
 sg13g2_xnor2_1 _16139_ (.Y(_09417_),
    .A(_00231_),
    .B(_09416_));
 sg13g2_inv_1 _16140_ (.Y(_09418_),
    .A(_00242_));
 sg13g2_a22oi_1 _16141_ (.Y(_09419_),
    .B1(_09345_),
    .B2(\cpu.dcache.r_tag[5][11] ),
    .A2(_09272_),
    .A1(\cpu.dcache.r_tag[1][11] ));
 sg13g2_a22oi_1 _16142_ (.Y(_09420_),
    .B1(net613),
    .B2(\cpu.dcache.r_tag[3][11] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][11] ));
 sg13g2_mux2_1 _16143_ (.A0(\cpu.dcache.r_tag[4][11] ),
    .A1(\cpu.dcache.r_tag[6][11] ),
    .S(net1034),
    .X(_09421_));
 sg13g2_a22oi_1 _16144_ (.Y(_09422_),
    .B1(_09421_),
    .B2(_09252_),
    .A2(net765),
    .A1(\cpu.dcache.r_tag[7][11] ));
 sg13g2_nand2b_1 _16145_ (.Y(_09423_),
    .B(_09255_),
    .A_N(_09422_));
 sg13g2_nand4_1 _16146_ (.B(_09419_),
    .C(_09420_),
    .A(_09260_),
    .Y(_09424_),
    .D(_09423_));
 sg13g2_o21ai_1 _16147_ (.B1(_09424_),
    .Y(_09425_),
    .A1(_09418_),
    .A2(net549));
 sg13g2_xor2_1 _16148_ (.B(_09425_),
    .A(_00241_),
    .X(_09426_));
 sg13g2_or4_1 _16149_ (.A(_09401_),
    .B(_09409_),
    .C(_09417_),
    .D(_09426_),
    .X(_09427_));
 sg13g2_buf_1 _16150_ (.A(net1026),
    .X(_09428_));
 sg13g2_mux4_1 _16151_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net777),
    .X(_09429_));
 sg13g2_mux4_1 _16152_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net777),
    .X(_09430_));
 sg13g2_mux4_1 _16153_ (.S0(_09230_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net777),
    .X(_09431_));
 sg13g2_mux4_1 _16154_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(_09227_),
    .X(_09432_));
 sg13g2_mux4_1 _16155_ (.S0(_08740_),
    .A0(_09429_),
    .A1(_09430_),
    .A2(_09431_),
    .A3(_09432_),
    .S1(net767),
    .X(_09433_));
 sg13g2_nand2_1 _16156_ (.Y(_09434_),
    .A(_08364_),
    .B(_09433_));
 sg13g2_buf_2 _16157_ (.A(_09224_),
    .X(_09435_));
 sg13g2_buf_2 _16158_ (.A(_09226_),
    .X(_09436_));
 sg13g2_mux4_1 _16159_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net763),
    .X(_09437_));
 sg13g2_mux4_1 _16160_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(net763),
    .X(_09438_));
 sg13g2_mux4_1 _16161_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net777),
    .X(_09439_));
 sg13g2_mux4_1 _16162_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(_09227_),
    .X(_09440_));
 sg13g2_mux4_1 _16163_ (.S0(_08740_),
    .A0(_09437_),
    .A1(_09438_),
    .A2(_09439_),
    .A3(_09440_),
    .S1(net774),
    .X(_09441_));
 sg13g2_o21ai_1 _16164_ (.B1(net1026),
    .Y(_09442_),
    .A1(_08513_),
    .A2(_09441_));
 sg13g2_o21ai_1 _16165_ (.B1(_09442_),
    .Y(_09443_),
    .A1(_09428_),
    .A2(_09434_));
 sg13g2_buf_1 _16166_ (.A(_09443_),
    .X(_09444_));
 sg13g2_a22oi_1 _16167_ (.Y(_09445_),
    .B1(net547),
    .B2(\cpu.dcache.r_tag[1][15] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][15] ));
 sg13g2_a22oi_1 _16168_ (.Y(_09446_),
    .B1(_09394_),
    .B2(\cpu.dcache.r_tag[4][15] ),
    .A2(net613),
    .A1(\cpu.dcache.r_tag[3][15] ));
 sg13g2_mux2_1 _16169_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(\cpu.dcache.r_tag[7][15] ),
    .S(net899),
    .X(_09447_));
 sg13g2_a22oi_1 _16170_ (.Y(_09448_),
    .B1(_09447_),
    .B2(net900),
    .A2(net894),
    .A1(\cpu.dcache.r_tag[6][15] ));
 sg13g2_nand2b_1 _16171_ (.Y(_09449_),
    .B(net893),
    .A_N(_09448_));
 sg13g2_and4_1 _16172_ (.A(net549),
    .B(_09445_),
    .C(_09446_),
    .D(_09449_),
    .X(_09450_));
 sg13g2_a21oi_1 _16173_ (.A1(_00246_),
    .A2(net615),
    .Y(_09451_),
    .B1(_09450_));
 sg13g2_xnor2_1 _16174_ (.Y(_09452_),
    .A(net438),
    .B(_09451_));
 sg13g2_mux4_1 _16175_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net763),
    .X(_09453_));
 sg13g2_mux4_1 _16176_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net763),
    .X(_09454_));
 sg13g2_mux4_1 _16177_ (.S0(_09230_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net763),
    .X(_09455_));
 sg13g2_mux4_1 _16178_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net763),
    .X(_09456_));
 sg13g2_buf_2 _16179_ (.A(net1112),
    .X(_09457_));
 sg13g2_mux4_1 _16180_ (.S0(net767),
    .A0(_09453_),
    .A1(_09454_),
    .A2(_09455_),
    .A3(_09456_),
    .S1(net1023),
    .X(_09458_));
 sg13g2_nand2_1 _16181_ (.Y(_09459_),
    .A(net683),
    .B(_09458_));
 sg13g2_mux4_1 _16182_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(net763),
    .X(_09460_));
 sg13g2_mux4_1 _16183_ (.S0(_09435_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net763),
    .X(_09461_));
 sg13g2_mux4_1 _16184_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(_09436_),
    .X(_09462_));
 sg13g2_mux4_1 _16185_ (.S0(net776),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(_09436_),
    .X(_09463_));
 sg13g2_mux4_1 _16186_ (.S0(net767),
    .A0(_09460_),
    .A1(_09461_),
    .A2(_09462_),
    .A3(_09463_),
    .S1(net1023),
    .X(_09464_));
 sg13g2_nand2_1 _16187_ (.Y(_09465_),
    .A(net674),
    .B(_09464_));
 sg13g2_a21oi_1 _16188_ (.A1(_09459_),
    .A2(_09465_),
    .Y(_09466_),
    .B1(_08435_));
 sg13g2_buf_1 _16189_ (.A(_09466_),
    .X(_09467_));
 sg13g2_a22oi_1 _16190_ (.Y(_09468_),
    .B1(net547),
    .B2(\cpu.dcache.r_tag[1][23] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][23] ));
 sg13g2_a22oi_1 _16191_ (.Y(_09469_),
    .B1(_09285_),
    .B2(\cpu.dcache.r_tag[6][23] ),
    .A2(net613),
    .A1(\cpu.dcache.r_tag[3][23] ));
 sg13g2_mux2_1 _16192_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(\cpu.dcache.r_tag[7][23] ),
    .S(_09089_),
    .X(_09470_));
 sg13g2_a22oi_1 _16193_ (.Y(_09471_),
    .B1(_09470_),
    .B2(net900),
    .A2(_09289_),
    .A1(\cpu.dcache.r_tag[4][23] ));
 sg13g2_nand2b_1 _16194_ (.Y(_09472_),
    .B(_09293_),
    .A_N(_09471_));
 sg13g2_and4_1 _16195_ (.A(net549),
    .B(_09468_),
    .C(_09469_),
    .D(_09472_),
    .X(_09473_));
 sg13g2_a21oi_1 _16196_ (.A1(_00251_),
    .A2(net615),
    .Y(_09474_),
    .B1(_09473_));
 sg13g2_xnor2_1 _16197_ (.Y(_09475_),
    .A(net437),
    .B(_09474_));
 sg13g2_nand2_1 _16198_ (.Y(_09476_),
    .A(_09452_),
    .B(_09475_));
 sg13g2_nor4_1 _16199_ (.A(_09356_),
    .B(_09388_),
    .C(_09427_),
    .D(_09476_),
    .Y(_09477_));
 sg13g2_buf_1 _16200_ (.A(net774),
    .X(_09478_));
 sg13g2_buf_2 _16201_ (.A(_09226_),
    .X(_09479_));
 sg13g2_mux4_1 _16202_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net762),
    .X(_09480_));
 sg13g2_mux4_1 _16203_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net762),
    .X(_09481_));
 sg13g2_mux4_1 _16204_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net762),
    .X(_09482_));
 sg13g2_mux4_1 _16205_ (.S0(_09435_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net762),
    .X(_09483_));
 sg13g2_mux4_1 _16206_ (.S0(_08740_),
    .A0(_09480_),
    .A1(_09481_),
    .A2(_09482_),
    .A3(_09483_),
    .S1(net1023),
    .X(_09484_));
 sg13g2_nand2_1 _16207_ (.Y(_09485_),
    .A(_08364_),
    .B(_09484_));
 sg13g2_mux4_1 _16208_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net762),
    .X(_09486_));
 sg13g2_mux4_1 _16209_ (.S0(_09336_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(_09479_),
    .X(_09487_));
 sg13g2_mux4_1 _16210_ (.S0(net764),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net762),
    .X(_09488_));
 sg13g2_mux4_1 _16211_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(net762),
    .X(_09489_));
 sg13g2_mux4_1 _16212_ (.S0(_08740_),
    .A0(_09486_),
    .A1(_09487_),
    .A2(_09488_),
    .A3(_09489_),
    .S1(net1023),
    .X(_09490_));
 sg13g2_o21ai_1 _16213_ (.B1(net774),
    .Y(_09491_),
    .A1(_08513_),
    .A2(_09490_));
 sg13g2_o21ai_1 _16214_ (.B1(_09491_),
    .Y(_09492_),
    .A1(_09478_),
    .A2(_09485_));
 sg13g2_buf_1 _16215_ (.A(_09492_),
    .X(_09493_));
 sg13g2_a22oi_1 _16216_ (.Y(_09494_),
    .B1(_09345_),
    .B2(\cpu.dcache.r_tag[5][14] ),
    .A2(net547),
    .A1(\cpu.dcache.r_tag[1][14] ));
 sg13g2_a22oi_1 _16217_ (.Y(_09495_),
    .B1(_09281_),
    .B2(\cpu.dcache.r_tag[3][14] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][14] ));
 sg13g2_mux2_1 _16218_ (.A0(\cpu.dcache.r_tag[4][14] ),
    .A1(\cpu.dcache.r_tag[6][14] ),
    .S(net899),
    .X(_09496_));
 sg13g2_a22oi_1 _16219_ (.Y(_09497_),
    .B1(_09496_),
    .B2(net892),
    .A2(net765),
    .A1(\cpu.dcache.r_tag[7][14] ));
 sg13g2_nand2b_1 _16220_ (.Y(_09498_),
    .B(net893),
    .A_N(_09497_));
 sg13g2_and4_1 _16221_ (.A(net549),
    .B(_09494_),
    .C(_09495_),
    .D(_09498_),
    .X(_09499_));
 sg13g2_a21oi_1 _16222_ (.A1(_00245_),
    .A2(_09257_),
    .Y(_09500_),
    .B1(_09499_));
 sg13g2_xor2_1 _16223_ (.B(_09500_),
    .A(net436),
    .X(_09501_));
 sg13g2_mux4_1 _16224_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net768),
    .X(_09502_));
 sg13g2_mux4_1 _16225_ (.S0(net769),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net768),
    .X(_09503_));
 sg13g2_mux4_1 _16226_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net768),
    .X(_09504_));
 sg13g2_mux4_1 _16227_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net768),
    .X(_09505_));
 sg13g2_mux4_1 _16228_ (.S0(_09331_),
    .A0(_09502_),
    .A1(_09503_),
    .A2(_09504_),
    .A3(_09505_),
    .S1(net1023),
    .X(_09506_));
 sg13g2_nand2_1 _16229_ (.Y(_09507_),
    .A(net683),
    .B(_09506_));
 sg13g2_mux4_1 _16230_ (.S0(_09325_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net768),
    .X(_09508_));
 sg13g2_mux4_1 _16231_ (.S0(_09325_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(_09328_),
    .X(_09509_));
 sg13g2_mux4_1 _16232_ (.S0(net766),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(net762),
    .X(_09510_));
 sg13g2_mux4_1 _16233_ (.S0(_09336_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(_09479_),
    .X(_09511_));
 sg13g2_mux4_1 _16234_ (.S0(net767),
    .A0(_09508_),
    .A1(_09509_),
    .A2(_09510_),
    .A3(_09511_),
    .S1(_09457_),
    .X(_09512_));
 sg13g2_nand2_1 _16235_ (.Y(_09513_),
    .A(net674),
    .B(_09512_));
 sg13g2_a21oi_2 _16236_ (.B1(_08435_),
    .Y(_09514_),
    .A2(_09513_),
    .A1(_09507_));
 sg13g2_buf_1 _16237_ (.A(_09514_),
    .X(_09515_));
 sg13g2_a22oi_1 _16238_ (.Y(_09516_),
    .B1(_09274_),
    .B2(\cpu.dcache.r_tag[1][16] ),
    .A2(_09268_),
    .A1(\cpu.dcache.r_tag[2][16] ));
 sg13g2_a22oi_1 _16239_ (.Y(_09517_),
    .B1(net612),
    .B2(\cpu.dcache.r_tag[6][16] ),
    .A2(net613),
    .A1(\cpu.dcache.r_tag[3][16] ));
 sg13g2_mux2_1 _16240_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(\cpu.dcache.r_tag[7][16] ),
    .S(net899),
    .X(_09518_));
 sg13g2_a22oi_1 _16241_ (.Y(_09519_),
    .B1(_09518_),
    .B2(net900),
    .A2(_09290_),
    .A1(\cpu.dcache.r_tag[4][16] ));
 sg13g2_nand2b_1 _16242_ (.Y(_09520_),
    .B(net893),
    .A_N(_09519_));
 sg13g2_and4_1 _16243_ (.A(net549),
    .B(_09516_),
    .C(_09517_),
    .D(_09520_),
    .X(_09521_));
 sg13g2_a21oi_1 _16244_ (.A1(_00247_),
    .A2(net550),
    .Y(_09522_),
    .B1(_09521_));
 sg13g2_xor2_1 _16245_ (.B(_09522_),
    .A(net435),
    .X(_09523_));
 sg13g2_mux4_1 _16246_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net775),
    .X(_09524_));
 sg13g2_mux4_1 _16247_ (.S0(net778),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net775),
    .X(_09525_));
 sg13g2_mux4_1 _16248_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net770),
    .X(_09526_));
 sg13g2_mux4_1 _16249_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net770),
    .X(_09527_));
 sg13g2_mux4_1 _16250_ (.S0(net774),
    .A0(_09524_),
    .A1(_09525_),
    .A2(_09526_),
    .A3(_09527_),
    .S1(net1026),
    .X(_09528_));
 sg13g2_nand2_1 _16251_ (.Y(_09529_),
    .A(net683),
    .B(_09528_));
 sg13g2_mux4_1 _16252_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(net775),
    .X(_09530_));
 sg13g2_mux4_1 _16253_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net775),
    .X(_09531_));
 sg13g2_mux4_1 _16254_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net770),
    .X(_09532_));
 sg13g2_mux4_1 _16255_ (.S0(net771),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net770),
    .X(_09533_));
 sg13g2_mux4_1 _16256_ (.S0(net774),
    .A0(_09530_),
    .A1(_09531_),
    .A2(_09532_),
    .A3(_09533_),
    .S1(net1026),
    .X(_09534_));
 sg13g2_nand2_1 _16257_ (.Y(_09535_),
    .A(net674),
    .B(_09534_));
 sg13g2_a21oi_2 _16258_ (.B1(_08436_),
    .Y(_09536_),
    .A2(_09535_),
    .A1(_09529_));
 sg13g2_buf_1 _16259_ (.A(_09536_),
    .X(_09537_));
 sg13g2_a22oi_1 _16260_ (.Y(_09538_),
    .B1(_09281_),
    .B2(\cpu.dcache.r_tag[3][21] ),
    .A2(_09268_),
    .A1(\cpu.dcache.r_tag[2][21] ));
 sg13g2_a22oi_1 _16261_ (.Y(_09539_),
    .B1(net545),
    .B2(\cpu.dcache.r_tag[5][21] ),
    .A2(_09274_),
    .A1(\cpu.dcache.r_tag[1][21] ));
 sg13g2_mux2_1 _16262_ (.A0(\cpu.dcache.r_tag[4][21] ),
    .A1(\cpu.dcache.r_tag[6][21] ),
    .S(net783),
    .X(_09540_));
 sg13g2_a22oi_1 _16263_ (.Y(_09541_),
    .B1(_09540_),
    .B2(_09351_),
    .A2(net765),
    .A1(\cpu.dcache.r_tag[7][21] ));
 sg13g2_nand2b_1 _16264_ (.Y(_09542_),
    .B(_09294_),
    .A_N(_09541_));
 sg13g2_nand4_1 _16265_ (.B(_09538_),
    .C(_09539_),
    .A(_09262_),
    .Y(_09543_),
    .D(_09542_));
 sg13g2_o21ai_1 _16266_ (.B1(_09543_),
    .Y(_09544_),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .A2(net494));
 sg13g2_xnor2_1 _16267_ (.Y(_09545_),
    .A(_09537_),
    .B(_09544_));
 sg13g2_buf_2 _16268_ (.A(_08754_),
    .X(_09546_));
 sg13g2_mux4_1 _16269_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net777),
    .X(_09547_));
 sg13g2_mux4_1 _16270_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net777),
    .X(_09548_));
 sg13g2_buf_1 _16271_ (.A(_09226_),
    .X(_09549_));
 sg13g2_mux4_1 _16272_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net761),
    .X(_09550_));
 sg13g2_mux4_1 _16273_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(net761),
    .X(_09551_));
 sg13g2_mux4_1 _16274_ (.S0(_09331_),
    .A0(_09547_),
    .A1(_09548_),
    .A2(_09550_),
    .A3(_09551_),
    .S1(net1023),
    .X(_09552_));
 sg13g2_nand2_1 _16275_ (.Y(_09553_),
    .A(_08832_),
    .B(_09552_));
 sg13g2_mux4_1 _16276_ (.S0(_09546_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(net761),
    .X(_09554_));
 sg13g2_mux4_1 _16277_ (.S0(_09546_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net777),
    .X(_09555_));
 sg13g2_buf_2 _16278_ (.A(_08754_),
    .X(_09556_));
 sg13g2_mux4_1 _16279_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(_09549_),
    .X(_09557_));
 sg13g2_mux4_1 _16280_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(_09549_),
    .X(_09558_));
 sg13g2_mux4_1 _16281_ (.S0(net767),
    .A0(_09554_),
    .A1(_09555_),
    .A2(_09557_),
    .A3(_09558_),
    .S1(net1023),
    .X(_09559_));
 sg13g2_nand2_1 _16282_ (.Y(_09560_),
    .A(_09245_),
    .B(_09559_));
 sg13g2_a21oi_1 _16283_ (.A1(_09553_),
    .A2(_09560_),
    .Y(_09561_),
    .B1(_08435_));
 sg13g2_buf_1 _16284_ (.A(_09561_),
    .X(_09562_));
 sg13g2_inv_1 _16285_ (.Y(_09563_),
    .A(_00250_));
 sg13g2_a22oi_1 _16286_ (.Y(_09564_),
    .B1(_09345_),
    .B2(\cpu.dcache.r_tag[5][19] ),
    .A2(net547),
    .A1(\cpu.dcache.r_tag[1][19] ));
 sg13g2_a22oi_1 _16287_ (.Y(_09565_),
    .B1(net613),
    .B2(\cpu.dcache.r_tag[3][19] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][19] ));
 sg13g2_mux2_1 _16288_ (.A0(\cpu.dcache.r_tag[4][19] ),
    .A1(\cpu.dcache.r_tag[6][19] ),
    .S(net899),
    .X(_09566_));
 sg13g2_a22oi_1 _16289_ (.Y(_09567_),
    .B1(_09566_),
    .B2(_09252_),
    .A2(_09349_),
    .A1(\cpu.dcache.r_tag[7][19] ));
 sg13g2_nand2b_1 _16290_ (.Y(_09568_),
    .B(net893),
    .A_N(_09567_));
 sg13g2_nand4_1 _16291_ (.B(_09564_),
    .C(_09565_),
    .A(net549),
    .Y(_09569_),
    .D(_09568_));
 sg13g2_o21ai_1 _16292_ (.B1(_09569_),
    .Y(_09570_),
    .A1(_09563_),
    .A2(net494));
 sg13g2_xor2_1 _16293_ (.B(_09570_),
    .A(net433),
    .X(_09571_));
 sg13g2_mux4_1 _16294_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net761),
    .X(_09572_));
 sg13g2_mux4_1 _16295_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net761),
    .X(_09573_));
 sg13g2_buf_1 _16296_ (.A(_09226_),
    .X(_09574_));
 sg13g2_mux4_1 _16297_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net760),
    .X(_09575_));
 sg13g2_mux4_1 _16298_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net760),
    .X(_09576_));
 sg13g2_mux4_1 _16299_ (.S0(net767),
    .A0(_09572_),
    .A1(_09573_),
    .A2(_09575_),
    .A3(_09576_),
    .S1(net1023),
    .X(_09577_));
 sg13g2_nand2_1 _16300_ (.Y(_09578_),
    .A(net683),
    .B(_09577_));
 sg13g2_mux4_1 _16301_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(net761),
    .X(_09579_));
 sg13g2_mux4_1 _16302_ (.S0(net889),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(net761),
    .X(_09580_));
 sg13g2_mux4_1 _16303_ (.S0(_09556_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(_09574_),
    .X(_09581_));
 sg13g2_mux4_1 _16304_ (.S0(_09556_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(_09574_),
    .X(_09582_));
 sg13g2_mux4_1 _16305_ (.S0(net902),
    .A0(_09579_),
    .A1(_09580_),
    .A2(_09581_),
    .A3(_09582_),
    .S1(net1112),
    .X(_09583_));
 sg13g2_nand2_1 _16306_ (.Y(_09584_),
    .A(_09245_),
    .B(_09583_));
 sg13g2_a21oi_1 _16307_ (.A1(_09578_),
    .A2(_09584_),
    .Y(_09585_),
    .B1(_08435_));
 sg13g2_buf_1 _16308_ (.A(_09585_),
    .X(_09586_));
 sg13g2_a22oi_1 _16309_ (.Y(_09587_),
    .B1(net547),
    .B2(\cpu.dcache.r_tag[1][17] ),
    .A2(_09267_),
    .A1(\cpu.dcache.r_tag[2][17] ));
 sg13g2_a22oi_1 _16310_ (.Y(_09588_),
    .B1(_09285_),
    .B2(\cpu.dcache.r_tag[6][17] ),
    .A2(_09280_),
    .A1(\cpu.dcache.r_tag[3][17] ));
 sg13g2_mux2_1 _16311_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(\cpu.dcache.r_tag[7][17] ),
    .S(net899),
    .X(_09589_));
 sg13g2_a22oi_1 _16312_ (.Y(_09590_),
    .B1(_09589_),
    .B2(net1035),
    .A2(_09289_),
    .A1(\cpu.dcache.r_tag[4][17] ));
 sg13g2_nand2b_1 _16313_ (.Y(_09591_),
    .B(_09293_),
    .A_N(_09590_));
 sg13g2_and4_1 _16314_ (.A(_09261_),
    .B(_09587_),
    .C(_09588_),
    .D(_09591_),
    .X(_09592_));
 sg13g2_a21oi_1 _16315_ (.A1(_00248_),
    .A2(_09257_),
    .Y(_09593_),
    .B1(_09592_));
 sg13g2_xnor2_1 _16316_ (.Y(_09594_),
    .A(net432),
    .B(_09593_));
 sg13g2_mux4_1 _16317_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net760),
    .X(_09595_));
 sg13g2_mux4_1 _16318_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net761),
    .X(_09596_));
 sg13g2_buf_2 _16319_ (.A(_08754_),
    .X(_09597_));
 sg13g2_mux4_1 _16320_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net895),
    .X(_09598_));
 sg13g2_mux4_1 _16321_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net895),
    .X(_09599_));
 sg13g2_mux4_1 _16322_ (.S0(net902),
    .A0(_09595_),
    .A1(_09596_),
    .A2(_09598_),
    .A3(_09599_),
    .S1(net1112),
    .X(_09600_));
 sg13g2_nand2_1 _16323_ (.Y(_09601_),
    .A(net683),
    .B(_09600_));
 sg13g2_mux4_1 _16324_ (.S0(_09597_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net760),
    .X(_09602_));
 sg13g2_mux4_1 _16325_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net760),
    .X(_09603_));
 sg13g2_mux4_1 _16326_ (.S0(_09597_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(_09233_),
    .X(_09604_));
 sg13g2_mux4_1 _16327_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(_09233_),
    .X(_09605_));
 sg13g2_mux4_1 _16328_ (.S0(net902),
    .A0(_09602_),
    .A1(_09603_),
    .A2(_09604_),
    .A3(_09605_),
    .S1(net1112),
    .X(_09606_));
 sg13g2_nand2_1 _16329_ (.Y(_09607_),
    .A(net674),
    .B(_09606_));
 sg13g2_a21oi_2 _16330_ (.B1(_08435_),
    .Y(_09608_),
    .A2(_09607_),
    .A1(_09601_));
 sg13g2_buf_1 _16331_ (.A(_09608_),
    .X(_09609_));
 sg13g2_a22oi_1 _16332_ (.Y(_09610_),
    .B1(net613),
    .B2(\cpu.dcache.r_tag[3][22] ),
    .A2(net614),
    .A1(\cpu.dcache.r_tag[2][22] ));
 sg13g2_a22oi_1 _16333_ (.Y(_09611_),
    .B1(_09345_),
    .B2(\cpu.dcache.r_tag[5][22] ),
    .A2(_09273_),
    .A1(\cpu.dcache.r_tag[1][22] ));
 sg13g2_mux2_1 _16334_ (.A0(\cpu.dcache.r_tag[4][22] ),
    .A1(\cpu.dcache.r_tag[6][22] ),
    .S(net899),
    .X(_09612_));
 sg13g2_a22oi_1 _16335_ (.Y(_09613_),
    .B1(_09612_),
    .B2(_09252_),
    .A2(_09349_),
    .A1(\cpu.dcache.r_tag[7][22] ));
 sg13g2_nand2b_1 _16336_ (.Y(_09614_),
    .B(net893),
    .A_N(_09613_));
 sg13g2_nand4_1 _16337_ (.B(_09610_),
    .C(_09611_),
    .A(_09261_),
    .Y(_09615_),
    .D(_09614_));
 sg13g2_o21ai_1 _16338_ (.B1(_09615_),
    .Y(_09616_),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .A2(net494));
 sg13g2_xor2_1 _16339_ (.B(_09616_),
    .A(net431),
    .X(_09617_));
 sg13g2_mux4_1 _16340_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net760),
    .X(_09618_));
 sg13g2_mux4_1 _16341_ (.S0(net888),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net760),
    .X(_09619_));
 sg13g2_mux4_1 _16342_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net895),
    .X(_09620_));
 sg13g2_mux4_1 _16343_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net895),
    .X(_09621_));
 sg13g2_mux4_1 _16344_ (.S0(_08744_),
    .A0(_09618_),
    .A1(_09619_),
    .A2(_09620_),
    .A3(_09621_),
    .S1(_08749_),
    .X(_09622_));
 sg13g2_nand2_1 _16345_ (.Y(_09623_),
    .A(net683),
    .B(_09622_));
 sg13g2_mux4_1 _16346_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net895),
    .X(_09624_));
 sg13g2_mux4_1 _16347_ (.S0(net887),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net760),
    .X(_09625_));
 sg13g2_mux4_1 _16348_ (.S0(_09224_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net895),
    .X(_09626_));
 sg13g2_mux4_1 _16349_ (.S0(_09224_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net895),
    .X(_09627_));
 sg13g2_mux4_1 _16350_ (.S0(_08744_),
    .A0(_09624_),
    .A1(_09625_),
    .A2(_09626_),
    .A3(_09627_),
    .S1(_08749_),
    .X(_09628_));
 sg13g2_nand2_1 _16351_ (.Y(_09629_),
    .A(_08740_),
    .B(_09628_));
 sg13g2_a21oi_2 _16352_ (.B1(_08435_),
    .Y(_09630_),
    .A2(_09629_),
    .A1(_09623_));
 sg13g2_buf_1 _16353_ (.A(_09630_),
    .X(_09631_));
 sg13g2_a22oi_1 _16354_ (.Y(_09632_),
    .B1(_09273_),
    .B2(\cpu.dcache.r_tag[1][20] ),
    .A2(_09267_),
    .A1(\cpu.dcache.r_tag[2][20] ));
 sg13g2_a22oi_1 _16355_ (.Y(_09633_),
    .B1(_09285_),
    .B2(\cpu.dcache.r_tag[6][20] ),
    .A2(_09280_),
    .A1(\cpu.dcache.r_tag[3][20] ));
 sg13g2_mux2_1 _16356_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(\cpu.dcache.r_tag[7][20] ),
    .S(net899),
    .X(_09634_));
 sg13g2_a22oi_1 _16357_ (.Y(_09635_),
    .B1(_09634_),
    .B2(_09083_),
    .A2(_09290_),
    .A1(\cpu.dcache.r_tag[4][20] ));
 sg13g2_nand2b_1 _16358_ (.Y(_09636_),
    .B(net893),
    .A_N(_09635_));
 sg13g2_nand4_1 _16359_ (.B(_09632_),
    .C(_09633_),
    .A(net549),
    .Y(_09637_),
    .D(_09636_));
 sg13g2_o21ai_1 _16360_ (.B1(_09637_),
    .Y(_09638_),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .A2(net494));
 sg13g2_xor2_1 _16361_ (.B(_09638_),
    .A(net430),
    .X(_09639_));
 sg13g2_nand4_1 _16362_ (.B(_09594_),
    .C(_09617_),
    .A(_09571_),
    .Y(_09640_),
    .D(_09639_));
 sg13g2_nor4_1 _16363_ (.A(_09501_),
    .B(_09523_),
    .C(_09545_),
    .D(_09640_),
    .Y(_09641_));
 sg13g2_nand4_1 _16364_ (.B(_09324_),
    .C(_09477_),
    .A(_09298_),
    .Y(_09642_),
    .D(_09641_));
 sg13g2_mux4_1 _16365_ (.S0(net784),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(_09091_),
    .X(_09643_));
 sg13g2_mux4_1 _16366_ (.S0(net784),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net783),
    .X(_09644_));
 sg13g2_mux2_1 _16367_ (.A0(_09643_),
    .A1(_09644_),
    .S(net891),
    .X(_09645_));
 sg13g2_mux4_1 _16368_ (.S0(_09084_),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(net681),
    .X(_09646_));
 sg13g2_mux4_1 _16369_ (.S0(net784),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(net681),
    .X(_09647_));
 sg13g2_mux2_1 _16370_ (.A0(_09646_),
    .A1(_09647_),
    .S(net891),
    .X(_09648_));
 sg13g2_and3_1 _16371_ (.X(_09649_),
    .A(_09078_),
    .B(_09645_),
    .C(_09648_));
 sg13g2_buf_1 _16372_ (.A(_09649_),
    .X(_09650_));
 sg13g2_o21ai_1 _16373_ (.B1(_09650_),
    .Y(_09651_),
    .A1(_09223_),
    .A2(_09642_));
 sg13g2_nor2b_1 _16374_ (.A(_09642_),
    .B_N(_09645_),
    .Y(_09652_));
 sg13g2_buf_1 _16375_ (.A(_09652_),
    .X(_09653_));
 sg13g2_or3_1 _16376_ (.A(_09223_),
    .B(_09650_),
    .C(_09653_),
    .X(_09654_));
 sg13g2_buf_1 _16377_ (.A(_09654_),
    .X(_09655_));
 sg13g2_inv_1 _16378_ (.Y(_09656_),
    .A(_09107_));
 sg13g2_nand2_1 _16379_ (.Y(_09657_),
    .A(net886),
    .B(_09078_));
 sg13g2_a221oi_1 _16380_ (.B2(_09655_),
    .C1(_09657_),
    .B1(_09651_),
    .A1(_08764_),
    .Y(_09658_),
    .A2(_09103_));
 sg13g2_a21o_1 _16381_ (.A2(_08732_),
    .A1(_08734_),
    .B1(_09658_),
    .X(_09659_));
 sg13g2_inv_1 _16382_ (.Y(_09660_),
    .A(_09659_));
 sg13g2_nand2_1 _16383_ (.Y(_09661_),
    .A(\cpu.qspi.r_state[17] ),
    .B(_09660_));
 sg13g2_buf_1 _16384_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09662_));
 sg13g2_buf_1 _16385_ (.A(\cpu.qspi.r_ind ),
    .X(_09663_));
 sg13g2_buf_1 _16386_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09664_));
 sg13g2_buf_2 _16387_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09665_));
 sg13g2_buf_1 _16388_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09666_));
 sg13g2_nor3_1 _16389_ (.A(_09664_),
    .B(_09665_),
    .C(_09666_),
    .Y(_09667_));
 sg13g2_nor2b_1 _16390_ (.A(\cpu.qspi.r_count[3] ),
    .B_N(_09667_),
    .Y(_09668_));
 sg13g2_and2_1 _16391_ (.A(_00252_),
    .B(_09668_),
    .X(_09669_));
 sg13g2_buf_1 _16392_ (.A(_09669_),
    .X(_09670_));
 sg13g2_buf_1 _16393_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09671_));
 sg13g2_a221oi_1 _16394_ (.B2(_09671_),
    .C1(\cpu.qspi.r_state[1] ),
    .B1(_09670_),
    .A1(_09662_),
    .Y(_09672_),
    .A2(_09663_));
 sg13g2_a21oi_1 _16395_ (.A1(_09661_),
    .A2(_09672_),
    .Y(_00026_),
    .B1(net618));
 sg13g2_buf_2 _16396_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09673_));
 sg13g2_nand2_1 _16397_ (.Y(_09674_),
    .A(_00252_),
    .B(_09668_));
 sg13g2_buf_1 _16398_ (.A(_09674_),
    .X(_09675_));
 sg13g2_nand2_1 _16399_ (.Y(_09676_),
    .A(_09673_),
    .B(_09675_));
 sg13g2_buf_1 _16400_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09677_));
 sg13g2_nand2b_1 _16401_ (.Y(_09678_),
    .B(_08830_),
    .A_N(_09651_));
 sg13g2_buf_1 _16402_ (.A(_09678_),
    .X(_09679_));
 sg13g2_inv_1 _16403_ (.Y(_09680_),
    .A(net107));
 sg13g2_nand2_1 _16404_ (.Y(_09681_),
    .A(_09677_),
    .B(_09680_));
 sg13g2_a21oi_1 _16405_ (.A1(_09676_),
    .A2(_09681_),
    .Y(_00025_),
    .B1(_09184_));
 sg13g2_buf_1 _16406_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09682_));
 sg13g2_buf_1 _16407_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09683_));
 sg13g2_a21oi_1 _16408_ (.A1(_09682_),
    .A2(_09670_),
    .Y(_09684_),
    .B1(_09683_));
 sg13g2_nor2_1 _16409_ (.A(net617),
    .B(_09684_),
    .Y(_00022_));
 sg13g2_buf_1 _16410_ (.A(_00277_),
    .X(_09685_));
 sg13g2_buf_1 _16411_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09686_));
 sg13g2_nand2_1 _16412_ (.Y(_09687_),
    .A(net1102),
    .B(net671));
 sg13g2_a21oi_1 _16413_ (.A1(_09685_),
    .A2(_09687_),
    .Y(_00023_),
    .B1(_09184_));
 sg13g2_inv_1 _16414_ (.Y(_09688_),
    .A(\cpu.qspi.r_quad[0] ));
 sg13g2_buf_1 _16415_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09689_));
 sg13g2_buf_1 _16416_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09690_));
 sg13g2_nor2_1 _16417_ (.A(_08830_),
    .B(_08449_),
    .Y(_09691_));
 sg13g2_a21oi_1 _16418_ (.A1(_08830_),
    .A2(net437),
    .Y(_09692_),
    .B1(_09691_));
 sg13g2_nor3_1 _16419_ (.A(_09689_),
    .B(_09690_),
    .C(_09692_),
    .Y(_09693_));
 sg13g2_buf_1 _16420_ (.A(_09693_),
    .X(_09694_));
 sg13g2_nor2_1 _16421_ (.A(_09689_),
    .B(_09692_),
    .Y(_09695_));
 sg13g2_a21oi_1 _16422_ (.A1(_09689_),
    .A2(net107),
    .Y(_09696_),
    .B1(_09695_));
 sg13g2_nor2b_1 _16423_ (.A(_09696_),
    .B_N(_09690_),
    .Y(_09697_));
 sg13g2_buf_1 _16424_ (.A(_09697_),
    .X(_09698_));
 sg13g2_or2_1 _16425_ (.X(_09699_),
    .B(net69),
    .A(net324));
 sg13g2_buf_2 _16426_ (.A(_09699_),
    .X(_09700_));
 sg13g2_a22oi_1 _16427_ (.Y(_09701_),
    .B1(net69),
    .B2(\cpu.qspi.r_quad[1] ),
    .A2(net324),
    .A1(\cpu.qspi.r_quad[2] ));
 sg13g2_o21ai_1 _16428_ (.B1(_09701_),
    .Y(_09702_),
    .A1(_09688_),
    .A2(_09700_));
 sg13g2_buf_2 _16429_ (.A(_09702_),
    .X(_09703_));
 sg13g2_inv_1 _16430_ (.Y(_09704_),
    .A(_09703_));
 sg13g2_and2_1 _16431_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09659_),
    .X(_09705_));
 sg13g2_a22oi_1 _16432_ (.Y(_09706_),
    .B1(_09704_),
    .B2(_09705_),
    .A2(net671),
    .A1(_09682_));
 sg13g2_nor2_1 _16433_ (.A(net617),
    .B(_09706_),
    .Y(_00028_));
 sg13g2_nand2_1 _16434_ (.Y(_09707_),
    .A(_09671_),
    .B(_09675_));
 sg13g2_buf_1 _16435_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09708_));
 sg13g2_nand2_1 _16436_ (.Y(_09709_),
    .A(net1101),
    .B(_09670_));
 sg13g2_buf_1 _16437_ (.A(_09183_),
    .X(_09710_));
 sg13g2_a21oi_1 _16438_ (.A1(_09707_),
    .A2(_09709_),
    .Y(_00027_),
    .B1(_09710_));
 sg13g2_inv_1 _16439_ (.Y(_09711_),
    .A(_09663_));
 sg13g2_a21o_1 _16440_ (.A2(_09711_),
    .A1(_09662_),
    .B1(net679),
    .X(_00021_));
 sg13g2_nor2_1 _16441_ (.A(_08334_),
    .B(net191),
    .Y(_09712_));
 sg13g2_nand2_1 _16442_ (.Y(_09713_),
    .A(_08989_),
    .B(_09712_));
 sg13g2_buf_1 _16443_ (.A(\cpu.dec.r_op[10] ),
    .X(_09714_));
 sg13g2_nand2_1 _16444_ (.Y(_09715_),
    .A(_09714_),
    .B(net108));
 sg13g2_o21ai_1 _16445_ (.B1(_09715_),
    .Y(_00011_),
    .A1(net92),
    .A2(_09713_));
 sg13g2_buf_2 _16446_ (.A(\cpu.dec.r_op[1] ),
    .X(_09716_));
 sg13g2_a21oi_1 _16447_ (.A1(_08143_),
    .A2(_08204_),
    .Y(_09717_),
    .B1(_08221_));
 sg13g2_buf_1 _16448_ (.A(_09717_),
    .X(_09718_));
 sg13g2_nor2_1 _16449_ (.A(_09718_),
    .B(_08248_),
    .Y(_09719_));
 sg13g2_buf_1 _16450_ (.A(_09719_),
    .X(_09720_));
 sg13g2_nor2b_1 _16451_ (.A(net190),
    .B_N(_08990_),
    .Y(_09721_));
 sg13g2_and2_1 _16452_ (.A(_08880_),
    .B(_09721_),
    .X(_09722_));
 sg13g2_inv_1 _16453_ (.Y(_09723_),
    .A(net346));
 sg13g2_buf_1 _16454_ (.A(_08986_),
    .X(_09724_));
 sg13g2_nand3_1 _16455_ (.B(_09723_),
    .C(net343),
    .A(_09720_),
    .Y(_09725_));
 sg13g2_nor2_1 _16456_ (.A(_08949_),
    .B(_09725_),
    .Y(_09726_));
 sg13g2_a21oi_1 _16457_ (.A1(_09720_),
    .A2(_09722_),
    .Y(_09727_),
    .B1(_09726_));
 sg13g2_nor3_1 _16458_ (.A(net109),
    .B(_08889_),
    .C(_09727_),
    .Y(_09728_));
 sg13g2_a21o_1 _16459_ (.A2(net110),
    .A1(_09716_),
    .B1(_09728_),
    .X(_00012_));
 sg13g2_buf_1 _16460_ (.A(_08223_),
    .X(_09729_));
 sg13g2_buf_1 _16461_ (.A(_08886_),
    .X(_09730_));
 sg13g2_buf_1 _16462_ (.A(_08334_),
    .X(_09731_));
 sg13g2_nand3_1 _16463_ (.B(net189),
    .C(_09722_),
    .A(net166),
    .Y(_09732_));
 sg13g2_o21ai_1 _16464_ (.B1(_09732_),
    .Y(_09733_),
    .A1(net166),
    .A2(net189));
 sg13g2_nand4_1 _16465_ (.B(net147),
    .C(net191),
    .A(_09729_),
    .Y(_09734_),
    .D(_09733_));
 sg13g2_buf_1 _16466_ (.A(\cpu.dec.r_op[9] ),
    .X(_09735_));
 sg13g2_buf_1 _16467_ (.A(_09735_),
    .X(_09736_));
 sg13g2_nand2_1 _16468_ (.Y(_09737_),
    .A(_09736_),
    .B(net108));
 sg13g2_o21ai_1 _16469_ (.B1(_09737_),
    .Y(_00020_),
    .A1(net92),
    .A2(_09734_));
 sg13g2_buf_2 _16470_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09738_));
 sg13g2_a21oi_1 _16471_ (.A1(_09708_),
    .A2(net671),
    .Y(_09739_),
    .B1(_09738_));
 sg13g2_nor2_1 _16472_ (.A(net617),
    .B(_09739_),
    .Y(_00024_));
 sg13g2_nor2_1 _16473_ (.A(_08271_),
    .B(_08884_),
    .Y(_09740_));
 sg13g2_buf_1 _16474_ (.A(_09740_),
    .X(_09741_));
 sg13g2_nor2_1 _16475_ (.A(_08223_),
    .B(_08248_),
    .Y(_09742_));
 sg13g2_nand2_1 _16476_ (.Y(_09743_),
    .A(_09741_),
    .B(_09742_));
 sg13g2_buf_1 _16477_ (.A(\cpu.dec.r_op[8] ),
    .X(_09744_));
 sg13g2_nand2_1 _16478_ (.Y(_09745_),
    .A(_09744_),
    .B(_08997_));
 sg13g2_o21ai_1 _16479_ (.B1(_09745_),
    .Y(_00019_),
    .A1(_08928_),
    .A2(_09743_));
 sg13g2_a21oi_1 _16480_ (.A1(_08919_),
    .A2(_09721_),
    .Y(_09746_),
    .B1(_08335_));
 sg13g2_nor4_1 _16481_ (.A(_08251_),
    .B(_08311_),
    .C(_08887_),
    .D(_09746_),
    .Y(_09747_));
 sg13g2_buf_1 _16482_ (.A(\cpu.dec.r_op[2] ),
    .X(_09748_));
 sg13g2_buf_1 _16483_ (.A(net1099),
    .X(_09749_));
 sg13g2_nand3_1 _16484_ (.B(_08668_),
    .C(_08718_),
    .A(_08709_),
    .Y(_09750_));
 sg13g2_nand4_1 _16485_ (.B(_08688_),
    .C(_08691_),
    .A(_08678_),
    .Y(_09751_),
    .D(_08728_));
 sg13g2_nor2_1 _16486_ (.A(_09750_),
    .B(_09751_),
    .Y(_09752_));
 sg13g2_nand4_1 _16487_ (.B(_08485_),
    .C(_08551_),
    .A(_08458_),
    .Y(_09753_),
    .D(_09752_));
 sg13g2_nor3_1 _16488_ (.A(_08409_),
    .B(_08434_),
    .C(_09753_),
    .Y(_09754_));
 sg13g2_inv_1 _16489_ (.Y(_09755_),
    .A(_08506_));
 sg13g2_inv_1 _16490_ (.Y(_09756_),
    .A(_08572_));
 sg13g2_nor4_1 _16491_ (.A(_09755_),
    .B(_08592_),
    .C(_08657_),
    .D(_09756_),
    .Y(_09757_));
 sg13g2_nor2_1 _16492_ (.A(_08615_),
    .B(_08636_),
    .Y(_09758_));
 sg13g2_nand4_1 _16493_ (.B(_09757_),
    .C(_08529_),
    .A(_09754_),
    .Y(_09759_),
    .D(_09758_));
 sg13g2_nand3b_1 _16494_ (.B(_08733_),
    .C(_08837_),
    .Y(_09760_),
    .A_N(_09759_));
 sg13g2_buf_2 _16495_ (.A(_09760_),
    .X(_09761_));
 sg13g2_buf_1 _16496_ (.A(_09761_),
    .X(_09762_));
 sg13g2_mux2_1 _16497_ (.A0(_09747_),
    .A1(net1021),
    .S(net91),
    .X(_00013_));
 sg13g2_nand2b_1 _16498_ (.Y(_09763_),
    .B(_08969_),
    .A_N(_08986_));
 sg13g2_nand2_1 _16499_ (.Y(_09764_),
    .A(_08919_),
    .B(_09721_));
 sg13g2_o21ai_1 _16500_ (.B1(_09764_),
    .Y(_09765_),
    .A1(_08949_),
    .A2(_09763_));
 sg13g2_and2_1 _16501_ (.A(_08925_),
    .B(_09765_),
    .X(_09766_));
 sg13g2_buf_1 _16502_ (.A(\cpu.dec.r_op[7] ),
    .X(_09767_));
 sg13g2_buf_1 _16503_ (.A(_08840_),
    .X(_09768_));
 sg13g2_mux2_1 _16504_ (.A0(_09766_),
    .A1(_09767_),
    .S(net106),
    .X(_00018_));
 sg13g2_buf_1 _16505_ (.A(\cpu.uart.r_div[11] ),
    .X(_09769_));
 sg13g2_nor3_2 _16506_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09770_));
 sg13g2_nor2b_1 _16507_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09770_),
    .Y(_09771_));
 sg13g2_nor2b_1 _16508_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09771_),
    .Y(_09772_));
 sg13g2_nor2b_1 _16509_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09772_),
    .Y(_09773_));
 sg13g2_nor2b_1 _16510_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09773_),
    .Y(_09774_));
 sg13g2_nand2b_1 _16511_ (.Y(_09775_),
    .B(_09774_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16512_ (.A(\cpu.uart.r_div[8] ),
    .B(_09775_),
    .Y(_09776_));
 sg13g2_nand2b_1 _16513_ (.Y(_09777_),
    .B(_09776_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16514_ (.A(_09777_),
    .X(_09778_));
 sg13g2_nor3_1 _16515_ (.A(_09769_),
    .B(\cpu.uart.r_div[10] ),
    .C(_09778_),
    .Y(_09779_));
 sg13g2_buf_1 _16516_ (.A(_09779_),
    .X(_09780_));
 sg13g2_nor2_1 _16517_ (.A(net896),
    .B(net342),
    .Y(_09781_));
 sg13g2_buf_1 _16518_ (.A(_09781_),
    .X(_09782_));
 sg13g2_buf_1 _16519_ (.A(net248),
    .X(_09783_));
 sg13g2_mux2_1 _16520_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00279_),
    .S(net213),
    .X(_00079_));
 sg13g2_xnor2_1 _16521_ (.Y(_09784_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16522_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09784_),
    .S(_09783_),
    .X(_00082_));
 sg13g2_o21ai_1 _16523_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09785_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16524_ (.A(_09770_),
    .B_N(_09785_),
    .Y(_09786_));
 sg13g2_nor2_1 _16525_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net248),
    .Y(_09787_));
 sg13g2_a21oi_1 _16526_ (.A1(_09783_),
    .A2(_09786_),
    .Y(_00083_),
    .B1(_09787_));
 sg13g2_xnor2_1 _16527_ (.Y(_09788_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09770_));
 sg13g2_nor2_1 _16528_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net248),
    .Y(_09789_));
 sg13g2_a21oi_1 _16529_ (.A1(net213),
    .A2(_09788_),
    .Y(_00084_),
    .B1(_09789_));
 sg13g2_xnor2_1 _16530_ (.Y(_09790_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09771_));
 sg13g2_nor2_1 _16531_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net248),
    .Y(_09791_));
 sg13g2_a21oi_1 _16532_ (.A1(net213),
    .A2(_09790_),
    .Y(_00085_),
    .B1(_09791_));
 sg13g2_xnor2_1 _16533_ (.Y(_09792_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09772_));
 sg13g2_nor2_1 _16534_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net248),
    .Y(_09793_));
 sg13g2_a21oi_1 _16535_ (.A1(net213),
    .A2(_09792_),
    .Y(_00086_),
    .B1(_09793_));
 sg13g2_xnor2_1 _16536_ (.Y(_09794_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09773_));
 sg13g2_nor2_1 _16537_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net248),
    .Y(_09795_));
 sg13g2_a21oi_1 _16538_ (.A1(net213),
    .A2(_09794_),
    .Y(_00087_),
    .B1(_09795_));
 sg13g2_xnor2_1 _16539_ (.Y(_09796_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09774_));
 sg13g2_nor2_1 _16540_ (.A(\cpu.uart.r_div_value[7] ),
    .B(_09782_),
    .Y(_09797_));
 sg13g2_a21oi_1 _16541_ (.A1(net213),
    .A2(_09796_),
    .Y(_00088_),
    .B1(_09797_));
 sg13g2_xor2_1 _16542_ (.B(_09775_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09798_));
 sg13g2_nor2_1 _16543_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net248),
    .Y(_09799_));
 sg13g2_a21oi_1 _16544_ (.A1(net213),
    .A2(_09798_),
    .Y(_00089_),
    .B1(_09799_));
 sg13g2_xnor2_1 _16545_ (.Y(_09800_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09776_));
 sg13g2_nor2_1 _16546_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net248),
    .Y(_09801_));
 sg13g2_a21oi_1 _16547_ (.A1(net213),
    .A2(_09800_),
    .Y(_00090_),
    .B1(_09801_));
 sg13g2_buf_1 _16548_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09802_));
 sg13g2_inv_1 _16549_ (.Y(_09803_),
    .A(_09802_));
 sg13g2_nand2_1 _16550_ (.Y(_09804_),
    .A(net781),
    .B(_09778_));
 sg13g2_o21ai_1 _16551_ (.B1(_09804_),
    .Y(_09805_),
    .A1(_09769_),
    .A2(_09802_));
 sg13g2_inv_1 _16552_ (.Y(_09806_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16553_ (.A(_09806_),
    .B(net779),
    .C(_09778_),
    .Y(_09807_));
 sg13g2_a221oi_1 _16554_ (.B2(_09806_),
    .C1(_09807_),
    .B1(_09805_),
    .A1(_09803_),
    .Y(_00080_),
    .A2(net679));
 sg13g2_nor2_1 _16555_ (.A(\cpu.uart.r_div[10] ),
    .B(_09778_),
    .Y(_09808_));
 sg13g2_nand2_1 _16556_ (.Y(_09809_),
    .A(_09769_),
    .B(net781));
 sg13g2_o21ai_1 _16557_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09810_),
    .A1(net779),
    .A2(net342));
 sg13g2_o21ai_1 _16558_ (.B1(_09810_),
    .Y(_00081_),
    .A1(_09808_),
    .A2(_09809_));
 sg13g2_inv_2 _16559_ (.Y(_09811_),
    .A(_09079_));
 sg13g2_buf_1 _16560_ (.A(_09811_),
    .X(_09812_));
 sg13g2_buf_1 _16561_ (.A(net885),
    .X(_09813_));
 sg13g2_buf_1 _16562_ (.A(net772),
    .X(_09814_));
 sg13g2_buf_1 _16563_ (.A(net765),
    .X(_09815_));
 sg13g2_nand2_1 _16564_ (.Y(_09816_),
    .A(net670),
    .B(net669));
 sg13g2_buf_2 _16565_ (.A(_09816_),
    .X(_09817_));
 sg13g2_buf_2 _16566_ (.A(\cpu.addr[5] ),
    .X(_09818_));
 sg13g2_nor3_2 _16567_ (.A(_09818_),
    .B(net1038),
    .C(_09013_),
    .Y(_09819_));
 sg13g2_nand2_1 _16568_ (.Y(_09820_),
    .A(_09010_),
    .B(_09819_));
 sg13g2_buf_2 _16569_ (.A(_09820_),
    .X(_09821_));
 sg13g2_nor4_1 _16570_ (.A(net759),
    .B(_09109_),
    .C(_09817_),
    .D(_09821_),
    .Y(_09822_));
 sg13g2_buf_1 _16571_ (.A(_09822_),
    .X(_09823_));
 sg13g2_buf_1 _16572_ (.A(\cpu.intr.r_timer_count[12] ),
    .X(_09824_));
 sg13g2_buf_1 _16573_ (.A(\cpu.intr.r_timer_count[7] ),
    .X(_09825_));
 sg13g2_buf_2 _16574_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09826_));
 sg13g2_nor3_1 _16575_ (.A(_09826_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_09827_));
 sg13g2_nor2b_1 _16576_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_09827_),
    .Y(_09828_));
 sg13g2_nor2b_1 _16577_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09828_),
    .Y(_09829_));
 sg13g2_nor2b_1 _16578_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09829_),
    .Y(_09830_));
 sg13g2_nand2b_1 _16579_ (.Y(_09831_),
    .B(_09830_),
    .A_N(\cpu.intr.r_timer_count[6] ));
 sg13g2_nor3_1 _16580_ (.A(_09825_),
    .B(\cpu.intr.r_timer_count[8] ),
    .C(_09831_),
    .Y(_09832_));
 sg13g2_nor2b_1 _16581_ (.A(\cpu.intr.r_timer_count[9] ),
    .B_N(_09832_),
    .Y(_09833_));
 sg13g2_nor2b_1 _16582_ (.A(\cpu.intr.r_timer_count[10] ),
    .B_N(_09833_),
    .Y(_09834_));
 sg13g2_nand2b_1 _16583_ (.Y(_09835_),
    .B(_09834_),
    .A_N(\cpu.intr.r_timer_count[11] ));
 sg13g2_nor3_1 _16584_ (.A(\cpu.intr.r_timer_count[13] ),
    .B(_09824_),
    .C(_09835_),
    .Y(_09836_));
 sg13g2_nor2b_1 _16585_ (.A(\cpu.intr.r_timer_count[14] ),
    .B_N(_09836_),
    .Y(_09837_));
 sg13g2_nand2b_1 _16586_ (.Y(_09838_),
    .B(_09837_),
    .A_N(\cpu.intr.r_timer_count[15] ));
 sg13g2_buf_2 _16587_ (.A(_09838_),
    .X(_09839_));
 sg13g2_buf_1 _16588_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09840_));
 sg13g2_buf_1 _16589_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09841_));
 sg13g2_buf_1 _16590_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09842_));
 sg13g2_or4_1 _16591_ (.A(_09840_),
    .B(_09841_),
    .C(_09842_),
    .D(\cpu.intr.r_timer_count[19] ),
    .X(_09843_));
 sg13g2_or2_1 _16592_ (.X(_09844_),
    .B(_09843_),
    .A(_09839_));
 sg13g2_buf_2 _16593_ (.A(_09844_),
    .X(_09845_));
 sg13g2_buf_1 _16594_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_09846_));
 sg13g2_buf_1 _16595_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09847_));
 sg13g2_buf_1 _16596_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_09848_));
 sg13g2_buf_1 _16597_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09849_));
 sg13g2_or4_1 _16598_ (.A(_09846_),
    .B(_09847_),
    .C(_09848_),
    .D(_09849_),
    .X(_09850_));
 sg13g2_buf_1 _16599_ (.A(_09850_),
    .X(_09851_));
 sg13g2_or2_1 _16600_ (.X(_09852_),
    .B(_09851_),
    .A(_09845_));
 sg13g2_buf_2 _16601_ (.A(_09852_),
    .X(_09853_));
 sg13g2_inv_1 _16602_ (.Y(_09854_),
    .A(_09853_));
 sg13g2_nor2_1 _16603_ (.A(_09823_),
    .B(_09854_),
    .Y(_09855_));
 sg13g2_buf_1 _16604_ (.A(_09855_),
    .X(_09856_));
 sg13g2_buf_1 _16605_ (.A(_09856_),
    .X(_09857_));
 sg13g2_mux2_1 _16606_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(_00285_),
    .S(net68),
    .X(_00055_));
 sg13g2_xnor2_1 _16607_ (.Y(_09858_),
    .A(_09826_),
    .B(\cpu.intr.r_timer_count[0] ));
 sg13g2_mux2_1 _16608_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(_09858_),
    .S(net68),
    .X(_00066_));
 sg13g2_buf_1 _16609_ (.A(_09856_),
    .X(_09859_));
 sg13g2_o21ai_1 _16610_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_09860_),
    .A1(_09826_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16611_ (.A(_09827_),
    .B_N(_09860_),
    .Y(_09861_));
 sg13g2_nor2_1 _16612_ (.A(\cpu.intr.r_timer_reload[2] ),
    .B(net68),
    .Y(_09862_));
 sg13g2_a21oi_1 _16613_ (.A1(net67),
    .A2(_09861_),
    .Y(_00071_),
    .B1(_09862_));
 sg13g2_xnor2_1 _16614_ (.Y(_09863_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09827_));
 sg13g2_nor2_1 _16615_ (.A(\cpu.intr.r_timer_reload[3] ),
    .B(net68),
    .Y(_09864_));
 sg13g2_a21oi_1 _16616_ (.A1(net67),
    .A2(_09863_),
    .Y(_00072_),
    .B1(_09864_));
 sg13g2_xnor2_1 _16617_ (.Y(_09865_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09828_));
 sg13g2_nor2_1 _16618_ (.A(\cpu.intr.r_timer_reload[4] ),
    .B(net68),
    .Y(_09866_));
 sg13g2_a21oi_1 _16619_ (.A1(net67),
    .A2(_09865_),
    .Y(_00073_),
    .B1(_09866_));
 sg13g2_xnor2_1 _16620_ (.Y(_09867_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09829_));
 sg13g2_nor2_1 _16621_ (.A(\cpu.intr.r_timer_reload[5] ),
    .B(net68),
    .Y(_09868_));
 sg13g2_a21oi_1 _16622_ (.A1(net67),
    .A2(_09867_),
    .Y(_00074_),
    .B1(_09868_));
 sg13g2_xnor2_1 _16623_ (.Y(_09869_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09830_));
 sg13g2_buf_1 _16624_ (.A(_09856_),
    .X(_09870_));
 sg13g2_nor2_1 _16625_ (.A(\cpu.intr.r_timer_reload[6] ),
    .B(net66),
    .Y(_09871_));
 sg13g2_a21oi_1 _16626_ (.A1(net67),
    .A2(_09869_),
    .Y(_00075_),
    .B1(_09871_));
 sg13g2_xor2_1 _16627_ (.B(_09831_),
    .A(_09825_),
    .X(_09872_));
 sg13g2_nor2_1 _16628_ (.A(\cpu.intr.r_timer_reload[7] ),
    .B(net66),
    .Y(_09873_));
 sg13g2_a21oi_1 _16629_ (.A1(net67),
    .A2(_09872_),
    .Y(_00076_),
    .B1(_09873_));
 sg13g2_nor2_1 _16630_ (.A(_09825_),
    .B(_09831_),
    .Y(_09874_));
 sg13g2_xnor2_1 _16631_ (.Y(_09875_),
    .A(\cpu.intr.r_timer_count[8] ),
    .B(_09874_));
 sg13g2_nor2_1 _16632_ (.A(\cpu.intr.r_timer_reload[8] ),
    .B(net66),
    .Y(_09876_));
 sg13g2_a21oi_1 _16633_ (.A1(net67),
    .A2(_09875_),
    .Y(_00077_),
    .B1(_09876_));
 sg13g2_xnor2_1 _16634_ (.Y(_09877_),
    .A(\cpu.intr.r_timer_count[9] ),
    .B(_09832_));
 sg13g2_nor2_1 _16635_ (.A(\cpu.intr.r_timer_reload[9] ),
    .B(net66),
    .Y(_09878_));
 sg13g2_a21oi_1 _16636_ (.A1(net67),
    .A2(_09877_),
    .Y(_00078_),
    .B1(_09878_));
 sg13g2_xnor2_1 _16637_ (.Y(_09879_),
    .A(\cpu.intr.r_timer_count[10] ),
    .B(_09833_));
 sg13g2_nor2_1 _16638_ (.A(\cpu.intr.r_timer_reload[10] ),
    .B(net66),
    .Y(_09880_));
 sg13g2_a21oi_1 _16639_ (.A1(_09859_),
    .A2(_09879_),
    .Y(_00056_),
    .B1(_09880_));
 sg13g2_xnor2_1 _16640_ (.Y(_09881_),
    .A(\cpu.intr.r_timer_count[11] ),
    .B(_09834_));
 sg13g2_nor2_1 _16641_ (.A(\cpu.intr.r_timer_reload[11] ),
    .B(net66),
    .Y(_09882_));
 sg13g2_a21oi_1 _16642_ (.A1(_09859_),
    .A2(_09881_),
    .Y(_00057_),
    .B1(_09882_));
 sg13g2_xor2_1 _16643_ (.B(_09835_),
    .A(_09824_),
    .X(_09883_));
 sg13g2_nor2_1 _16644_ (.A(\cpu.intr.r_timer_reload[12] ),
    .B(net66),
    .Y(_09884_));
 sg13g2_a21oi_1 _16645_ (.A1(net68),
    .A2(_09883_),
    .Y(_00058_),
    .B1(_09884_));
 sg13g2_o21ai_1 _16646_ (.B1(\cpu.intr.r_timer_count[13] ),
    .Y(_09885_),
    .A1(_09824_),
    .A2(_09835_));
 sg13g2_nor2b_1 _16647_ (.A(_09836_),
    .B_N(_09885_),
    .Y(_09886_));
 sg13g2_nor2_1 _16648_ (.A(\cpu.intr.r_timer_reload[13] ),
    .B(net66),
    .Y(_09887_));
 sg13g2_a21oi_1 _16649_ (.A1(net68),
    .A2(_09886_),
    .Y(_00059_),
    .B1(_09887_));
 sg13g2_xnor2_1 _16650_ (.Y(_09888_),
    .A(\cpu.intr.r_timer_count[14] ),
    .B(_09836_));
 sg13g2_nor2_1 _16651_ (.A(\cpu.intr.r_timer_reload[14] ),
    .B(_09870_),
    .Y(_09889_));
 sg13g2_a21oi_1 _16652_ (.A1(_09857_),
    .A2(_09888_),
    .Y(_00060_),
    .B1(_09889_));
 sg13g2_xnor2_1 _16653_ (.Y(_09890_),
    .A(\cpu.intr.r_timer_count[15] ),
    .B(_09837_));
 sg13g2_nor2_1 _16654_ (.A(\cpu.intr.r_timer_reload[15] ),
    .B(_09870_),
    .Y(_09891_));
 sg13g2_a21oi_1 _16655_ (.A1(_09857_),
    .A2(_09890_),
    .Y(_00061_),
    .B1(_09891_));
 sg13g2_nor3_1 _16656_ (.A(\cpu.intr.r_timer_reload[16] ),
    .B(_09843_),
    .C(_09851_),
    .Y(_09892_));
 sg13g2_nor3_1 _16657_ (.A(_09841_),
    .B(_09839_),
    .C(_09892_),
    .Y(_09893_));
 sg13g2_a21o_1 _16658_ (.A2(_09839_),
    .A1(_09841_),
    .B1(_09893_),
    .X(_09894_));
 sg13g2_buf_1 _16659_ (.A(\cpu.dcache.wdata[0] ),
    .X(_09895_));
 sg13g2_buf_1 _16660_ (.A(_09895_),
    .X(_09896_));
 sg13g2_buf_1 _16661_ (.A(net1020),
    .X(_09897_));
 sg13g2_buf_1 _16662_ (.A(_09823_),
    .X(_09898_));
 sg13g2_mux2_1 _16663_ (.A0(_09894_),
    .A1(net884),
    .S(net105),
    .X(_00062_));
 sg13g2_buf_1 _16664_ (.A(_09823_),
    .X(_09899_));
 sg13g2_nor3_1 _16665_ (.A(_09840_),
    .B(_09841_),
    .C(_09839_),
    .Y(_09900_));
 sg13g2_o21ai_1 _16666_ (.B1(_09840_),
    .Y(_09901_),
    .A1(_09841_),
    .A2(_09839_));
 sg13g2_nand2b_1 _16667_ (.Y(_09902_),
    .B(_09901_),
    .A_N(_09900_));
 sg13g2_o21ai_1 _16668_ (.B1(_09902_),
    .Y(_09903_),
    .A1(\cpu.intr.r_timer_reload[17] ),
    .A2(_09853_));
 sg13g2_buf_1 _16669_ (.A(\cpu.dcache.wdata[1] ),
    .X(_09904_));
 sg13g2_buf_1 _16670_ (.A(_09904_),
    .X(_09905_));
 sg13g2_nand2_1 _16671_ (.Y(_09906_),
    .A(_09905_),
    .B(net105));
 sg13g2_o21ai_1 _16672_ (.B1(_09906_),
    .Y(_00063_),
    .A1(net104),
    .A2(_09903_));
 sg13g2_xor2_1 _16673_ (.B(_09900_),
    .A(_09842_),
    .X(_09907_));
 sg13g2_o21ai_1 _16674_ (.B1(_09907_),
    .Y(_09908_),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .A2(_09853_));
 sg13g2_buf_1 _16675_ (.A(\cpu.dcache.wdata[2] ),
    .X(_09909_));
 sg13g2_buf_1 _16676_ (.A(_09909_),
    .X(_09910_));
 sg13g2_nand2_1 _16677_ (.Y(_09911_),
    .A(net1018),
    .B(net105));
 sg13g2_o21ai_1 _16678_ (.B1(_09911_),
    .Y(_00064_),
    .A1(net104),
    .A2(_09908_));
 sg13g2_nor2b_1 _16679_ (.A(_09842_),
    .B_N(_09900_),
    .Y(_09912_));
 sg13g2_xor2_1 _16680_ (.B(_09912_),
    .A(\cpu.intr.r_timer_count[19] ),
    .X(_09913_));
 sg13g2_o21ai_1 _16681_ (.B1(_09913_),
    .Y(_09914_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09853_));
 sg13g2_buf_1 _16682_ (.A(\cpu.dcache.wdata[3] ),
    .X(_09915_));
 sg13g2_buf_1 _16683_ (.A(net1098),
    .X(_09916_));
 sg13g2_nand2_1 _16684_ (.Y(_09917_),
    .A(net1017),
    .B(net105));
 sg13g2_o21ai_1 _16685_ (.B1(_09917_),
    .Y(_00065_),
    .A1(net104),
    .A2(_09914_));
 sg13g2_nor2_1 _16686_ (.A(\cpu.intr.r_timer_reload[20] ),
    .B(_09851_),
    .Y(_09918_));
 sg13g2_nor3_1 _16687_ (.A(_09846_),
    .B(_09845_),
    .C(_09918_),
    .Y(_09919_));
 sg13g2_a21oi_1 _16688_ (.A1(_09846_),
    .A2(_09845_),
    .Y(_09920_),
    .B1(_09919_));
 sg13g2_buf_2 _16689_ (.A(\cpu.dcache.wdata[4] ),
    .X(_09921_));
 sg13g2_buf_1 _16690_ (.A(_09921_),
    .X(_09922_));
 sg13g2_nand2_1 _16691_ (.Y(_09923_),
    .A(net1016),
    .B(_09898_));
 sg13g2_o21ai_1 _16692_ (.B1(_09923_),
    .Y(_00067_),
    .A1(net104),
    .A2(_09920_));
 sg13g2_nor2_1 _16693_ (.A(_09846_),
    .B(_09845_),
    .Y(_09924_));
 sg13g2_xor2_1 _16694_ (.B(_09924_),
    .A(_09847_),
    .X(_09925_));
 sg13g2_o21ai_1 _16695_ (.B1(_09925_),
    .Y(_09926_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09853_));
 sg13g2_buf_2 _16696_ (.A(\cpu.dcache.wdata[5] ),
    .X(_09927_));
 sg13g2_buf_1 _16697_ (.A(_09927_),
    .X(_09928_));
 sg13g2_nand2_1 _16698_ (.Y(_09929_),
    .A(net1015),
    .B(_09823_));
 sg13g2_o21ai_1 _16699_ (.B1(_09929_),
    .Y(_00068_),
    .A1(_09898_),
    .A2(_09926_));
 sg13g2_nor3_1 _16700_ (.A(_09846_),
    .B(_09847_),
    .C(_09845_),
    .Y(_09930_));
 sg13g2_xor2_1 _16701_ (.B(_09930_),
    .A(_09848_),
    .X(_09931_));
 sg13g2_o21ai_1 _16702_ (.B1(_09931_),
    .Y(_09932_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_09853_));
 sg13g2_buf_2 _16703_ (.A(\cpu.dcache.wdata[6] ),
    .X(_09933_));
 sg13g2_buf_1 _16704_ (.A(_09933_),
    .X(_09934_));
 sg13g2_nand2_1 _16705_ (.Y(_09935_),
    .A(net1014),
    .B(_09823_));
 sg13g2_o21ai_1 _16706_ (.B1(_09935_),
    .Y(_00069_),
    .A1(net105),
    .A2(_09932_));
 sg13g2_nor2b_1 _16707_ (.A(_09848_),
    .B_N(_09930_),
    .Y(_09936_));
 sg13g2_nand2_1 _16708_ (.Y(_09937_),
    .A(\cpu.intr.r_timer_reload[23] ),
    .B(_09936_));
 sg13g2_nand2b_1 _16709_ (.Y(_09938_),
    .B(_09849_),
    .A_N(_09936_));
 sg13g2_o21ai_1 _16710_ (.B1(_09938_),
    .Y(_09939_),
    .A1(_09849_),
    .A2(_09937_));
 sg13g2_buf_2 _16711_ (.A(\cpu.dcache.wdata[7] ),
    .X(_09940_));
 sg13g2_buf_1 _16712_ (.A(_09940_),
    .X(_09941_));
 sg13g2_mux2_1 _16713_ (.A0(_09939_),
    .A1(net1013),
    .S(net105),
    .X(_00070_));
 sg13g2_buf_1 _16714_ (.A(net782),
    .X(_09942_));
 sg13g2_buf_1 _16715_ (.A(net668),
    .X(_09943_));
 sg13g2_buf_1 _16716_ (.A(net609),
    .X(_09944_));
 sg13g2_nor2b_1 _16717_ (.A(_09944_),
    .B_N(net1020),
    .Y(_09945_));
 sg13g2_nand2_1 _16718_ (.Y(_09946_),
    .A(_09130_),
    .B(_09283_));
 sg13g2_buf_1 _16719_ (.A(_09946_),
    .X(_09947_));
 sg13g2_nor3_1 _16720_ (.A(_09109_),
    .B(_09947_),
    .C(_09821_),
    .Y(_09948_));
 sg13g2_buf_1 _16721_ (.A(_09948_),
    .X(_09949_));
 sg13g2_buf_1 _16722_ (.A(_09949_),
    .X(_09950_));
 sg13g2_mux2_1 _16723_ (.A0(_00286_),
    .A1(_09945_),
    .S(net103),
    .X(_00036_));
 sg13g2_buf_1 _16724_ (.A(net1019),
    .X(_09951_));
 sg13g2_buf_2 _16725_ (.A(net759),
    .X(_09952_));
 sg13g2_and2_1 _16726_ (.A(net667),
    .B(net124),
    .X(_09953_));
 sg13g2_buf_1 _16727_ (.A(_09953_),
    .X(_09954_));
 sg13g2_buf_1 _16728_ (.A(_09954_),
    .X(_09955_));
 sg13g2_nor2_1 _16729_ (.A(_09109_),
    .B(_09821_),
    .Y(_09956_));
 sg13g2_buf_1 _16730_ (.A(_09956_),
    .X(_09957_));
 sg13g2_nand2_1 _16731_ (.Y(_09958_),
    .A(net1106),
    .B(net892));
 sg13g2_buf_1 _16732_ (.A(_09958_),
    .X(_09959_));
 sg13g2_nor3_1 _16733_ (.A(net891),
    .B(net619),
    .C(net666),
    .Y(_09960_));
 sg13g2_buf_1 _16734_ (.A(_09960_),
    .X(_09961_));
 sg13g2_buf_1 _16735_ (.A(_09961_),
    .X(_09962_));
 sg13g2_buf_1 _16736_ (.A(_09962_),
    .X(_09963_));
 sg13g2_and2_1 _16737_ (.A(net123),
    .B(net375),
    .X(_09964_));
 sg13g2_buf_1 _16738_ (.A(_09964_),
    .X(_09965_));
 sg13g2_buf_1 _16739_ (.A(net90),
    .X(_09966_));
 sg13g2_buf_1 _16740_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_09967_));
 sg13g2_buf_2 _16741_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_09968_));
 sg13g2_xnor2_1 _16742_ (.Y(_09969_),
    .A(_09967_),
    .B(_09968_));
 sg13g2_nor3_1 _16743_ (.A(net79),
    .B(net78),
    .C(_09969_),
    .Y(_09970_));
 sg13g2_a21o_1 _16744_ (.A2(net79),
    .A1(net883),
    .B1(_09970_),
    .X(_00043_));
 sg13g2_buf_1 _16745_ (.A(_09949_),
    .X(_09971_));
 sg13g2_buf_1 _16746_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_09972_));
 sg13g2_nand2_1 _16747_ (.Y(_09973_),
    .A(_09967_),
    .B(_09968_));
 sg13g2_xor2_1 _16748_ (.B(_09973_),
    .A(_09972_),
    .X(_09974_));
 sg13g2_buf_1 _16749_ (.A(net667),
    .X(_09975_));
 sg13g2_buf_1 _16750_ (.A(net608),
    .X(_09976_));
 sg13g2_nand3_1 _16751_ (.B(net1018),
    .C(net103),
    .A(net543),
    .Y(_09977_));
 sg13g2_o21ai_1 _16752_ (.B1(_09977_),
    .Y(_00044_),
    .A1(net102),
    .A2(_09974_));
 sg13g2_buf_1 _16753_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_09978_));
 sg13g2_nand2_1 _16754_ (.Y(_09979_),
    .A(_09968_),
    .B(_09972_));
 sg13g2_nor2_1 _16755_ (.A(_00286_),
    .B(_09979_),
    .Y(_09980_));
 sg13g2_xnor2_1 _16756_ (.Y(_09981_),
    .A(_09978_),
    .B(_09980_));
 sg13g2_nand3_1 _16757_ (.B(net1017),
    .C(net103),
    .A(net543),
    .Y(_09982_));
 sg13g2_o21ai_1 _16758_ (.B1(_09982_),
    .Y(_00045_),
    .A1(net102),
    .A2(_09981_));
 sg13g2_buf_2 _16759_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_09983_));
 sg13g2_nand4_1 _16760_ (.B(_09968_),
    .C(_09972_),
    .A(_09967_),
    .Y(_09984_),
    .D(_09978_));
 sg13g2_xor2_1 _16761_ (.B(_09984_),
    .A(_09983_),
    .X(_09985_));
 sg13g2_nand3_1 _16762_ (.B(net1016),
    .C(net103),
    .A(net543),
    .Y(_09986_));
 sg13g2_o21ai_1 _16763_ (.B1(_09986_),
    .Y(_00046_),
    .A1(net102),
    .A2(_09985_));
 sg13g2_buf_1 _16764_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_09987_));
 sg13g2_and3_1 _16765_ (.X(_09988_),
    .A(_09978_),
    .B(_09983_),
    .C(_09980_));
 sg13g2_xnor2_1 _16766_ (.Y(_09989_),
    .A(_09987_),
    .B(_09988_));
 sg13g2_nand3_1 _16767_ (.B(net1015),
    .C(net103),
    .A(net543),
    .Y(_09990_));
 sg13g2_o21ai_1 _16768_ (.B1(_09990_),
    .Y(_00047_),
    .A1(net102),
    .A2(_09989_));
 sg13g2_buf_1 _16769_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_09991_));
 sg13g2_nand2_1 _16770_ (.Y(_09992_),
    .A(_09983_),
    .B(_09987_));
 sg13g2_nor2_1 _16771_ (.A(_09984_),
    .B(_09992_),
    .Y(_09993_));
 sg13g2_xnor2_1 _16772_ (.Y(_09994_),
    .A(_09991_),
    .B(_09993_));
 sg13g2_nand3_1 _16773_ (.B(net1014),
    .C(net103),
    .A(net543),
    .Y(_09995_));
 sg13g2_o21ai_1 _16774_ (.B1(_09995_),
    .Y(_00048_),
    .A1(net102),
    .A2(_09994_));
 sg13g2_buf_2 _16775_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_09996_));
 sg13g2_nand3_1 _16776_ (.B(_09991_),
    .C(_09988_),
    .A(_09987_),
    .Y(_09997_));
 sg13g2_buf_1 _16777_ (.A(_09997_),
    .X(_09998_));
 sg13g2_xor2_1 _16778_ (.B(_09998_),
    .A(_09996_),
    .X(_09999_));
 sg13g2_buf_1 _16779_ (.A(_09940_),
    .X(_10000_));
 sg13g2_buf_1 _16780_ (.A(net124),
    .X(_10001_));
 sg13g2_nand3_1 _16781_ (.B(net1012),
    .C(net101),
    .A(net543),
    .Y(_10002_));
 sg13g2_o21ai_1 _16782_ (.B1(_10002_),
    .Y(_00049_),
    .A1(net102),
    .A2(_09999_));
 sg13g2_buf_2 _16783_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10003_));
 sg13g2_and2_1 _16784_ (.A(_09991_),
    .B(_09993_),
    .X(_10004_));
 sg13g2_buf_1 _16785_ (.A(_10004_),
    .X(_10005_));
 sg13g2_nand2_1 _16786_ (.Y(_10006_),
    .A(_09996_),
    .B(_10005_));
 sg13g2_xor2_1 _16787_ (.B(_10006_),
    .A(_10003_),
    .X(_10007_));
 sg13g2_buf_2 _16788_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10008_));
 sg13g2_nand3_1 _16789_ (.B(_10008_),
    .C(net101),
    .A(net543),
    .Y(_10009_));
 sg13g2_o21ai_1 _16790_ (.B1(_10009_),
    .Y(_00050_),
    .A1(_09971_),
    .A2(_10007_));
 sg13g2_buf_1 _16791_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10010_));
 sg13g2_nand3_1 _16792_ (.B(_10003_),
    .C(_10005_),
    .A(_09996_),
    .Y(_10011_));
 sg13g2_xor2_1 _16793_ (.B(_10011_),
    .A(_10010_),
    .X(_10012_));
 sg13g2_buf_2 _16794_ (.A(\cpu.dcache.wdata[9] ),
    .X(_10013_));
 sg13g2_nand3_1 _16795_ (.B(_10013_),
    .C(net101),
    .A(net543),
    .Y(_10014_));
 sg13g2_o21ai_1 _16796_ (.B1(_10014_),
    .Y(_00051_),
    .A1(net102),
    .A2(_10012_));
 sg13g2_buf_1 _16797_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10015_));
 sg13g2_nand4_1 _16798_ (.B(_10003_),
    .C(_10010_),
    .A(_09996_),
    .Y(_10016_),
    .D(_10005_));
 sg13g2_xor2_1 _16799_ (.B(_10016_),
    .A(_10015_),
    .X(_10017_));
 sg13g2_buf_2 _16800_ (.A(\cpu.dcache.wdata[10] ),
    .X(_10018_));
 sg13g2_nand3_1 _16801_ (.B(_10018_),
    .C(net101),
    .A(net608),
    .Y(_10019_));
 sg13g2_o21ai_1 _16802_ (.B1(_10019_),
    .Y(_00037_),
    .A1(_09971_),
    .A2(_10017_));
 sg13g2_buf_2 _16803_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10020_));
 sg13g2_and4_1 _16804_ (.A(_09996_),
    .B(_10003_),
    .C(_10010_),
    .D(_10015_),
    .X(_10021_));
 sg13g2_buf_1 _16805_ (.A(_10021_),
    .X(_10022_));
 sg13g2_nor2b_1 _16806_ (.A(_09998_),
    .B_N(_10022_),
    .Y(_10023_));
 sg13g2_xnor2_1 _16807_ (.Y(_10024_),
    .A(_10020_),
    .B(_10023_));
 sg13g2_buf_2 _16808_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10025_));
 sg13g2_nand3_1 _16809_ (.B(_10025_),
    .C(net101),
    .A(net608),
    .Y(_10026_));
 sg13g2_o21ai_1 _16810_ (.B1(_10026_),
    .Y(_00038_),
    .A1(net102),
    .A2(_10024_));
 sg13g2_buf_1 _16811_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10027_));
 sg13g2_nand3_1 _16812_ (.B(_10005_),
    .C(_10022_),
    .A(_10020_),
    .Y(_10028_));
 sg13g2_xor2_1 _16813_ (.B(_10028_),
    .A(_10027_),
    .X(_10029_));
 sg13g2_buf_2 _16814_ (.A(\cpu.dcache.wdata[12] ),
    .X(_10030_));
 sg13g2_nand3_1 _16815_ (.B(_10030_),
    .C(_10001_),
    .A(net608),
    .Y(_10031_));
 sg13g2_o21ai_1 _16816_ (.B1(_10031_),
    .Y(_00039_),
    .A1(net103),
    .A2(_10029_));
 sg13g2_buf_2 _16817_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10032_));
 sg13g2_nand3_1 _16818_ (.B(_10027_),
    .C(_10022_),
    .A(_10020_),
    .Y(_10033_));
 sg13g2_nor2_1 _16819_ (.A(_09998_),
    .B(_10033_),
    .Y(_10034_));
 sg13g2_xnor2_1 _16820_ (.Y(_10035_),
    .A(_10032_),
    .B(_10034_));
 sg13g2_buf_2 _16821_ (.A(\cpu.dcache.wdata[13] ),
    .X(_10036_));
 sg13g2_nand3_1 _16822_ (.B(_10036_),
    .C(_10001_),
    .A(net608),
    .Y(_10037_));
 sg13g2_o21ai_1 _16823_ (.B1(_10037_),
    .Y(_00040_),
    .A1(net103),
    .A2(_10035_));
 sg13g2_buf_2 _16824_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10038_));
 sg13g2_and4_1 _16825_ (.A(_10020_),
    .B(_10027_),
    .C(_10005_),
    .D(_10022_),
    .X(_10039_));
 sg13g2_buf_1 _16826_ (.A(_10039_),
    .X(_10040_));
 sg13g2_nand2_1 _16827_ (.Y(_10041_),
    .A(_10032_),
    .B(_10040_));
 sg13g2_xor2_1 _16828_ (.B(_10041_),
    .A(_10038_),
    .X(_10042_));
 sg13g2_buf_2 _16829_ (.A(\cpu.dcache.wdata[14] ),
    .X(_10043_));
 sg13g2_nand3_1 _16830_ (.B(_10043_),
    .C(net101),
    .A(net608),
    .Y(_10044_));
 sg13g2_o21ai_1 _16831_ (.B1(_10044_),
    .Y(_00041_),
    .A1(_09950_),
    .A2(_10042_));
 sg13g2_buf_1 _16832_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10045_));
 sg13g2_nand3_1 _16833_ (.B(_10038_),
    .C(_10034_),
    .A(_10032_),
    .Y(_10046_));
 sg13g2_xor2_1 _16834_ (.B(_10046_),
    .A(_10045_),
    .X(_10047_));
 sg13g2_buf_2 _16835_ (.A(\cpu.dcache.wdata[15] ),
    .X(_10048_));
 sg13g2_nand3_1 _16836_ (.B(_10048_),
    .C(net101),
    .A(net608),
    .Y(_10049_));
 sg13g2_o21ai_1 _16837_ (.B1(_10049_),
    .Y(_00042_),
    .A1(_09950_),
    .A2(_10047_));
 sg13g2_buf_1 _16838_ (.A(\cpu.ex.r_mult[0] ),
    .X(_10050_));
 sg13g2_buf_1 _16839_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10051_));
 sg13g2_buf_8 _16840_ (.A(_10051_),
    .X(_10052_));
 sg13g2_buf_2 _16841_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10053_));
 sg13g2_buf_1 _16842_ (.A(_10053_),
    .X(_10054_));
 sg13g2_buf_1 _16843_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10055_));
 sg13g2_buf_1 _16844_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10056_));
 sg13g2_buf_2 _16845_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10057_));
 sg13g2_inv_1 _16846_ (.Y(_10058_),
    .A(_10057_));
 sg13g2_nor2_1 _16847_ (.A(net1096),
    .B(_10058_),
    .Y(_10059_));
 sg13g2_nand4_1 _16848_ (.B(net1010),
    .C(net1097),
    .A(net1011),
    .Y(_10060_),
    .D(_10059_));
 sg13g2_buf_2 _16849_ (.A(_10060_),
    .X(_10061_));
 sg13g2_buf_1 _16850_ (.A(\cpu.ex.r_set_cc ),
    .X(_10062_));
 sg13g2_nand2_1 _16851_ (.Y(_10063_),
    .A(net1097),
    .B(_10062_));
 sg13g2_buf_1 _16852_ (.A(_10063_),
    .X(_10064_));
 sg13g2_and2_1 _16853_ (.A(_10061_),
    .B(_10064_),
    .X(_10065_));
 sg13g2_buf_1 _16854_ (.A(_10065_),
    .X(_10066_));
 sg13g2_nor2_2 _16855_ (.A(_09209_),
    .B(net1103),
    .Y(_10067_));
 sg13g2_nand2_2 _16856_ (.Y(_10068_),
    .A(_09207_),
    .B(_10067_));
 sg13g2_nand2_1 _16857_ (.Y(_10069_),
    .A(_10066_),
    .B(_10068_));
 sg13g2_buf_1 _16858_ (.A(_10069_),
    .X(_10070_));
 sg13g2_buf_1 _16859_ (.A(net428),
    .X(_10071_));
 sg13g2_buf_2 _16860_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10072_));
 sg13g2_inv_2 _16861_ (.Y(_10073_),
    .A(_10072_));
 sg13g2_buf_1 _16862_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10074_));
 sg13g2_buf_1 _16863_ (.A(net1095),
    .X(_10075_));
 sg13g2_buf_1 _16864_ (.A(_10075_),
    .X(_10076_));
 sg13g2_nand2_1 _16865_ (.Y(_10077_),
    .A(_08658_),
    .B(net882));
 sg13g2_buf_1 _16866_ (.A(\cpu.addr[11] ),
    .X(_10078_));
 sg13g2_buf_8 _16867_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10079_));
 sg13g2_xor2_1 _16868_ (.B(_10079_),
    .A(_10057_),
    .X(_10080_));
 sg13g2_buf_1 _16869_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10081_));
 sg13g2_xor2_1 _16870_ (.B(net1092),
    .A(_10052_),
    .X(_10082_));
 sg13g2_or2_1 _16871_ (.X(_10083_),
    .B(_10082_),
    .A(_10080_));
 sg13g2_buf_1 _16872_ (.A(_10083_),
    .X(_10084_));
 sg13g2_inv_1 _16873_ (.Y(_10085_),
    .A(net1097));
 sg13g2_buf_2 _16874_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10086_));
 sg13g2_xor2_1 _16875_ (.B(_10086_),
    .A(_10056_),
    .X(_10087_));
 sg13g2_buf_2 _16876_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10088_));
 sg13g2_xor2_1 _16877_ (.B(_10088_),
    .A(_10053_),
    .X(_10089_));
 sg13g2_nor4_1 _16878_ (.A(_10051_),
    .B(_10053_),
    .C(net1096),
    .D(_10057_),
    .Y(_10090_));
 sg13g2_or4_1 _16879_ (.A(_10085_),
    .B(_10087_),
    .C(_10089_),
    .D(_10090_),
    .X(_10091_));
 sg13g2_buf_1 _16880_ (.A(_10091_),
    .X(_10092_));
 sg13g2_nor2_1 _16881_ (.A(_10084_),
    .B(_10092_),
    .Y(_10093_));
 sg13g2_buf_2 _16882_ (.A(_10093_),
    .X(_10094_));
 sg13g2_buf_8 _16883_ (.A(_10094_),
    .X(_10095_));
 sg13g2_nor2_1 _16884_ (.A(_10080_),
    .B(_10082_),
    .Y(_10096_));
 sg13g2_nor4_1 _16885_ (.A(_10085_),
    .B(_10087_),
    .C(_10089_),
    .D(_10090_),
    .Y(_10097_));
 sg13g2_buf_8 _16886_ (.A(_10088_),
    .X(_10098_));
 sg13g2_nor2_1 _16887_ (.A(_10098_),
    .B(net1092),
    .Y(_10099_));
 sg13g2_buf_1 _16888_ (.A(_10099_),
    .X(_10100_));
 sg13g2_buf_8 _16889_ (.A(_10086_),
    .X(_10101_));
 sg13g2_nor2_1 _16890_ (.A(net1007),
    .B(_10079_),
    .Y(_10102_));
 sg13g2_buf_2 _16891_ (.A(_10102_),
    .X(_10103_));
 sg13g2_a22oi_1 _16892_ (.Y(_10104_),
    .B1(_10100_),
    .B2(_10103_),
    .A2(_10097_),
    .A1(_10096_));
 sg13g2_buf_1 _16893_ (.A(_10104_),
    .X(_10105_));
 sg13g2_buf_8 _16894_ (.A(_10105_),
    .X(_10106_));
 sg13g2_and2_1 _16895_ (.A(_10088_),
    .B(net1092),
    .X(_10107_));
 sg13g2_buf_1 _16896_ (.A(_10107_),
    .X(_10108_));
 sg13g2_inv_1 _16897_ (.Y(_10109_),
    .A(_00269_));
 sg13g2_a22oi_1 _16898_ (.Y(_10110_),
    .B1(_10108_),
    .B2(_10109_),
    .A2(net758),
    .A1(\cpu.ex.r_12[11] ));
 sg13g2_and2_1 _16899_ (.A(net1007),
    .B(net1093),
    .X(_10111_));
 sg13g2_buf_1 _16900_ (.A(_10111_),
    .X(_10112_));
 sg13g2_buf_1 _16901_ (.A(_10112_),
    .X(_10113_));
 sg13g2_nor2b_1 _16902_ (.A(_10110_),
    .B_N(net665),
    .Y(_10114_));
 sg13g2_buf_2 _16903_ (.A(net1092),
    .X(_10115_));
 sg13g2_buf_1 _16904_ (.A(_10115_),
    .X(_10116_));
 sg13g2_buf_1 _16905_ (.A(_10116_),
    .X(_10117_));
 sg13g2_buf_1 _16906_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10118_));
 sg13g2_buf_2 _16907_ (.A(net1093),
    .X(_10119_));
 sg13g2_buf_1 _16908_ (.A(net1005),
    .X(_10120_));
 sg13g2_buf_1 _16909_ (.A(_10101_),
    .X(_10121_));
 sg13g2_buf_1 _16910_ (.A(net879),
    .X(_10122_));
 sg13g2_mux4_1 _16911_ (.S0(net880),
    .A0(_10118_),
    .A1(\cpu.ex.r_stmp[11] ),
    .A2(\cpu.ex.r_10[11] ),
    .A3(\cpu.ex.r_14[11] ),
    .S1(net756),
    .X(_10123_));
 sg13g2_nand2_1 _16912_ (.Y(_10124_),
    .A(_10117_),
    .B(_10123_));
 sg13g2_inv_1 _16913_ (.Y(_10125_),
    .A(net1005));
 sg13g2_buf_1 _16914_ (.A(_10125_),
    .X(_10126_));
 sg13g2_nor2b_1 _16915_ (.A(_10081_),
    .B_N(_10086_),
    .Y(_10127_));
 sg13g2_buf_1 _16916_ (.A(_10127_),
    .X(_10128_));
 sg13g2_buf_1 _16917_ (.A(_10128_),
    .X(_10129_));
 sg13g2_nand3_1 _16918_ (.B(net755),
    .C(net754),
    .A(\cpu.ex.r_8[11] ),
    .Y(_10130_));
 sg13g2_buf_1 _16919_ (.A(net1008),
    .X(_10131_));
 sg13g2_buf_1 _16920_ (.A(net878),
    .X(_10132_));
 sg13g2_buf_1 _16921_ (.A(net753),
    .X(_10133_));
 sg13g2_a21oi_1 _16922_ (.A1(_10124_),
    .A2(_10130_),
    .Y(_10134_),
    .B1(net664));
 sg13g2_nor2b_1 _16923_ (.A(net1007),
    .B_N(net1092),
    .Y(_10135_));
 sg13g2_buf_1 _16924_ (.A(_10135_),
    .X(_10136_));
 sg13g2_buf_1 _16925_ (.A(_10136_),
    .X(_10137_));
 sg13g2_a22oi_1 _16926_ (.Y(_10138_),
    .B1(net663),
    .B2(\cpu.ex.r_epc[11] ),
    .A2(net754),
    .A1(\cpu.ex.r_9[11] ));
 sg13g2_nor2b_1 _16927_ (.A(net1093),
    .B_N(_10088_),
    .Y(_10139_));
 sg13g2_buf_1 _16928_ (.A(_10139_),
    .X(_10140_));
 sg13g2_nor2b_1 _16929_ (.A(_10138_),
    .B_N(net877),
    .Y(_10141_));
 sg13g2_inv_2 _16930_ (.Y(_10142_),
    .A(net1008));
 sg13g2_buf_1 _16931_ (.A(_10142_),
    .X(_10143_));
 sg13g2_buf_1 _16932_ (.A(net752),
    .X(_10144_));
 sg13g2_a221oi_1 _16933_ (.B2(\cpu.ex.r_13[11] ),
    .C1(_10117_),
    .B1(_10113_),
    .A1(\cpu.ex.r_lr[11] ),
    .Y(_10145_),
    .A2(_10103_));
 sg13g2_nor2b_1 _16934_ (.A(net1005),
    .B_N(net1007),
    .Y(_10146_));
 sg13g2_buf_1 _16935_ (.A(_10146_),
    .X(_10147_));
 sg13g2_buf_1 _16936_ (.A(net1007),
    .X(_10148_));
 sg13g2_buf_1 _16937_ (.A(_10119_),
    .X(_10149_));
 sg13g2_nor2b_1 _16938_ (.A(net876),
    .B_N(net875),
    .Y(_10150_));
 sg13g2_buf_8 _16939_ (.A(net1006),
    .X(_10151_));
 sg13g2_inv_2 _16940_ (.Y(_10152_),
    .A(net874));
 sg13g2_buf_8 _16941_ (.A(_10152_),
    .X(_10153_));
 sg13g2_a221oi_1 _16942_ (.B2(\cpu.ex.r_mult[27] ),
    .C1(net661),
    .B1(_10150_),
    .A1(\cpu.ex.r_11[11] ),
    .Y(_10154_),
    .A2(net751));
 sg13g2_nor3_1 _16943_ (.A(net662),
    .B(_10145_),
    .C(_10154_),
    .Y(_10155_));
 sg13g2_or4_1 _16944_ (.A(_10114_),
    .B(_10134_),
    .C(_10141_),
    .D(_10155_),
    .X(_10156_));
 sg13g2_buf_2 _16945_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10157_));
 sg13g2_inv_1 _16946_ (.Y(_10158_),
    .A(_10157_));
 sg13g2_buf_1 _16947_ (.A(_10158_),
    .X(_10159_));
 sg13g2_a221oi_1 _16948_ (.B2(_10156_),
    .C1(net873),
    .B1(net541),
    .A1(net1094),
    .Y(_10160_),
    .A2(net492));
 sg13g2_buf_1 _16949_ (.A(_10157_),
    .X(_10161_));
 sg13g2_nor2_1 _16950_ (.A(net1004),
    .B(\cpu.dec.imm[11] ),
    .Y(_10162_));
 sg13g2_buf_2 _16951_ (.A(\cpu.dec.r_rs2_inv ),
    .X(_10163_));
 sg13g2_nor2_1 _16952_ (.A(net1095),
    .B(_10163_),
    .Y(_10164_));
 sg13g2_buf_1 _16953_ (.A(_10164_),
    .X(_10165_));
 sg13g2_o21ai_1 _16954_ (.B1(_10165_),
    .Y(_10166_),
    .A1(_10160_),
    .A2(_10162_));
 sg13g2_buf_1 _16955_ (.A(_10166_),
    .X(_10167_));
 sg13g2_and2_1 _16956_ (.A(_10077_),
    .B(_10167_),
    .X(_10168_));
 sg13g2_buf_2 _16957_ (.A(_10168_),
    .X(_10169_));
 sg13g2_buf_1 _16958_ (.A(_00301_),
    .X(_10170_));
 sg13g2_a21oi_1 _16959_ (.A1(_10073_),
    .A2(_10169_),
    .Y(_10171_),
    .B1(_10170_));
 sg13g2_or3_1 _16960_ (.A(_09196_),
    .B(_09210_),
    .C(\cpu.ex.r_mult_off[2] ),
    .X(_10172_));
 sg13g2_o21ai_1 _16961_ (.B1(\cpu.ex.r_mult_off[2] ),
    .Y(_10173_),
    .A1(_09196_),
    .A2(_09210_));
 sg13g2_and3_1 _16962_ (.X(_10174_),
    .A(_09207_),
    .B(_10172_),
    .C(_10173_));
 sg13g2_buf_2 _16963_ (.A(_10174_),
    .X(_10175_));
 sg13g2_buf_2 _16964_ (.A(\cpu.br ),
    .X(_10176_));
 sg13g2_xor2_1 _16965_ (.B(_09210_),
    .A(_09196_),
    .X(_10177_));
 sg13g2_and2_1 _16966_ (.A(_09207_),
    .B(_10177_),
    .X(_10178_));
 sg13g2_buf_2 _16967_ (.A(_10178_),
    .X(_10179_));
 sg13g2_inv_2 _16968_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_10179_));
 sg13g2_nor2_1 _16969_ (.A(net495),
    .B(\cpu.ex.c_mult_off[1] ),
    .Y(_10180_));
 sg13g2_nor2_1 _16970_ (.A(_09018_),
    .B(_09075_),
    .Y(_10181_));
 sg13g2_nand2_1 _16971_ (.Y(_10182_),
    .A(net379),
    .B(_10181_));
 sg13g2_buf_1 _16972_ (.A(_10182_),
    .X(_10183_));
 sg13g2_nand4_1 _16973_ (.B(_10176_),
    .C(_10180_),
    .A(_08738_),
    .Y(_10184_),
    .D(_10183_));
 sg13g2_inv_1 _16974_ (.Y(_10185_),
    .A(_09071_));
 sg13g2_nor2_1 _16975_ (.A(_10185_),
    .B(_09074_),
    .Y(_10186_));
 sg13g2_o21ai_1 _16976_ (.B1(_10186_),
    .Y(_10187_),
    .A1(_09060_),
    .A2(_09070_));
 sg13g2_a21oi_1 _16977_ (.A1(_09073_),
    .A2(_09040_),
    .Y(_10188_),
    .B1(_09018_));
 sg13g2_buf_1 _16978_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10189_));
 sg13g2_buf_1 _16979_ (.A(_10189_),
    .X(_10190_));
 sg13g2_buf_2 _16980_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10191_));
 sg13g2_buf_1 _16981_ (.A(_10191_),
    .X(_10192_));
 sg13g2_nor2_1 _16982_ (.A(net1003),
    .B(net1002),
    .Y(_10193_));
 sg13g2_buf_2 _16983_ (.A(_10193_),
    .X(_10194_));
 sg13g2_buf_2 _16984_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10195_));
 sg13g2_buf_8 _16985_ (.A(_10195_),
    .X(_10196_));
 sg13g2_buf_1 _16986_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10197_));
 sg13g2_nor2_1 _16987_ (.A(_10196_),
    .B(_10197_),
    .Y(_10198_));
 sg13g2_buf_2 _16988_ (.A(_10198_),
    .X(_10199_));
 sg13g2_a21oi_1 _16989_ (.A1(_10194_),
    .A2(_10199_),
    .Y(_10200_),
    .B1(_00273_));
 sg13g2_and3_1 _16990_ (.X(_10201_),
    .A(_10187_),
    .B(_10188_),
    .C(_10200_));
 sg13g2_buf_2 _16991_ (.A(_10201_),
    .X(_10202_));
 sg13g2_inv_1 _16992_ (.Y(_10203_),
    .A(_10176_));
 sg13g2_a21oi_1 _16993_ (.A1(net379),
    .A2(_10202_),
    .Y(_10204_),
    .B1(_10203_));
 sg13g2_buf_2 _16994_ (.A(_10204_),
    .X(_10205_));
 sg13g2_buf_2 _16995_ (.A(_00200_),
    .X(_10206_));
 sg13g2_inv_1 _16996_ (.Y(_10207_),
    .A(_10206_));
 sg13g2_nand2_1 _16997_ (.Y(_10208_),
    .A(_10207_),
    .B(_10179_));
 sg13g2_o21ai_1 _16998_ (.B1(_10208_),
    .Y(_10209_),
    .A1(_00191_),
    .A2(_10179_));
 sg13g2_nand3_1 _16999_ (.B(_10205_),
    .C(_10209_),
    .A(net495),
    .Y(_10210_));
 sg13g2_nand2b_1 _17000_ (.Y(_10211_),
    .B(net1097),
    .A_N(_10090_));
 sg13g2_xnor2_1 _17001_ (.Y(_10212_),
    .A(net1096),
    .B(_10195_));
 sg13g2_xnor2_1 _17002_ (.Y(_10213_),
    .A(_10053_),
    .B(_10189_));
 sg13g2_nand2_1 _17003_ (.Y(_10214_),
    .A(_10212_),
    .B(_10213_));
 sg13g2_xnor2_1 _17004_ (.Y(_10215_),
    .A(_10057_),
    .B(net1091));
 sg13g2_xnor2_1 _17005_ (.Y(_10216_),
    .A(net1011),
    .B(_10191_));
 sg13g2_nand2_1 _17006_ (.Y(_10217_),
    .A(_10215_),
    .B(_10216_));
 sg13g2_or3_1 _17007_ (.A(_10211_),
    .B(_10214_),
    .C(_10217_),
    .X(_10218_));
 sg13g2_buf_1 _17008_ (.A(_10218_),
    .X(_10219_));
 sg13g2_buf_1 _17009_ (.A(_10219_),
    .X(_10220_));
 sg13g2_buf_1 _17010_ (.A(_10220_),
    .X(_10221_));
 sg13g2_nor2_1 _17011_ (.A(_09090_),
    .B(net491),
    .Y(_10222_));
 sg13g2_nor3_1 _17012_ (.A(_10211_),
    .B(_10214_),
    .C(_10217_),
    .Y(_10223_));
 sg13g2_buf_1 _17013_ (.A(_10223_),
    .X(_10224_));
 sg13g2_inv_1 _17014_ (.Y(_10225_),
    .A(_10192_));
 sg13g2_buf_1 _17015_ (.A(_10225_),
    .X(_10226_));
 sg13g2_buf_8 _17016_ (.A(net1091),
    .X(_10227_));
 sg13g2_inv_2 _17017_ (.Y(_10228_),
    .A(net1000));
 sg13g2_buf_1 _17018_ (.A(_10228_),
    .X(_10229_));
 sg13g2_nor2b_1 _17019_ (.A(net1003),
    .B_N(net1001),
    .Y(_10230_));
 sg13g2_buf_1 _17020_ (.A(_10230_),
    .X(_10231_));
 sg13g2_and2_1 _17021_ (.A(net749),
    .B(net748),
    .X(_10232_));
 sg13g2_buf_1 _17022_ (.A(net1001),
    .X(_10233_));
 sg13g2_buf_8 _17023_ (.A(_10233_),
    .X(_10234_));
 sg13g2_buf_8 _17024_ (.A(net747),
    .X(_10235_));
 sg13g2_buf_8 _17025_ (.A(_10190_),
    .X(_10236_));
 sg13g2_buf_8 _17026_ (.A(_10236_),
    .X(_10237_));
 sg13g2_buf_8 _17027_ (.A(net1000),
    .X(_10238_));
 sg13g2_buf_1 _17028_ (.A(_10238_),
    .X(_10239_));
 sg13g2_nand2_1 _17029_ (.Y(_10240_),
    .A(net746),
    .B(net745));
 sg13g2_nor2_1 _17030_ (.A(net660),
    .B(_10240_),
    .Y(_10241_));
 sg13g2_buf_2 _17031_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10242_));
 sg13g2_a22oi_1 _17032_ (.Y(_10243_),
    .B1(_10241_),
    .B2(_10242_),
    .A2(_10232_),
    .A1(\cpu.ex.r_8[3] ));
 sg13g2_buf_1 _17033_ (.A(_10199_),
    .X(_10244_));
 sg13g2_buf_1 _17034_ (.A(_10237_),
    .X(_10245_));
 sg13g2_buf_1 _17035_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10246_));
 sg13g2_nor2b_1 _17036_ (.A(net658),
    .B_N(_10246_),
    .Y(_10247_));
 sg13g2_buf_1 _17037_ (.A(net749),
    .X(_10248_));
 sg13g2_nor2_1 _17038_ (.A(net657),
    .B(_00261_),
    .Y(_10249_));
 sg13g2_and2_1 _17039_ (.A(net871),
    .B(net872),
    .X(_10250_));
 sg13g2_buf_1 _17040_ (.A(_10250_),
    .X(_10251_));
 sg13g2_a221oi_1 _17041_ (.B2(_10251_),
    .C1(net750),
    .B1(_10249_),
    .A1(net659),
    .Y(_10252_),
    .A2(_10247_));
 sg13g2_a21oi_1 _17042_ (.A1(_10226_),
    .A2(_10243_),
    .Y(_10253_),
    .B1(_10252_));
 sg13g2_inv_1 _17043_ (.Y(_10254_),
    .A(net1001));
 sg13g2_buf_1 _17044_ (.A(_10254_),
    .X(_10255_));
 sg13g2_nor2b_1 _17045_ (.A(net871),
    .B_N(net1000),
    .Y(_10256_));
 sg13g2_buf_1 _17046_ (.A(_10256_),
    .X(_10257_));
 sg13g2_buf_8 _17047_ (.A(net1002),
    .X(_10258_));
 sg13g2_buf_8 _17048_ (.A(net869),
    .X(_10259_));
 sg13g2_mux2_1 _17049_ (.A0(\cpu.ex.r_12[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net743),
    .X(_10260_));
 sg13g2_inv_1 _17050_ (.Y(_10261_),
    .A(\cpu.ex.r_10[3] ));
 sg13g2_nand2b_1 _17051_ (.Y(_10262_),
    .B(_10191_),
    .A_N(_10189_));
 sg13g2_buf_2 _17052_ (.A(_10262_),
    .X(_10263_));
 sg13g2_nand3b_1 _17053_ (.B(\cpu.ex.r_9[3] ),
    .C(net746),
    .Y(_10264_),
    .A_N(net743));
 sg13g2_o21ai_1 _17054_ (.B1(_10264_),
    .Y(_10265_),
    .A1(_10261_),
    .A2(_10263_));
 sg13g2_buf_1 _17055_ (.A(net870),
    .X(_10266_));
 sg13g2_nand3b_1 _17056_ (.B(_10266_),
    .C(\cpu.ex.r_13[3] ),
    .Y(_10267_),
    .A_N(net743));
 sg13g2_nand3b_1 _17057_ (.B(\cpu.ex.r_11[3] ),
    .C(net743),
    .Y(_10268_),
    .A_N(net745));
 sg13g2_inv_1 _17058_ (.Y(_10269_),
    .A(net1003));
 sg13g2_buf_1 _17059_ (.A(_10269_),
    .X(_10270_));
 sg13g2_a21oi_1 _17060_ (.A1(_10267_),
    .A2(_10268_),
    .Y(_10271_),
    .B1(net741));
 sg13g2_a221oi_1 _17061_ (.B2(net657),
    .C1(_10271_),
    .B1(_10265_),
    .A1(_10257_),
    .Y(_10272_),
    .A2(_10260_));
 sg13g2_nor2_1 _17062_ (.A(_10255_),
    .B(_10272_),
    .Y(_10273_));
 sg13g2_nor2_1 _17063_ (.A(net749),
    .B(_10263_),
    .Y(_10274_));
 sg13g2_buf_1 _17064_ (.A(net745),
    .X(_10275_));
 sg13g2_nor2_1 _17065_ (.A(_10270_),
    .B(net656),
    .Y(_10276_));
 sg13g2_buf_2 _17066_ (.A(net869),
    .X(_10277_));
 sg13g2_mux2_1 _17067_ (.A0(\cpu.ex.r_lr[3] ),
    .A1(\cpu.ex.r_epc[3] ),
    .S(_10277_),
    .X(_10278_));
 sg13g2_a22oi_1 _17068_ (.Y(_10279_),
    .B1(_10276_),
    .B2(_10278_),
    .A2(_10274_),
    .A1(\cpu.ex.r_stmp[3] ));
 sg13g2_and2_1 _17069_ (.A(net871),
    .B(net1002),
    .X(_10280_));
 sg13g2_buf_1 _17070_ (.A(_10280_),
    .X(_10281_));
 sg13g2_a22oi_1 _17071_ (.Y(_10282_),
    .B1(_10281_),
    .B2(\cpu.ex.r_mult[19] ),
    .A2(_10194_),
    .A1(net1115));
 sg13g2_nand2b_1 _17072_ (.Y(_10283_),
    .B(net656),
    .A_N(_10282_));
 sg13g2_a21oi_1 _17073_ (.A1(_10279_),
    .A2(_10283_),
    .Y(_10284_),
    .B1(net660));
 sg13g2_nor4_2 _17074_ (.A(net607),
    .B(_10253_),
    .C(_10273_),
    .Y(_10285_),
    .D(_10284_));
 sg13g2_nand2_1 _17075_ (.Y(_10286_),
    .A(net495),
    .B(\cpu.ex.c_mult_off[1] ));
 sg13g2_nor3_1 _17076_ (.A(_10222_),
    .B(_10285_),
    .C(_10286_),
    .Y(_10287_));
 sg13g2_buf_1 _17077_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10288_));
 sg13g2_mux2_1 _17078_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.mmu_read[1] ),
    .S(net870),
    .X(_10289_));
 sg13g2_a22oi_1 _17079_ (.Y(_10290_),
    .B1(_10289_),
    .B2(net658),
    .A2(_10257_),
    .A1(_10288_));
 sg13g2_nand3_1 _17080_ (.B(\cpu.ex.r_8[1] ),
    .C(net748),
    .A(net749),
    .Y(_10291_));
 sg13g2_o21ai_1 _17081_ (.B1(_10291_),
    .Y(_10292_),
    .A1(net660),
    .A2(_10290_));
 sg13g2_nand3_1 _17082_ (.B(\cpu.ex.r_11[1] ),
    .C(_10251_),
    .A(net657),
    .Y(_10293_));
 sg13g2_buf_1 _17083_ (.A(net872),
    .X(_10294_));
 sg13g2_mux2_1 _17084_ (.A0(\cpu.ex.r_stmp[1] ),
    .A1(\cpu.ex.r_14[1] ),
    .S(_10294_),
    .X(_10295_));
 sg13g2_nand2_1 _17085_ (.Y(_10296_),
    .A(_10257_),
    .B(_10295_));
 sg13g2_nand3_1 _17086_ (.B(_10293_),
    .C(_10296_),
    .A(net740),
    .Y(_10297_));
 sg13g2_o21ai_1 _17087_ (.B1(_10297_),
    .Y(_10298_),
    .A1(net740),
    .A2(_10292_));
 sg13g2_nand2_1 _17088_ (.Y(_10299_),
    .A(net743),
    .B(_10234_));
 sg13g2_nor2_1 _17089_ (.A(net871),
    .B(_10227_),
    .Y(_10300_));
 sg13g2_buf_2 _17090_ (.A(_10300_),
    .X(_10301_));
 sg13g2_and2_1 _17091_ (.A(net1003),
    .B(net1091),
    .X(_10302_));
 sg13g2_buf_2 _17092_ (.A(_10302_),
    .X(_10303_));
 sg13g2_inv_1 _17093_ (.Y(_10304_),
    .A(_00259_));
 sg13g2_a22oi_1 _17094_ (.Y(_10305_),
    .B1(_10303_),
    .B2(_10304_),
    .A2(_10301_),
    .A1(\cpu.ex.r_10[1] ));
 sg13g2_nor2_1 _17095_ (.A(_10299_),
    .B(_10305_),
    .Y(_10306_));
 sg13g2_and2_1 _17096_ (.A(net870),
    .B(\cpu.ex.r_mult[17] ),
    .X(_10307_));
 sg13g2_a21oi_1 _17097_ (.A1(net749),
    .A2(\cpu.ex.r_epc[1] ),
    .Y(_10308_),
    .B1(_10307_));
 sg13g2_nand2_1 _17098_ (.Y(_10309_),
    .A(net744),
    .B(net655));
 sg13g2_nor2b_1 _17099_ (.A(net1002),
    .B_N(_10195_),
    .Y(_10310_));
 sg13g2_buf_1 _17100_ (.A(_10310_),
    .X(_10311_));
 sg13g2_nand3_1 _17101_ (.B(_10257_),
    .C(_10311_),
    .A(\cpu.ex.r_12[1] ),
    .Y(_10312_));
 sg13g2_o21ai_1 _17102_ (.B1(_10312_),
    .Y(_10313_),
    .A1(_10308_),
    .A2(_10309_));
 sg13g2_buf_8 _17103_ (.A(_10238_),
    .X(_10314_));
 sg13g2_nand2b_1 _17104_ (.Y(_10315_),
    .B(_10314_),
    .A_N(\cpu.ex.r_13[1] ));
 sg13g2_o21ai_1 _17105_ (.B1(_10315_),
    .Y(_10316_),
    .A1(_10239_),
    .A2(\cpu.ex.r_9[1] ));
 sg13g2_nand2_1 _17106_ (.Y(_10317_),
    .A(net746),
    .B(_10311_));
 sg13g2_buf_1 _17107_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10318_));
 sg13g2_nor2b_1 _17108_ (.A(net871),
    .B_N(net1002),
    .Y(_10319_));
 sg13g2_buf_1 _17109_ (.A(_10319_),
    .X(_10320_));
 sg13g2_nand3_1 _17110_ (.B(net659),
    .C(net654),
    .A(_10318_),
    .Y(_10321_));
 sg13g2_o21ai_1 _17111_ (.B1(_10321_),
    .Y(_10322_),
    .A1(_10316_),
    .A2(_10317_));
 sg13g2_nor4_2 _17112_ (.A(net607),
    .B(_10306_),
    .C(_10313_),
    .Y(_10323_),
    .D(_10322_));
 sg13g2_nor2_1 _17113_ (.A(_09079_),
    .B(net540),
    .Y(_10324_));
 sg13g2_a21oi_2 _17114_ (.B1(_10324_),
    .Y(_10325_),
    .A2(_10323_),
    .A1(_10298_));
 sg13g2_and2_1 _17115_ (.A(_09208_),
    .B(_10179_),
    .X(_10326_));
 sg13g2_nor2_1 _17116_ (.A(_08767_),
    .B(_10220_),
    .Y(_10327_));
 sg13g2_nor2b_1 _17117_ (.A(_10195_),
    .B_N(net1091),
    .Y(_10328_));
 sg13g2_buf_2 _17118_ (.A(_10328_),
    .X(_10329_));
 sg13g2_mux2_1 _17119_ (.A0(\cpu.ex.r_8[0] ),
    .A1(\cpu.ex.r_12[0] ),
    .S(net870),
    .X(_10330_));
 sg13g2_a22oi_1 _17120_ (.Y(_10331_),
    .B1(_10330_),
    .B2(net747),
    .A2(_10329_),
    .A1(_09073_));
 sg13g2_nand2b_1 _17121_ (.Y(_10332_),
    .B(_10194_),
    .A_N(_10331_));
 sg13g2_nand2_2 _17122_ (.Y(_10333_),
    .A(_10195_),
    .B(net1091));
 sg13g2_nor2_1 _17123_ (.A(_10333_),
    .B(_10263_),
    .Y(_10334_));
 sg13g2_mux2_1 _17124_ (.A0(\cpu.ex.r_9[0] ),
    .A1(\cpu.ex.r_13[0] ),
    .S(net870),
    .X(_10335_));
 sg13g2_nand2b_1 _17125_ (.Y(_10336_),
    .B(net871),
    .A_N(net1002));
 sg13g2_buf_1 _17126_ (.A(_10336_),
    .X(_10337_));
 sg13g2_nor2_1 _17127_ (.A(net744),
    .B(_10337_),
    .Y(_10338_));
 sg13g2_nand3b_1 _17128_ (.B(\cpu.ex.r_10[0] ),
    .C(net872),
    .Y(_10339_),
    .A_N(net870));
 sg13g2_nand3b_1 _17129_ (.B(net870),
    .C(\cpu.ex.r_stmp[0] ),
    .Y(_10340_),
    .A_N(net872));
 sg13g2_a21oi_1 _17130_ (.A1(_10339_),
    .A2(_10340_),
    .Y(_10341_),
    .B1(_10263_));
 sg13g2_a221oi_1 _17131_ (.B2(_10338_),
    .C1(_10341_),
    .B1(_10335_),
    .A1(\cpu.ex.r_14[0] ),
    .Y(_10342_),
    .A2(_10334_));
 sg13g2_buf_1 _17132_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10343_));
 sg13g2_mux4_1 _17133_ (.S0(net872),
    .A0(_10343_),
    .A1(\cpu.ex.r_11[0] ),
    .A2(\cpu.ex.r_mult[16] ),
    .A3(\cpu.ex.r_15[0] ),
    .S1(net738),
    .X(_10344_));
 sg13g2_nand2_1 _17134_ (.Y(_10345_),
    .A(net655),
    .B(_10344_));
 sg13g2_and4_1 _17135_ (.A(_10219_),
    .B(_10332_),
    .C(_10342_),
    .D(_10345_),
    .X(_10346_));
 sg13g2_buf_1 _17136_ (.A(_10346_),
    .X(_10347_));
 sg13g2_nor4_1 _17137_ (.A(_09208_),
    .B(\cpu.ex.c_mult_off[1] ),
    .C(_10327_),
    .D(_10347_),
    .Y(_10348_));
 sg13g2_a21o_1 _17138_ (.A2(_10326_),
    .A1(_10325_),
    .B1(_10348_),
    .X(_10349_));
 sg13g2_a21o_1 _17139_ (.A2(_10202_),
    .A1(_08836_),
    .B1(_10203_),
    .X(_10350_));
 sg13g2_buf_8 _17140_ (.A(_10350_),
    .X(_10351_));
 sg13g2_o21ai_1 _17141_ (.B1(_10351_),
    .Y(_10352_),
    .A1(_10287_),
    .A2(_10349_));
 sg13g2_nor2_1 _17142_ (.A(net495),
    .B(_10179_),
    .Y(_10353_));
 sg13g2_nand2_1 _17143_ (.Y(_10354_),
    .A(_09351_),
    .B(net607));
 sg13g2_mux2_1 _17144_ (.A0(\cpu.ex.r_9[2] ),
    .A1(\cpu.ex.r_13[2] ),
    .S(net742),
    .X(_10355_));
 sg13g2_nand2_1 _17145_ (.Y(_10356_),
    .A(\cpu.ex.r_10[2] ),
    .B(_10301_));
 sg13g2_o21ai_1 _17146_ (.B1(_10356_),
    .Y(_10357_),
    .A1(_00260_),
    .A2(_10240_));
 sg13g2_and2_1 _17147_ (.A(_10191_),
    .B(_10195_),
    .X(_10358_));
 sg13g2_buf_1 _17148_ (.A(_10358_),
    .X(_10359_));
 sg13g2_a22oi_1 _17149_ (.Y(_10360_),
    .B1(_10357_),
    .B2(_10359_),
    .A2(_10355_),
    .A1(_10338_));
 sg13g2_nor2_1 _17150_ (.A(net869),
    .B(net872),
    .Y(_10361_));
 sg13g2_a22oi_1 _17151_ (.Y(_10362_),
    .B1(_10361_),
    .B2(_08366_),
    .A2(_10359_),
    .A1(\cpu.ex.r_14[2] ));
 sg13g2_buf_1 _17152_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10363_));
 sg13g2_nor2b_1 _17153_ (.A(net1002),
    .B_N(net871),
    .Y(_10364_));
 sg13g2_buf_2 _17154_ (.A(_10364_),
    .X(_10365_));
 sg13g2_nand3_1 _17155_ (.B(_10363_),
    .C(_10365_),
    .A(net744),
    .Y(_10366_));
 sg13g2_o21ai_1 _17156_ (.B1(_10366_),
    .Y(_10367_),
    .A1(_10245_),
    .A2(_10362_));
 sg13g2_nand2_1 _17157_ (.Y(_10368_),
    .A(_10275_),
    .B(_10367_));
 sg13g2_nor2b_1 _17158_ (.A(_10233_),
    .B_N(_10236_),
    .Y(_10369_));
 sg13g2_buf_2 _17159_ (.A(_10369_),
    .X(_10370_));
 sg13g2_a22oi_1 _17160_ (.Y(_10371_),
    .B1(_10370_),
    .B2(\cpu.ex.r_lr[2] ),
    .A2(net748),
    .A1(\cpu.ex.r_8[2] ));
 sg13g2_nor2_1 _17161_ (.A(_10191_),
    .B(net1091),
    .Y(_10372_));
 sg13g2_buf_2 _17162_ (.A(_10372_),
    .X(_10373_));
 sg13g2_nor2b_1 _17163_ (.A(_10371_),
    .B_N(_10373_),
    .Y(_10374_));
 sg13g2_nand2_1 _17164_ (.Y(_10375_),
    .A(_10190_),
    .B(_10191_));
 sg13g2_buf_2 _17165_ (.A(_10375_),
    .X(_10376_));
 sg13g2_nor2b_1 _17166_ (.A(net1000),
    .B_N(net872),
    .Y(_10377_));
 sg13g2_buf_2 _17167_ (.A(_10377_),
    .X(_10378_));
 sg13g2_a22oi_1 _17168_ (.Y(_10379_),
    .B1(_10378_),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10199_),
    .A1(\cpu.ex.r_epc[2] ));
 sg13g2_nor2_1 _17169_ (.A(_10376_),
    .B(_10379_),
    .Y(_10380_));
 sg13g2_nand2_1 _17170_ (.Y(_10381_),
    .A(net741),
    .B(net745));
 sg13g2_nor2b_1 _17171_ (.A(_10196_),
    .B_N(_10192_),
    .Y(_10382_));
 sg13g2_buf_1 _17172_ (.A(_10382_),
    .X(_10383_));
 sg13g2_a22oi_1 _17173_ (.Y(_10384_),
    .B1(_10383_),
    .B2(\cpu.ex.r_stmp[2] ),
    .A2(_10311_),
    .A1(\cpu.ex.r_12[2] ));
 sg13g2_nor2_1 _17174_ (.A(_10381_),
    .B(_10384_),
    .Y(_10385_));
 sg13g2_buf_1 _17175_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10386_));
 sg13g2_a22oi_1 _17176_ (.Y(_10387_),
    .B1(_10303_),
    .B2(\cpu.ex.r_mult[18] ),
    .A2(_10301_),
    .A1(_10386_));
 sg13g2_buf_1 _17177_ (.A(_10383_),
    .X(_10388_));
 sg13g2_nor2b_1 _17178_ (.A(_10387_),
    .B_N(net653),
    .Y(_10389_));
 sg13g2_nor4_1 _17179_ (.A(_10374_),
    .B(_10380_),
    .C(_10385_),
    .D(_10389_),
    .Y(_10390_));
 sg13g2_nand4_1 _17180_ (.B(_10360_),
    .C(_10368_),
    .A(net540),
    .Y(_10391_),
    .D(_10390_));
 sg13g2_buf_1 _17181_ (.A(_10391_),
    .X(_10392_));
 sg13g2_nand3_1 _17182_ (.B(_10354_),
    .C(_10392_),
    .A(_10353_),
    .Y(_10393_));
 sg13g2_buf_1 _17183_ (.A(_00297_),
    .X(_10394_));
 sg13g2_nand2b_1 _17184_ (.Y(_10395_),
    .B(_10353_),
    .A_N(_10394_));
 sg13g2_mux2_1 _17185_ (.A0(_10393_),
    .A1(_10395_),
    .S(_10205_),
    .X(_10396_));
 sg13g2_nand4_1 _17186_ (.B(_10210_),
    .C(_10352_),
    .A(_10184_),
    .Y(_10397_),
    .D(_10396_));
 sg13g2_buf_2 _17187_ (.A(_00294_),
    .X(_10398_));
 sg13g2_buf_2 _17188_ (.A(_00296_),
    .X(_10399_));
 sg13g2_mux2_1 _17189_ (.A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_10[7] ),
    .S(net740),
    .X(_10400_));
 sg13g2_nand2_1 _17190_ (.Y(_10401_),
    .A(net750),
    .B(\cpu.ex.r_9[7] ));
 sg13g2_nand2_1 _17191_ (.Y(_10402_),
    .A(_10294_),
    .B(_10228_));
 sg13g2_a21oi_1 _17192_ (.A1(net658),
    .A2(_10401_),
    .Y(_10403_),
    .B1(_10402_));
 sg13g2_o21ai_1 _17193_ (.B1(_10403_),
    .Y(_10404_),
    .A1(net658),
    .A2(_10400_));
 sg13g2_mux2_1 _17194_ (.A0(\cpu.ex.r_lr[7] ),
    .A1(\cpu.ex.r_epc[7] ),
    .S(net740),
    .X(_10405_));
 sg13g2_buf_1 _17195_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10406_));
 sg13g2_a21oi_1 _17196_ (.A1(_10259_),
    .A2(_10406_),
    .Y(_10407_),
    .B1(net658));
 sg13g2_nor2b_1 _17197_ (.A(_10407_),
    .B_N(net659),
    .Y(_10408_));
 sg13g2_o21ai_1 _17198_ (.B1(_10408_),
    .Y(_10409_),
    .A1(net741),
    .A2(_10405_));
 sg13g2_nand3_1 _17199_ (.B(_10404_),
    .C(_10409_),
    .A(net540),
    .Y(_10410_));
 sg13g2_nand2b_1 _17200_ (.Y(_10411_),
    .B(net743),
    .A_N(_00265_));
 sg13g2_nand2_1 _17201_ (.Y(_10412_),
    .A(net750),
    .B(\cpu.ex.r_13[7] ));
 sg13g2_nand2_1 _17202_ (.Y(_10413_),
    .A(net746),
    .B(net747));
 sg13g2_a21oi_1 _17203_ (.A1(_10411_),
    .A2(_10412_),
    .Y(_10414_),
    .B1(_10413_));
 sg13g2_nor2_1 _17204_ (.A(net746),
    .B(net739),
    .Y(_10415_));
 sg13g2_buf_1 _17205_ (.A(\cpu.dec.user_io ),
    .X(_10416_));
 sg13g2_mux2_1 _17206_ (.A0(_10416_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net869),
    .X(_10417_));
 sg13g2_and2_1 _17207_ (.A(_10415_),
    .B(_10417_),
    .X(_10418_));
 sg13g2_o21ai_1 _17208_ (.B1(net656),
    .Y(_10419_),
    .A1(_10414_),
    .A2(_10418_));
 sg13g2_buf_1 _17209_ (.A(_10311_),
    .X(_10420_));
 sg13g2_nand3_1 _17210_ (.B(_10257_),
    .C(net652),
    .A(\cpu.ex.r_12[7] ),
    .Y(_10421_));
 sg13g2_nand3_1 _17211_ (.B(net655),
    .C(_10378_),
    .A(\cpu.ex.r_11[7] ),
    .Y(_10422_));
 sg13g2_a22oi_1 _17212_ (.Y(_10423_),
    .B1(_10370_),
    .B2(\cpu.ex.r_mult[23] ),
    .A2(net748),
    .A1(\cpu.ex.r_14[7] ));
 sg13g2_and2_1 _17213_ (.A(net1002),
    .B(net1000),
    .X(_10424_));
 sg13g2_buf_2 _17214_ (.A(_10424_),
    .X(_10425_));
 sg13g2_nand2b_1 _17215_ (.Y(_10426_),
    .B(_10425_),
    .A_N(_10423_));
 sg13g2_nand4_1 _17216_ (.B(_10421_),
    .C(_10422_),
    .A(_10419_),
    .Y(_10427_),
    .D(_10426_));
 sg13g2_nand2b_1 _17217_ (.Y(_10428_),
    .B(net607),
    .A_N(_09013_));
 sg13g2_o21ai_1 _17218_ (.B1(_10428_),
    .Y(_10429_),
    .A1(_10410_),
    .A2(_10427_));
 sg13g2_buf_1 _17219_ (.A(_10429_),
    .X(_10430_));
 sg13g2_inv_2 _17220_ (.Y(_10431_),
    .A(_09818_));
 sg13g2_a22oi_1 _17221_ (.Y(_10432_),
    .B1(net653),
    .B2(\cpu.ex.r_mult[21] ),
    .A2(net652),
    .A1(\cpu.ex.r_13[5] ));
 sg13g2_inv_1 _17222_ (.Y(_10433_),
    .A(_10432_));
 sg13g2_inv_1 _17223_ (.Y(_10434_),
    .A(_00263_));
 sg13g2_nand2_1 _17224_ (.Y(_10435_),
    .A(net742),
    .B(_10434_));
 sg13g2_nand3_1 _17225_ (.B(\cpu.ex.r_lr[5] ),
    .C(net659),
    .A(net750),
    .Y(_10436_));
 sg13g2_o21ai_1 _17226_ (.B1(_10436_),
    .Y(_10437_),
    .A1(_10299_),
    .A2(_10435_));
 sg13g2_mux2_1 _17227_ (.A0(\cpu.ex.r_8[5] ),
    .A1(\cpu.ex.r_9[5] ),
    .S(net871),
    .X(_10438_));
 sg13g2_a22oi_1 _17228_ (.Y(_10439_),
    .B1(_10438_),
    .B2(net750),
    .A2(net654),
    .A1(\cpu.ex.r_10[5] ));
 sg13g2_and2_1 _17229_ (.A(net1001),
    .B(net1000),
    .X(_10440_));
 sg13g2_buf_2 _17230_ (.A(_10440_),
    .X(_10441_));
 sg13g2_nand3_1 _17231_ (.B(_10441_),
    .C(net654),
    .A(\cpu.ex.r_14[5] ),
    .Y(_10442_));
 sg13g2_o21ai_1 _17232_ (.B1(_10442_),
    .Y(_10443_),
    .A1(_10402_),
    .A2(_10439_));
 sg13g2_a221oi_1 _17233_ (.B2(net658),
    .C1(_10443_),
    .B1(_10437_),
    .A1(_10303_),
    .Y(_10444_),
    .A2(_10433_));
 sg13g2_nand4_1 _17234_ (.B(net656),
    .C(\cpu.ex.r_12[5] ),
    .A(_10235_),
    .Y(_10445_),
    .D(_10194_));
 sg13g2_nor2_1 _17235_ (.A(net745),
    .B(_10376_),
    .Y(_10446_));
 sg13g2_nand3_1 _17236_ (.B(\cpu.ex.r_11[5] ),
    .C(_10446_),
    .A(net660),
    .Y(_10447_));
 sg13g2_buf_1 _17237_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10448_));
 sg13g2_and2_1 _17238_ (.A(net870),
    .B(\cpu.ex.r_stmp[5] ),
    .X(_10449_));
 sg13g2_a21oi_1 _17239_ (.A1(_10229_),
    .A2(_10448_),
    .Y(_10450_),
    .B1(_10449_));
 sg13g2_nor2b_1 _17240_ (.A(net738),
    .B_N(\cpu.ex.r_epc[5] ),
    .Y(_10451_));
 sg13g2_o21ai_1 _17241_ (.B1(_10383_),
    .Y(_10452_),
    .A1(_10269_),
    .A2(_10451_));
 sg13g2_a21o_1 _17242_ (.A2(_10450_),
    .A1(net741),
    .B1(_10452_),
    .X(_10453_));
 sg13g2_and4_1 _17243_ (.A(_10219_),
    .B(_10445_),
    .C(_10447_),
    .D(_10453_),
    .X(_10454_));
 sg13g2_a22oi_1 _17244_ (.Y(_10455_),
    .B1(_10444_),
    .B2(_10454_),
    .A2(net607),
    .A1(_10431_));
 sg13g2_buf_1 _17245_ (.A(_10455_),
    .X(_10456_));
 sg13g2_inv_1 _17246_ (.Y(_10457_),
    .A(_10456_));
 sg13g2_mux4_1 _17247_ (.S0(_10179_),
    .A0(_10398_),
    .A1(_10399_),
    .A2(_10430_),
    .A3(_10457_),
    .S1(_10351_),
    .X(_10458_));
 sg13g2_nand2_1 _17248_ (.Y(_10459_),
    .A(net495),
    .B(_10458_));
 sg13g2_a21o_1 _17249_ (.A2(_09024_),
    .A1(_08781_),
    .B1(_09025_),
    .X(_10460_));
 sg13g2_nand2_1 _17250_ (.Y(_10461_),
    .A(net891),
    .B(_10224_));
 sg13g2_buf_1 _17251_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10462_));
 sg13g2_mux2_1 _17252_ (.A0(_10462_),
    .A1(\cpu.ex.r_stmp[4] ),
    .S(net1091),
    .X(_10463_));
 sg13g2_a22oi_1 _17253_ (.Y(_10464_),
    .B1(_10463_),
    .B2(_10269_),
    .A2(_10303_),
    .A1(\cpu.ex.r_mult[20] ));
 sg13g2_nand2b_1 _17254_ (.Y(_10465_),
    .B(_10383_),
    .A_N(_10464_));
 sg13g2_nand2b_1 _17255_ (.Y(_10466_),
    .B(_10227_),
    .A_N(_00262_));
 sg13g2_nand2b_1 _17256_ (.Y(_10467_),
    .B(\cpu.ex.r_11[4] ),
    .A_N(net1000));
 sg13g2_nand3_1 _17257_ (.B(_10466_),
    .C(_10467_),
    .A(net1001),
    .Y(_10468_));
 sg13g2_nand2b_1 _17258_ (.Y(_10469_),
    .B(\cpu.ex.r_epc[4] ),
    .A_N(net1091));
 sg13g2_a21oi_1 _17259_ (.A1(_10254_),
    .A2(_10469_),
    .Y(_10470_),
    .B1(_10376_));
 sg13g2_and2_1 _17260_ (.A(_10225_),
    .B(_10329_),
    .X(_10471_));
 sg13g2_nor2_1 _17261_ (.A(_08736_),
    .B(net1003),
    .Y(_10472_));
 sg13g2_and4_1 _17262_ (.A(_10269_),
    .B(_10228_),
    .C(\cpu.ex.r_10[4] ),
    .D(_10359_),
    .X(_10473_));
 sg13g2_a221oi_1 _17263_ (.B2(_10472_),
    .C1(_10473_),
    .B1(_10471_),
    .A1(_10468_),
    .Y(_10474_),
    .A2(_10470_));
 sg13g2_nand2_1 _17264_ (.Y(_10475_),
    .A(net1001),
    .B(\cpu.ex.r_9[4] ));
 sg13g2_nand2b_1 _17265_ (.Y(_10476_),
    .B(\cpu.ex.r_lr[4] ),
    .A_N(net1001));
 sg13g2_nand3_1 _17266_ (.B(_10475_),
    .C(_10476_),
    .A(net1003),
    .Y(_10477_));
 sg13g2_a21oi_1 _17267_ (.A1(net1001),
    .A2(\cpu.ex.r_8[4] ),
    .Y(_10478_),
    .B1(net1003));
 sg13g2_nor2b_1 _17268_ (.A(_10478_),
    .B_N(_10373_),
    .Y(_10479_));
 sg13g2_mux2_1 _17269_ (.A0(\cpu.ex.r_12[4] ),
    .A1(\cpu.ex.r_13[4] ),
    .S(net1003),
    .X(_10480_));
 sg13g2_and3_1 _17270_ (.X(_10481_),
    .A(net1000),
    .B(_10311_),
    .C(_10480_));
 sg13g2_a221oi_1 _17271_ (.B2(_10479_),
    .C1(_10481_),
    .B1(_10477_),
    .A1(\cpu.ex.r_14[4] ),
    .Y(_10482_),
    .A2(_10334_));
 sg13g2_nand4_1 _17272_ (.B(_10465_),
    .C(_10474_),
    .A(_10219_),
    .Y(_10483_),
    .D(_10482_));
 sg13g2_buf_1 _17273_ (.A(_10483_),
    .X(_10484_));
 sg13g2_nand4_1 _17274_ (.B(_10202_),
    .C(_10461_),
    .A(_09023_),
    .Y(_10485_),
    .D(_10484_));
 sg13g2_nand3_1 _17275_ (.B(_10461_),
    .C(_10484_),
    .A(_10203_),
    .Y(_10486_));
 sg13g2_o21ai_1 _17276_ (.B1(_10486_),
    .Y(_10487_),
    .A1(_10460_),
    .A2(_10485_));
 sg13g2_buf_1 _17277_ (.A(_10487_),
    .X(_10488_));
 sg13g2_nand2b_1 _17278_ (.Y(_10489_),
    .B(_10176_),
    .A_N(_08144_));
 sg13g2_a21oi_2 _17279_ (.B1(_10489_),
    .Y(_10490_),
    .A2(_10202_),
    .A1(net379));
 sg13g2_nor2_1 _17280_ (.A(_10488_),
    .B(_10490_),
    .Y(_10491_));
 sg13g2_buf_2 _17281_ (.A(_10491_),
    .X(_10492_));
 sg13g2_inv_1 _17282_ (.Y(_10493_),
    .A(_00264_));
 sg13g2_a22oi_1 _17283_ (.Y(_10494_),
    .B1(_10415_),
    .B2(\cpu.ex.r_stmp[6] ),
    .A2(_10251_),
    .A1(_10493_));
 sg13g2_nand2b_1 _17284_ (.Y(_10495_),
    .B(_10425_),
    .A_N(_10494_));
 sg13g2_and2_1 _17285_ (.A(_10234_),
    .B(\cpu.ex.r_14[6] ),
    .X(_10496_));
 sg13g2_nor2_1 _17286_ (.A(net745),
    .B(_10337_),
    .Y(_10497_));
 sg13g2_and2_1 _17287_ (.A(net747),
    .B(\cpu.ex.r_9[6] ),
    .X(_10498_));
 sg13g2_a22oi_1 _17288_ (.Y(_10499_),
    .B1(_10497_),
    .B2(_10498_),
    .A2(_10496_),
    .A1(_10274_));
 sg13g2_nand3_1 _17289_ (.B(\cpu.ex.r_10[6] ),
    .C(net748),
    .A(_10228_),
    .Y(_10500_));
 sg13g2_buf_2 _17290_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10501_));
 sg13g2_nand3_1 _17291_ (.B(_10501_),
    .C(_10303_),
    .A(_10254_),
    .Y(_10502_));
 sg13g2_a21oi_1 _17292_ (.A1(_10500_),
    .A2(_10502_),
    .Y(_10503_),
    .B1(net750));
 sg13g2_a22oi_1 _17293_ (.Y(_10504_),
    .B1(net655),
    .B2(\cpu.ex.r_11[6] ),
    .A2(_10194_),
    .A1(\cpu.ex.r_8[6] ));
 sg13g2_nor2_1 _17294_ (.A(_10402_),
    .B(_10504_),
    .Y(_10505_));
 sg13g2_mux2_1 _17295_ (.A0(\cpu.ex.r_lr[6] ),
    .A1(\cpu.ex.r_epc[6] ),
    .S(_10258_),
    .X(_10506_));
 sg13g2_nand3_1 _17296_ (.B(_10199_),
    .C(_10506_),
    .A(_10237_),
    .Y(_10507_));
 sg13g2_nand3_1 _17297_ (.B(_10441_),
    .C(_10365_),
    .A(\cpu.ex.r_13[6] ),
    .Y(_10508_));
 sg13g2_nand2_1 _17298_ (.Y(_10509_),
    .A(_10507_),
    .B(_10508_));
 sg13g2_nand3_1 _17299_ (.B(\cpu.ex.r_12[6] ),
    .C(_10441_),
    .A(_10269_),
    .Y(_10510_));
 sg13g2_buf_1 _17300_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10511_));
 sg13g2_nand4_1 _17301_ (.B(_10258_),
    .C(_10511_),
    .A(_10269_),
    .Y(_10512_),
    .D(_10199_));
 sg13g2_o21ai_1 _17302_ (.B1(_10512_),
    .Y(_10513_),
    .A1(_10259_),
    .A2(_10510_));
 sg13g2_nor4_1 _17303_ (.A(_10503_),
    .B(_10505_),
    .C(_10509_),
    .D(_10513_),
    .Y(_10514_));
 sg13g2_nand4_1 _17304_ (.B(_10495_),
    .C(_10499_),
    .A(net540),
    .Y(_10515_),
    .D(_10514_));
 sg13g2_o21ai_1 _17305_ (.B1(_10515_),
    .Y(_10516_),
    .A1(_09010_),
    .A2(net540));
 sg13g2_mux2_1 _17306_ (.A0(_00295_),
    .A1(_10516_),
    .S(_10351_),
    .X(_10517_));
 sg13g2_buf_8 _17307_ (.A(_10517_),
    .X(_10518_));
 sg13g2_a221oi_1 _17308_ (.B2(_10353_),
    .C1(_10175_),
    .B1(net247),
    .A1(_10180_),
    .Y(_10519_),
    .A2(_10492_));
 sg13g2_xor2_1 _17309_ (.B(_10172_),
    .A(\cpu.ex.r_mult_off[3] ),
    .X(_10520_));
 sg13g2_and2_1 _17310_ (.A(_09207_),
    .B(_10520_),
    .X(_10521_));
 sg13g2_buf_1 _17311_ (.A(_10521_),
    .X(_10522_));
 sg13g2_inv_1 _17312_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(_10522_));
 sg13g2_a221oi_1 _17313_ (.B2(_10519_),
    .C1(\cpu.ex.c_mult_off[3] ),
    .B1(_10459_),
    .A1(_10175_),
    .Y(_10523_),
    .A2(_10397_));
 sg13g2_buf_1 _17314_ (.A(_10523_),
    .X(_10524_));
 sg13g2_buf_1 _17315_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10525_));
 sg13g2_nand3_1 _17316_ (.B(_10525_),
    .C(_10365_),
    .A(net742),
    .Y(_10526_));
 sg13g2_buf_1 _17317_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10527_));
 sg13g2_nand3_1 _17318_ (.B(_10527_),
    .C(net654),
    .A(net657),
    .Y(_10528_));
 sg13g2_a21oi_1 _17319_ (.A1(_10526_),
    .A2(_10528_),
    .Y(_10529_),
    .B1(net660));
 sg13g2_nand3_1 _17320_ (.B(\cpu.ex.r_12[12] ),
    .C(_10194_),
    .A(net742),
    .Y(_10530_));
 sg13g2_nand3_1 _17321_ (.B(\cpu.ex.r_11[12] ),
    .C(net655),
    .A(net657),
    .Y(_10531_));
 sg13g2_a21oi_1 _17322_ (.A1(_10530_),
    .A2(_10531_),
    .Y(_10532_),
    .B1(net744));
 sg13g2_mux2_1 _17323_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_9[12] ),
    .S(net739),
    .X(_10533_));
 sg13g2_nand3_1 _17324_ (.B(_10365_),
    .C(_10533_),
    .A(net657),
    .Y(_10534_));
 sg13g2_nand3_1 _17325_ (.B(_10194_),
    .C(_10378_),
    .A(\cpu.ex.r_8[12] ),
    .Y(_10535_));
 sg13g2_nand2_1 _17326_ (.Y(_10536_),
    .A(_10534_),
    .B(_10535_));
 sg13g2_a22oi_1 _17327_ (.Y(_10537_),
    .B1(_10365_),
    .B2(\cpu.ex.r_13[12] ),
    .A2(net654),
    .A1(\cpu.ex.r_14[12] ));
 sg13g2_nor2_1 _17328_ (.A(_10333_),
    .B(_10537_),
    .Y(_10538_));
 sg13g2_nor4_1 _17329_ (.A(_10529_),
    .B(_10532_),
    .C(_10536_),
    .D(_10538_),
    .Y(_10539_));
 sg13g2_a22oi_1 _17330_ (.Y(_10540_),
    .B1(_10378_),
    .B2(\cpu.ex.r_10[12] ),
    .A2(_10329_),
    .A1(\cpu.ex.r_stmp[12] ));
 sg13g2_inv_1 _17331_ (.Y(_10541_),
    .A(_00270_));
 sg13g2_mux2_1 _17332_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(\cpu.ex.r_mult[28] ),
    .S(net738),
    .X(_10542_));
 sg13g2_a221oi_1 _17333_ (.B2(net744),
    .C1(net741),
    .B1(_10542_),
    .A1(_10541_),
    .Y(_10543_),
    .A2(_10441_));
 sg13g2_a21oi_1 _17334_ (.A1(net741),
    .A2(_10540_),
    .Y(_10544_),
    .B1(_10543_));
 sg13g2_a21oi_1 _17335_ (.A1(net740),
    .A2(_10544_),
    .Y(_10545_),
    .B1(net607));
 sg13g2_a22oi_1 _17336_ (.Y(_10546_),
    .B1(_10539_),
    .B2(_10545_),
    .A2(net607),
    .A1(_08822_));
 sg13g2_inv_1 _17337_ (.Y(_10547_),
    .A(_10546_));
 sg13g2_nor2_1 _17338_ (.A(net747),
    .B(_10263_),
    .Y(_10548_));
 sg13g2_a22oi_1 _17339_ (.Y(_10549_),
    .B1(_10548_),
    .B2(\cpu.ex.r_stmp[14] ),
    .A2(_10338_),
    .A1(\cpu.ex.r_13[14] ));
 sg13g2_nor2_1 _17340_ (.A(net739),
    .B(_10337_),
    .Y(_10550_));
 sg13g2_and2_1 _17341_ (.A(net739),
    .B(\cpu.ex.r_10[14] ),
    .X(_10551_));
 sg13g2_a221oi_1 _17342_ (.B2(net654),
    .C1(net742),
    .B1(_10551_),
    .A1(\cpu.ex.r_lr[14] ),
    .Y(_10552_),
    .A2(_10550_));
 sg13g2_a21oi_1 _17343_ (.A1(net656),
    .A2(_10549_),
    .Y(_10553_),
    .B1(_10552_));
 sg13g2_buf_1 _17344_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10554_));
 sg13g2_a22oi_1 _17345_ (.Y(_10555_),
    .B1(_10303_),
    .B2(\cpu.ex.r_mult[30] ),
    .A2(_10301_),
    .A1(_10554_));
 sg13g2_nand2b_1 _17346_ (.Y(_10556_),
    .B(net653),
    .A_N(_10555_));
 sg13g2_inv_1 _17347_ (.Y(_10557_),
    .A(_00272_));
 sg13g2_a22oi_1 _17348_ (.Y(_10558_),
    .B1(_10441_),
    .B2(_10557_),
    .A2(_10199_),
    .A1(\cpu.ex.r_epc[14] ));
 sg13g2_nand2b_1 _17349_ (.Y(_10559_),
    .B(net655),
    .A_N(_10558_));
 sg13g2_inv_1 _17350_ (.Y(_10560_),
    .A(\cpu.ex.r_8[14] ));
 sg13g2_nand2_1 _17351_ (.Y(_10561_),
    .A(net738),
    .B(\cpu.ex.r_12[14] ));
 sg13g2_o21ai_1 _17352_ (.B1(_10561_),
    .Y(_10562_),
    .A1(net738),
    .A2(_10560_));
 sg13g2_nand3_1 _17353_ (.B(_10194_),
    .C(_10562_),
    .A(net747),
    .Y(_10563_));
 sg13g2_nand3_1 _17354_ (.B(_10559_),
    .C(_10563_),
    .A(_10556_),
    .Y(_10564_));
 sg13g2_a22oi_1 _17355_ (.Y(_10565_),
    .B1(_10497_),
    .B2(\cpu.ex.r_9[14] ),
    .A2(_10274_),
    .A1(\cpu.ex.r_14[14] ));
 sg13g2_buf_2 _17356_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10566_));
 sg13g2_nand3_1 _17357_ (.B(_10566_),
    .C(_10329_),
    .A(net750),
    .Y(_10567_));
 sg13g2_nand3_1 _17358_ (.B(\cpu.ex.r_11[14] ),
    .C(_10359_),
    .A(net749),
    .Y(_10568_));
 sg13g2_a21o_1 _17359_ (.A2(_10568_),
    .A1(_10567_),
    .B1(net741),
    .X(_10569_));
 sg13g2_o21ai_1 _17360_ (.B1(_10569_),
    .Y(_10570_),
    .A1(net744),
    .A2(_10565_));
 sg13g2_or4_1 _17361_ (.A(net607),
    .B(_10553_),
    .C(_10564_),
    .D(_10570_),
    .X(_10571_));
 sg13g2_o21ai_1 _17362_ (.B1(_10571_),
    .Y(_10572_),
    .A1(net774),
    .A2(net491));
 sg13g2_buf_1 _17363_ (.A(_10572_),
    .X(_10573_));
 sg13g2_nor2b_1 _17364_ (.A(_00271_),
    .B_N(net738),
    .Y(_10574_));
 sg13g2_nor2b_1 _17365_ (.A(net745),
    .B_N(\cpu.ex.r_11[13] ),
    .Y(_10575_));
 sg13g2_o21ai_1 _17366_ (.B1(net747),
    .Y(_10576_),
    .A1(_10574_),
    .A2(_10575_));
 sg13g2_nand2_1 _17367_ (.Y(_10577_),
    .A(\cpu.ex.r_epc[13] ),
    .B(net659));
 sg13g2_a21oi_1 _17368_ (.A1(_10576_),
    .A2(_10577_),
    .Y(_10578_),
    .B1(_10376_));
 sg13g2_buf_1 _17369_ (.A(\cpu.ex.r_sp[13] ),
    .X(_10579_));
 sg13g2_nand3_1 _17370_ (.B(_10579_),
    .C(net654),
    .A(net744),
    .Y(_10580_));
 sg13g2_nand3_1 _17371_ (.B(\cpu.ex.r_9[13] ),
    .C(net652),
    .A(net658),
    .Y(_10581_));
 sg13g2_a21oi_1 _17372_ (.A1(_10580_),
    .A2(_10581_),
    .Y(_10582_),
    .B1(net656));
 sg13g2_nand3_1 _17373_ (.B(_10441_),
    .C(_10365_),
    .A(\cpu.ex.r_13[13] ),
    .Y(_10583_));
 sg13g2_nand3b_1 _17374_ (.B(net739),
    .C(\cpu.ex.r_14[13] ),
    .Y(_10584_),
    .A_N(net746));
 sg13g2_buf_2 _17375_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10585_));
 sg13g2_nand3b_1 _17376_ (.B(_10585_),
    .C(net746),
    .Y(_10586_),
    .A_N(net739));
 sg13g2_nand2_1 _17377_ (.Y(_10587_),
    .A(net743),
    .B(_10239_));
 sg13g2_a21o_1 _17378_ (.A2(_10586_),
    .A1(_10584_),
    .B1(_10587_),
    .X(_10588_));
 sg13g2_nand3b_1 _17379_ (.B(\cpu.ex.r_10[13] ),
    .C(net739),
    .Y(_10589_),
    .A_N(net738));
 sg13g2_nand3b_1 _17380_ (.B(net738),
    .C(\cpu.ex.r_stmp[13] ),
    .Y(_10590_),
    .A_N(net739));
 sg13g2_a21o_1 _17381_ (.A2(_10590_),
    .A1(_10589_),
    .B1(_10263_),
    .X(_10591_));
 sg13g2_nand3_1 _17382_ (.B(_10588_),
    .C(_10591_),
    .A(_10583_),
    .Y(_10592_));
 sg13g2_a221oi_1 _17383_ (.B2(\cpu.ex.r_lr[13] ),
    .C1(net742),
    .B1(_10370_),
    .A1(\cpu.ex.r_8[13] ),
    .Y(_10593_),
    .A2(net748));
 sg13g2_buf_2 _17384_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10594_));
 sg13g2_a221oi_1 _17385_ (.B2(_10594_),
    .C1(net657),
    .B1(_10370_),
    .A1(\cpu.ex.r_12[13] ),
    .Y(_10595_),
    .A2(net748));
 sg13g2_nor3_1 _17386_ (.A(net740),
    .B(_10593_),
    .C(_10595_),
    .Y(_10596_));
 sg13g2_nor4_1 _17387_ (.A(_10578_),
    .B(_10582_),
    .C(_10592_),
    .D(_10596_),
    .Y(_10597_));
 sg13g2_nor2_1 _17388_ (.A(net676),
    .B(net540),
    .Y(_10598_));
 sg13g2_a21oi_1 _17389_ (.A1(net491),
    .A2(_10597_),
    .Y(_10599_),
    .B1(_10598_));
 sg13g2_inv_1 _17390_ (.Y(_10600_),
    .A(_10599_));
 sg13g2_nor2_1 _17391_ (.A(_09457_),
    .B(_10221_),
    .Y(_10601_));
 sg13g2_buf_1 _17392_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10602_));
 sg13g2_nand3_1 _17393_ (.B(_10602_),
    .C(net653),
    .A(net657),
    .Y(_10603_));
 sg13g2_nand3_1 _17394_ (.B(\cpu.ex.r_12[15] ),
    .C(net652),
    .A(net742),
    .Y(_10604_));
 sg13g2_nand2_1 _17395_ (.Y(_10605_),
    .A(_10603_),
    .B(_10604_));
 sg13g2_a22oi_1 _17396_ (.Y(_10606_),
    .B1(_10425_),
    .B2(\cpu.ex.r_14[15] ),
    .A2(_10373_),
    .A1(\cpu.ex.r_8[15] ));
 sg13g2_nor2_1 _17397_ (.A(net744),
    .B(_10606_),
    .Y(_10607_));
 sg13g2_o21ai_1 _17398_ (.B1(net741),
    .Y(_10608_),
    .A1(_10605_),
    .A2(_10607_));
 sg13g2_mux2_1 _17399_ (.A0(\cpu.ex.r_lr[15] ),
    .A1(\cpu.ex.r_9[15] ),
    .S(net747),
    .X(_10609_));
 sg13g2_mux2_1 _17400_ (.A0(\cpu.ex.r_epc[15] ),
    .A1(\cpu.ex.r_11[15] ),
    .S(net660),
    .X(_10610_));
 sg13g2_a22oi_1 _17401_ (.Y(_10611_),
    .B1(_10378_),
    .B2(\cpu.ex.r_10[15] ),
    .A2(_10329_),
    .A1(\cpu.ex.r_stmp[15] ));
 sg13g2_nor2_1 _17402_ (.A(_10263_),
    .B(_10611_),
    .Y(_10612_));
 sg13g2_a221oi_1 _17403_ (.B2(_10446_),
    .C1(_10612_),
    .B1(_10610_),
    .A1(_10497_),
    .Y(_10613_),
    .A2(_10609_));
 sg13g2_buf_1 _17404_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10614_));
 sg13g2_a22oi_1 _17405_ (.Y(_10615_),
    .B1(_10361_),
    .B2(_10614_),
    .A2(_10359_),
    .A1(\cpu.ex.r_15[15] ));
 sg13g2_a22oi_1 _17406_ (.Y(_10616_),
    .B1(net653),
    .B2(\cpu.ex.r_mult[31] ),
    .A2(net652),
    .A1(\cpu.ex.r_13[15] ));
 sg13g2_a21o_1 _17407_ (.A2(_10616_),
    .A1(_10615_),
    .B1(_10240_),
    .X(_10617_));
 sg13g2_nand4_1 _17408_ (.B(_10608_),
    .C(_10613_),
    .A(net491),
    .Y(_10618_),
    .D(_10617_));
 sg13g2_nand2b_1 _17409_ (.Y(_10619_),
    .B(_10618_),
    .A_N(_10601_));
 sg13g2_mux4_1 _17410_ (.S0(\cpu.ex.c_mult_off[1] ),
    .A0(_10547_),
    .A1(_10573_),
    .A2(_10600_),
    .A3(_10619_),
    .S1(net495),
    .X(_10620_));
 sg13g2_buf_1 _17411_ (.A(_00195_),
    .X(_10621_));
 sg13g2_mux4_1 _17412_ (.S0(_10179_),
    .A0(_10621_),
    .A1(_00289_),
    .A2(_00194_),
    .A3(_00196_),
    .S1(\cpu.ex.c_mult_off[0] ),
    .X(_10622_));
 sg13g2_inv_1 _17413_ (.Y(_10623_),
    .A(_10622_));
 sg13g2_a21oi_1 _17414_ (.A1(_10205_),
    .A2(_10623_),
    .Y(_10624_),
    .B1(_10175_));
 sg13g2_o21ai_1 _17415_ (.B1(_10624_),
    .Y(_10625_),
    .A1(_10205_),
    .A2(_10620_));
 sg13g2_buf_2 _17416_ (.A(_00292_),
    .X(_10626_));
 sg13g2_buf_2 _17417_ (.A(\cpu.addr[9] ),
    .X(_10627_));
 sg13g2_inv_1 _17418_ (.Y(_10628_),
    .A(\cpu.ex.r_9[9] ));
 sg13g2_buf_1 _17419_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10629_));
 sg13g2_nand3_1 _17420_ (.B(_10629_),
    .C(_10320_),
    .A(_10255_),
    .Y(_10630_));
 sg13g2_o21ai_1 _17421_ (.B1(_10630_),
    .Y(_10631_),
    .A1(_10628_),
    .A2(_10317_));
 sg13g2_nand3_1 _17422_ (.B(\cpu.ex.r_11[9] ),
    .C(_10251_),
    .A(_10229_),
    .Y(_10632_));
 sg13g2_nand3_1 _17423_ (.B(\cpu.ex.r_stmp[9] ),
    .C(_10329_),
    .A(_10270_),
    .Y(_10633_));
 sg13g2_nand2_1 _17424_ (.Y(_10634_),
    .A(_10632_),
    .B(_10633_));
 sg13g2_a22oi_1 _17425_ (.Y(_10635_),
    .B1(_10634_),
    .B2(net740),
    .A2(_10631_),
    .A1(_10248_));
 sg13g2_nor2_1 _17426_ (.A(_10333_),
    .B(_10337_),
    .Y(_10636_));
 sg13g2_and2_1 _17427_ (.A(net659),
    .B(net655),
    .X(_10637_));
 sg13g2_nor3_1 _17428_ (.A(_00267_),
    .B(_10333_),
    .C(_10376_),
    .Y(_10638_));
 sg13g2_a221oi_1 _17429_ (.B2(\cpu.ex.r_epc[9] ),
    .C1(_10638_),
    .B1(_10637_),
    .A1(\cpu.ex.r_13[9] ),
    .Y(_10639_),
    .A2(_10636_));
 sg13g2_a22oi_1 _17430_ (.Y(_10640_),
    .B1(_10425_),
    .B2(\cpu.ex.r_mult[25] ),
    .A2(_10373_),
    .A1(\cpu.ex.r_lr[9] ));
 sg13g2_inv_1 _17431_ (.Y(_10641_),
    .A(_10640_));
 sg13g2_mux4_1 _17432_ (.S0(net743),
    .A0(\cpu.ex.r_8[9] ),
    .A1(\cpu.ex.r_10[9] ),
    .A2(\cpu.ex.r_12[9] ),
    .A3(\cpu.ex.r_14[9] ),
    .S1(_10266_),
    .X(_10642_));
 sg13g2_a22oi_1 _17433_ (.Y(_10643_),
    .B1(_10642_),
    .B2(_10231_),
    .A2(_10641_),
    .A1(_10370_));
 sg13g2_nand4_1 _17434_ (.B(_10635_),
    .C(_10639_),
    .A(net540),
    .Y(_10644_),
    .D(_10643_));
 sg13g2_o21ai_1 _17435_ (.B1(_10644_),
    .Y(_10645_),
    .A1(_10627_),
    .A2(net491));
 sg13g2_mux2_1 _17436_ (.A0(_10626_),
    .A1(_10645_),
    .S(_10351_),
    .X(_10646_));
 sg13g2_buf_1 _17437_ (.A(_10646_),
    .X(_10647_));
 sg13g2_nand3_1 _17438_ (.B(_10326_),
    .C(_10647_),
    .A(_10175_),
    .Y(_10648_));
 sg13g2_a21oi_1 _17439_ (.A1(_10625_),
    .A2(_10648_),
    .Y(_10649_),
    .B1(_10522_));
 sg13g2_buf_1 _17440_ (.A(_10649_),
    .X(_10650_));
 sg13g2_inv_1 _17441_ (.Y(\cpu.ex.c_mult_off[2] ),
    .A(_10175_));
 sg13g2_buf_2 _17442_ (.A(_00291_),
    .X(_10651_));
 sg13g2_buf_1 _17443_ (.A(\cpu.addr[10] ),
    .X(_10652_));
 sg13g2_and2_1 _17444_ (.A(net869),
    .B(\cpu.ex.r_11[10] ),
    .X(_10653_));
 sg13g2_a21oi_1 _17445_ (.A1(net750),
    .A2(\cpu.ex.r_9[10] ),
    .Y(_10654_),
    .B1(_10653_));
 sg13g2_nor3_1 _17446_ (.A(net656),
    .B(_10413_),
    .C(_10654_),
    .Y(_10655_));
 sg13g2_nor3_1 _17447_ (.A(_00268_),
    .B(_10333_),
    .C(_10376_),
    .Y(_10656_));
 sg13g2_and2_1 _17448_ (.A(_10314_),
    .B(_10072_),
    .X(_10657_));
 sg13g2_a21oi_1 _17449_ (.A1(net749),
    .A2(\cpu.ex.r_epc[10] ),
    .Y(_10658_),
    .B1(_10657_));
 sg13g2_mux2_1 _17450_ (.A0(\cpu.ex.r_stmp[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(net872),
    .X(_10659_));
 sg13g2_nand3_1 _17451_ (.B(net654),
    .C(_10659_),
    .A(net742),
    .Y(_10660_));
 sg13g2_o21ai_1 _17452_ (.B1(_10660_),
    .Y(_10661_),
    .A1(_10309_),
    .A2(_10658_));
 sg13g2_buf_1 _17453_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10662_));
 sg13g2_a22oi_1 _17454_ (.Y(_10663_),
    .B1(net653),
    .B2(_10662_),
    .A2(net652),
    .A1(\cpu.ex.r_8[10] ));
 sg13g2_nor2b_1 _17455_ (.A(_10663_),
    .B_N(_10301_),
    .Y(_10664_));
 sg13g2_nor4_1 _17456_ (.A(_10655_),
    .B(_10656_),
    .C(_10661_),
    .D(_10664_),
    .Y(_10665_));
 sg13g2_nand3_1 _17457_ (.B(\cpu.ex.r_lr[10] ),
    .C(net659),
    .A(net658),
    .Y(_10666_));
 sg13g2_nand3_1 _17458_ (.B(\cpu.ex.r_12[10] ),
    .C(net748),
    .A(net656),
    .Y(_10667_));
 sg13g2_a21oi_1 _17459_ (.A1(_10666_),
    .A2(_10667_),
    .Y(_10668_),
    .B1(net740));
 sg13g2_inv_1 _17460_ (.Y(_10669_),
    .A(_10668_));
 sg13g2_nor2_1 _17461_ (.A(net749),
    .B(_10337_),
    .Y(_10670_));
 sg13g2_nor2_1 _17462_ (.A(net745),
    .B(_10263_),
    .Y(_10671_));
 sg13g2_a22oi_1 _17463_ (.Y(_10672_),
    .B1(_10671_),
    .B2(\cpu.ex.r_10[10] ),
    .A2(_10670_),
    .A1(\cpu.ex.r_13[10] ));
 sg13g2_nand2b_1 _17464_ (.Y(_10673_),
    .B(net660),
    .A_N(_10672_));
 sg13g2_nand4_1 _17465_ (.B(_10665_),
    .C(_10669_),
    .A(net491),
    .Y(_10674_),
    .D(_10673_));
 sg13g2_o21ai_1 _17466_ (.B1(_10674_),
    .Y(_10675_),
    .A1(net1089),
    .A2(net491));
 sg13g2_buf_2 _17467_ (.A(_00290_),
    .X(_10676_));
 sg13g2_nor2_1 _17468_ (.A(net1094),
    .B(_10221_),
    .Y(_10677_));
 sg13g2_a22oi_1 _17469_ (.Y(_10678_),
    .B1(_10415_),
    .B2(_10118_),
    .A2(_10251_),
    .A1(\cpu.ex.r_11[11] ));
 sg13g2_mux2_1 _17470_ (.A0(\cpu.ex.r_8[11] ),
    .A1(\cpu.ex.r_10[11] ),
    .S(net869),
    .X(_10679_));
 sg13g2_mux2_1 _17471_ (.A0(\cpu.ex.r_lr[11] ),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net869),
    .X(_10680_));
 sg13g2_a22oi_1 _17472_ (.Y(_10681_),
    .B1(_10680_),
    .B2(_10370_),
    .A2(_10679_),
    .A1(_10231_));
 sg13g2_o21ai_1 _17473_ (.B1(_10681_),
    .Y(_10682_),
    .A1(_10226_),
    .A2(_10678_));
 sg13g2_nand2_1 _17474_ (.Y(_10683_),
    .A(_10248_),
    .B(_10682_));
 sg13g2_a22oi_1 _17475_ (.Y(_10684_),
    .B1(_10388_),
    .B2(\cpu.ex.r_stmp[11] ),
    .A2(net652),
    .A1(\cpu.ex.r_12[11] ));
 sg13g2_nor2_1 _17476_ (.A(_10381_),
    .B(_10684_),
    .Y(_10685_));
 sg13g2_a22oi_1 _17477_ (.Y(_10686_),
    .B1(_10425_),
    .B2(_10109_),
    .A2(_10373_),
    .A1(\cpu.ex.r_9[11] ));
 sg13g2_nor2_1 _17478_ (.A(_10413_),
    .B(_10686_),
    .Y(_10687_));
 sg13g2_nor2_1 _17479_ (.A(_10685_),
    .B(_10687_),
    .Y(_10688_));
 sg13g2_a22oi_1 _17480_ (.Y(_10689_),
    .B1(net653),
    .B2(\cpu.ex.r_mult[27] ),
    .A2(net652),
    .A1(\cpu.ex.r_13[11] ));
 sg13g2_nor2_1 _17481_ (.A(_10240_),
    .B(_10689_),
    .Y(_10690_));
 sg13g2_a21oi_1 _17482_ (.A1(\cpu.ex.r_14[11] ),
    .A2(_10334_),
    .Y(_10691_),
    .B1(_10690_));
 sg13g2_nand4_1 _17483_ (.B(_10683_),
    .C(_10688_),
    .A(net491),
    .Y(_10692_),
    .D(_10691_));
 sg13g2_nand2b_1 _17484_ (.Y(_10693_),
    .B(_10692_),
    .A_N(_10677_));
 sg13g2_mux4_1 _17485_ (.S0(_10351_),
    .A0(_10651_),
    .A1(_10675_),
    .A2(_10676_),
    .A3(_10693_),
    .S1(\cpu.ex.c_mult_off[0] ),
    .X(_10694_));
 sg13g2_buf_2 _17486_ (.A(_00293_),
    .X(_10695_));
 sg13g2_nand2b_1 _17487_ (.Y(_10696_),
    .B(_10224_),
    .A_N(_09011_));
 sg13g2_buf_1 _17488_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10697_));
 sg13g2_a22oi_1 _17489_ (.Y(_10698_),
    .B1(net653),
    .B2(_10697_),
    .A2(_10420_),
    .A1(\cpu.ex.r_8[8] ));
 sg13g2_nand2b_1 _17490_ (.Y(_10699_),
    .B(_10301_),
    .A_N(_10698_));
 sg13g2_a22oi_1 _17491_ (.Y(_10700_),
    .B1(_10671_),
    .B2(\cpu.ex.r_10[8] ),
    .A2(_10670_),
    .A1(\cpu.ex.r_13[8] ));
 sg13g2_nand2b_1 _17492_ (.Y(_10701_),
    .B(net660),
    .A_N(_10700_));
 sg13g2_a22oi_1 _17493_ (.Y(_10702_),
    .B1(_10388_),
    .B2(\cpu.ex.r_stmp[8] ),
    .A2(_10420_),
    .A1(\cpu.ex.r_12[8] ));
 sg13g2_nor2_1 _17494_ (.A(_10381_),
    .B(_10702_),
    .Y(_10703_));
 sg13g2_inv_1 _17495_ (.Y(_10704_),
    .A(_00266_));
 sg13g2_a22oi_1 _17496_ (.Y(_10705_),
    .B1(_10425_),
    .B2(_10704_),
    .A2(_10373_),
    .A1(\cpu.ex.r_9[8] ));
 sg13g2_nor2_1 _17497_ (.A(_10413_),
    .B(_10705_),
    .Y(_10706_));
 sg13g2_mux2_1 _17498_ (.A0(\cpu.ex.r_lr[8] ),
    .A1(\cpu.ex.r_epc[8] ),
    .S(net869),
    .X(_10707_));
 sg13g2_nand3_1 _17499_ (.B(net659),
    .C(_10707_),
    .A(net746),
    .Y(_10708_));
 sg13g2_nand3_1 _17500_ (.B(_10441_),
    .C(_10320_),
    .A(\cpu.ex.r_14[8] ),
    .Y(_10709_));
 sg13g2_nand3_1 _17501_ (.B(net655),
    .C(_10378_),
    .A(\cpu.ex.r_11[8] ),
    .Y(_10710_));
 sg13g2_nand3_1 _17502_ (.B(_10281_),
    .C(_10329_),
    .A(\cpu.ex.r_mult[24] ),
    .Y(_10711_));
 sg13g2_nand4_1 _17503_ (.B(_10709_),
    .C(_10710_),
    .A(_10708_),
    .Y(_10712_),
    .D(_10711_));
 sg13g2_nor3_1 _17504_ (.A(_10703_),
    .B(_10706_),
    .C(_10712_),
    .Y(_10713_));
 sg13g2_nand4_1 _17505_ (.B(_10699_),
    .C(_10701_),
    .A(net540),
    .Y(_10714_),
    .D(_10713_));
 sg13g2_nand2_1 _17506_ (.Y(_10715_),
    .A(_10696_),
    .B(_10714_));
 sg13g2_mux2_1 _17507_ (.A0(_10695_),
    .A1(_10715_),
    .S(_10351_),
    .X(_10716_));
 sg13g2_buf_2 _17508_ (.A(_10716_),
    .X(_10717_));
 sg13g2_a22oi_1 _17509_ (.Y(_10718_),
    .B1(_10717_),
    .B2(_10180_),
    .A2(_10694_),
    .A1(\cpu.ex.c_mult_off[1] ));
 sg13g2_nor3_1 _17510_ (.A(_10522_),
    .B(\cpu.ex.c_mult_off[2] ),
    .C(_10718_),
    .Y(_10719_));
 sg13g2_buf_1 _17511_ (.A(_10719_),
    .X(_10720_));
 sg13g2_or3_1 _17512_ (.A(_10524_),
    .B(_10650_),
    .C(_10720_),
    .X(_10721_));
 sg13g2_buf_1 _17513_ (.A(_10721_),
    .X(_10722_));
 sg13g2_buf_1 _17514_ (.A(_09217_),
    .X(_10723_));
 sg13g2_nand2_1 _17515_ (.Y(_10724_),
    .A(_09202_),
    .B(net737));
 sg13g2_buf_1 _17516_ (.A(_10724_),
    .X(_10725_));
 sg13g2_or2_1 _17517_ (.X(_10726_),
    .B(_10163_),
    .A(net1095));
 sg13g2_buf_1 _17518_ (.A(_10726_),
    .X(_10727_));
 sg13g2_nor2_1 _17519_ (.A(_10159_),
    .B(_10727_),
    .Y(_10728_));
 sg13g2_and2_1 _17520_ (.A(net758),
    .B(net665),
    .X(_10729_));
 sg13g2_mux2_1 _17521_ (.A0(\cpu.ex.r_9[5] ),
    .A1(\cpu.ex.r_13[5] ),
    .S(_10120_),
    .X(_10730_));
 sg13g2_nand2b_1 _17522_ (.Y(_10731_),
    .B(_10101_),
    .A_N(_10115_));
 sg13g2_buf_1 _17523_ (.A(_10731_),
    .X(_10732_));
 sg13g2_nor2_1 _17524_ (.A(net752),
    .B(_10732_),
    .Y(_10733_));
 sg13g2_a22oi_1 _17525_ (.Y(_10734_),
    .B1(_10730_),
    .B2(_10733_),
    .A2(_10729_),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_inv_2 _17526_ (.Y(_10735_),
    .A(net879));
 sg13g2_mux4_1 _17527_ (.S0(_10126_),
    .A0(_10434_),
    .A1(\cpu.ex.r_11[5] ),
    .A2(\cpu.ex.r_mult[21] ),
    .A3(\cpu.ex.r_epc[5] ),
    .S1(_10735_),
    .X(_10736_));
 sg13g2_nand2_1 _17528_ (.Y(_10737_),
    .A(_10108_),
    .B(_10736_));
 sg13g2_nor2_1 _17529_ (.A(net1092),
    .B(net1093),
    .Y(_10738_));
 sg13g2_buf_2 _17530_ (.A(_10738_),
    .X(_10739_));
 sg13g2_and2_1 _17531_ (.A(net1092),
    .B(net1093),
    .X(_10740_));
 sg13g2_buf_1 _17532_ (.A(_10740_),
    .X(_10741_));
 sg13g2_buf_1 _17533_ (.A(_10741_),
    .X(_10742_));
 sg13g2_a22oi_1 _17534_ (.Y(_10743_),
    .B1(net736),
    .B2(\cpu.ex.r_14[5] ),
    .A2(_10739_),
    .A1(\cpu.ex.r_8[5] ));
 sg13g2_nor2b_1 _17535_ (.A(net1008),
    .B_N(net879),
    .Y(_10744_));
 sg13g2_buf_2 _17536_ (.A(_10744_),
    .X(_10745_));
 sg13g2_nand2b_1 _17537_ (.Y(_10746_),
    .B(_10745_),
    .A_N(_10743_));
 sg13g2_nor2b_1 _17538_ (.A(net878),
    .B_N(net881),
    .Y(_10747_));
 sg13g2_buf_2 _17539_ (.A(_10747_),
    .X(_10748_));
 sg13g2_nand3b_1 _17540_ (.B(net880),
    .C(\cpu.ex.r_stmp[5] ),
    .Y(_10749_),
    .A_N(net876));
 sg13g2_nand3b_1 _17541_ (.B(net756),
    .C(\cpu.ex.r_10[5] ),
    .Y(_10750_),
    .A_N(net880));
 sg13g2_nand2_1 _17542_ (.Y(_10751_),
    .A(_10749_),
    .B(_10750_));
 sg13g2_nand3b_1 _17543_ (.B(net753),
    .C(\cpu.ex.r_lr[5] ),
    .Y(_10752_),
    .A_N(net881));
 sg13g2_nand3b_1 _17544_ (.B(net881),
    .C(_10448_),
    .Y(_10753_),
    .A_N(net878));
 sg13g2_nand2_1 _17545_ (.Y(_10754_),
    .A(_10752_),
    .B(_10753_));
 sg13g2_a22oi_1 _17546_ (.Y(_10755_),
    .B1(_10754_),
    .B2(_10103_),
    .A2(_10751_),
    .A1(_10748_));
 sg13g2_nand4_1 _17547_ (.B(_10737_),
    .C(_10746_),
    .A(_10734_),
    .Y(_10756_),
    .D(_10755_));
 sg13g2_a22oi_1 _17548_ (.Y(_10757_),
    .B1(net541),
    .B2(_10756_),
    .A2(net492),
    .A1(_09818_));
 sg13g2_buf_2 _17549_ (.A(_10757_),
    .X(_10758_));
 sg13g2_nor2b_1 _17550_ (.A(_08701_),
    .B_N(net1095),
    .Y(_10759_));
 sg13g2_nor4_1 _17551_ (.A(net1004),
    .B(net1095),
    .C(_10163_),
    .D(\cpu.dec.imm[5] ),
    .Y(_10760_));
 sg13g2_or2_1 _17552_ (.X(_10761_),
    .B(_10760_),
    .A(_10759_));
 sg13g2_a21oi_1 _17553_ (.A1(_10728_),
    .A2(_10758_),
    .Y(_10762_),
    .B1(_10761_));
 sg13g2_buf_1 _17554_ (.A(_10762_),
    .X(_10763_));
 sg13g2_buf_1 _17555_ (.A(_00306_),
    .X(_10764_));
 sg13g2_and3_1 _17556_ (.X(_10765_),
    .A(\cpu.ex.r_10[4] ),
    .B(net874),
    .C(net879));
 sg13g2_a221oi_1 _17557_ (.B2(_10462_),
    .C1(_10765_),
    .B1(_10137_),
    .A1(\cpu.ex.r_8[4] ),
    .Y(_10766_),
    .A2(_10129_));
 sg13g2_nor2_1 _17558_ (.A(net1008),
    .B(net1005),
    .Y(_10767_));
 sg13g2_buf_1 _17559_ (.A(_10767_),
    .X(_10768_));
 sg13g2_nand2b_1 _17560_ (.Y(_10769_),
    .B(net735),
    .A_N(_10766_));
 sg13g2_nor2b_1 _17561_ (.A(net881),
    .B_N(net875),
    .Y(_10770_));
 sg13g2_nor2_1 _17562_ (.A(net1008),
    .B(net1007),
    .Y(_10771_));
 sg13g2_and3_1 _17563_ (.X(_10772_),
    .A(\cpu.ex.r_13[4] ),
    .B(net1008),
    .C(net879));
 sg13g2_a21o_1 _17564_ (.A2(_10771_),
    .A1(_08735_),
    .B1(_10772_),
    .X(_10773_));
 sg13g2_inv_1 _17565_ (.Y(_10774_),
    .A(\cpu.ex.r_12[4] ));
 sg13g2_nand3b_1 _17566_ (.B(net874),
    .C(\cpu.ex.r_stmp[4] ),
    .Y(_10775_),
    .A_N(net879));
 sg13g2_o21ai_1 _17567_ (.B1(_10775_),
    .Y(_10776_),
    .A1(_10774_),
    .A2(_10732_));
 sg13g2_nor2b_1 _17568_ (.A(_10088_),
    .B_N(net1093),
    .Y(_10777_));
 sg13g2_buf_2 _17569_ (.A(_10777_),
    .X(_10778_));
 sg13g2_nand3b_1 _17570_ (.B(_10149_),
    .C(\cpu.ex.r_mult[20] ),
    .Y(_10779_),
    .A_N(_10121_));
 sg13g2_nand3b_1 _17571_ (.B(_10121_),
    .C(\cpu.ex.r_11[4] ),
    .Y(_10780_),
    .A_N(_10119_));
 sg13g2_nand2_1 _17572_ (.Y(_10781_),
    .A(_10131_),
    .B(net874));
 sg13g2_a21oi_1 _17573_ (.A1(_10779_),
    .A2(_10780_),
    .Y(_10782_),
    .B1(_10781_));
 sg13g2_a221oi_1 _17574_ (.B2(_10778_),
    .C1(_10782_),
    .B1(_10776_),
    .A1(_10770_),
    .Y(_10783_),
    .A2(_10773_));
 sg13g2_nand3_1 _17575_ (.B(net878),
    .C(_10739_),
    .A(\cpu.ex.r_9[4] ),
    .Y(_10784_));
 sg13g2_nand3_1 _17576_ (.B(_10142_),
    .C(net736),
    .A(\cpu.ex.r_14[4] ),
    .Y(_10785_));
 sg13g2_a21o_1 _17577_ (.A2(_10785_),
    .A1(_10784_),
    .B1(_10735_),
    .X(_10786_));
 sg13g2_mux2_1 _17578_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_epc[4] ),
    .S(net1006),
    .X(_10787_));
 sg13g2_nor2b_1 _17579_ (.A(_00262_),
    .B_N(_10151_),
    .Y(_10788_));
 sg13g2_a22oi_1 _17580_ (.Y(_10789_),
    .B1(_10788_),
    .B2(_10112_),
    .A2(_10787_),
    .A1(_10103_));
 sg13g2_nand2b_1 _17581_ (.Y(_10790_),
    .B(net753),
    .A_N(_10789_));
 sg13g2_and4_1 _17582_ (.A(_10769_),
    .B(_10783_),
    .C(_10786_),
    .D(_10790_),
    .X(_10791_));
 sg13g2_nand2b_1 _17583_ (.Y(_10792_),
    .B(net1095),
    .A_N(\cpu.ex.pc[4] ));
 sg13g2_nand3_1 _17584_ (.B(net541),
    .C(_10792_),
    .A(_10157_),
    .Y(_10793_));
 sg13g2_nor4_1 _17585_ (.A(_09359_),
    .B(_10158_),
    .C(_10084_),
    .D(_10092_),
    .Y(_10794_));
 sg13g2_a21o_1 _17586_ (.A2(\cpu.dec.imm[4] ),
    .A1(net873),
    .B1(_10727_),
    .X(_10795_));
 sg13g2_o21ai_1 _17587_ (.B1(_10792_),
    .Y(_10796_),
    .A1(_10794_),
    .A2(_10795_));
 sg13g2_o21ai_1 _17588_ (.B1(_10796_),
    .Y(_10797_),
    .A1(_10791_),
    .A2(_10793_));
 sg13g2_buf_8 _17589_ (.A(_10797_),
    .X(_10798_));
 sg13g2_or2_1 _17590_ (.X(_10799_),
    .B(net373),
    .A(net1088));
 sg13g2_a21o_1 _17591_ (.A2(_10758_),
    .A1(_10728_),
    .B1(_10761_),
    .X(_10800_));
 sg13g2_buf_2 _17592_ (.A(_10800_),
    .X(_10801_));
 sg13g2_nand4_1 _17593_ (.B(_10783_),
    .C(_10786_),
    .A(_10769_),
    .Y(_10802_),
    .D(_10790_));
 sg13g2_nand2b_1 _17594_ (.Y(_10803_),
    .B(_10802_),
    .A_N(_10793_));
 sg13g2_and2_1 _17595_ (.A(_10796_),
    .B(_10803_),
    .X(_10804_));
 sg13g2_buf_1 _17596_ (.A(_10804_),
    .X(_10805_));
 sg13g2_nand3b_1 _17597_ (.B(_10801_),
    .C(_10805_),
    .Y(_10806_),
    .A_N(net1088));
 sg13g2_buf_2 _17598_ (.A(_00305_),
    .X(_10807_));
 sg13g2_a22oi_1 _17599_ (.Y(_10808_),
    .B1(_10806_),
    .B2(_10807_),
    .A2(_10799_),
    .A1(_10763_));
 sg13g2_buf_1 _17600_ (.A(_00308_),
    .X(_10809_));
 sg13g2_inv_1 _17601_ (.Y(_10810_),
    .A(_10809_));
 sg13g2_buf_1 _17602_ (.A(\cpu.dec.imm[2] ),
    .X(_10811_));
 sg13g2_nor4_1 _17603_ (.A(_10811_),
    .B(net1004),
    .C(net1095),
    .D(_10163_),
    .Y(_10812_));
 sg13g2_a21oi_2 _17604_ (.B1(_10812_),
    .Y(_10813_),
    .A2(net1009),
    .A1(_08159_));
 sg13g2_a21o_1 _17605_ (.A2(_10103_),
    .A1(_10100_),
    .B1(_10094_),
    .X(_10814_));
 sg13g2_buf_2 _17606_ (.A(_10814_),
    .X(_10815_));
 sg13g2_and2_1 _17607_ (.A(net754),
    .B(net877),
    .X(_10816_));
 sg13g2_mux2_1 _17608_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(_10363_),
    .S(net875),
    .X(_10817_));
 sg13g2_or2_1 _17609_ (.X(_10818_),
    .B(net1007),
    .A(net1006));
 sg13g2_nor2_1 _17610_ (.A(_10142_),
    .B(_10818_),
    .Y(_10819_));
 sg13g2_and2_1 _17611_ (.A(net1006),
    .B(net1007),
    .X(_10820_));
 sg13g2_buf_1 _17612_ (.A(_10820_),
    .X(_10821_));
 sg13g2_and3_1 _17613_ (.X(_10822_),
    .A(\cpu.ex.r_10[2] ),
    .B(net735),
    .C(_10821_));
 sg13g2_a221oi_1 _17614_ (.B2(_10819_),
    .C1(_10822_),
    .B1(_10817_),
    .A1(\cpu.ex.r_9[2] ),
    .Y(_10823_),
    .A2(_10816_));
 sg13g2_mux2_1 _17615_ (.A0(net1114),
    .A1(\cpu.ex.r_stmp[2] ),
    .S(net1006),
    .X(_10824_));
 sg13g2_a221oi_1 _17616_ (.B2(_10735_),
    .C1(net878),
    .B1(_10824_),
    .A1(\cpu.ex.r_12[2] ),
    .Y(_10825_),
    .A2(net754));
 sg13g2_buf_1 _17617_ (.A(net880),
    .X(_10826_));
 sg13g2_nand2_2 _17618_ (.Y(_10827_),
    .A(_10151_),
    .B(net879));
 sg13g2_o21ai_1 _17619_ (.B1(net878),
    .Y(_10828_),
    .A1(_00260_),
    .A2(_10827_));
 sg13g2_nand3b_1 _17620_ (.B(net734),
    .C(_10828_),
    .Y(_10829_),
    .A_N(_10825_));
 sg13g2_and2_1 _17621_ (.A(net1008),
    .B(net879),
    .X(_10830_));
 sg13g2_buf_1 _17622_ (.A(_10830_),
    .X(_10831_));
 sg13g2_nand3b_1 _17623_ (.B(net874),
    .C(\cpu.ex.r_11[2] ),
    .Y(_10832_),
    .A_N(net1005));
 sg13g2_nand3b_1 _17624_ (.B(net875),
    .C(\cpu.ex.r_13[2] ),
    .Y(_10833_),
    .A_N(net874));
 sg13g2_nand2_1 _17625_ (.Y(_10834_),
    .A(_10832_),
    .B(_10833_));
 sg13g2_inv_1 _17626_ (.Y(_10835_),
    .A(\cpu.ex.r_8[2] ));
 sg13g2_or2_1 _17627_ (.X(_10836_),
    .B(net1005),
    .A(net1006));
 sg13g2_buf_1 _17628_ (.A(_10836_),
    .X(_10837_));
 sg13g2_nand3_1 _17629_ (.B(net874),
    .C(net875),
    .A(\cpu.ex.r_14[2] ),
    .Y(_10838_));
 sg13g2_o21ai_1 _17630_ (.B1(_10838_),
    .Y(_10839_),
    .A1(_10835_),
    .A2(_10837_));
 sg13g2_a22oi_1 _17631_ (.Y(_10840_),
    .B1(_10839_),
    .B2(_10745_),
    .A2(_10834_),
    .A1(_10831_));
 sg13g2_mux2_1 _17632_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(\cpu.ex.r_mult[18] ),
    .S(net1005),
    .X(_10841_));
 sg13g2_a22oi_1 _17633_ (.Y(_10842_),
    .B1(_10841_),
    .B2(net753),
    .A2(net735),
    .A1(_10386_));
 sg13g2_nand2b_1 _17634_ (.Y(_10843_),
    .B(net663),
    .A_N(_10842_));
 sg13g2_and4_1 _17635_ (.A(_10823_),
    .B(_10829_),
    .C(_10840_),
    .D(_10843_),
    .X(_10844_));
 sg13g2_nand2_1 _17636_ (.Y(_10845_),
    .A(_10157_),
    .B(_10165_));
 sg13g2_a21oi_1 _17637_ (.A1(_09082_),
    .A2(_10094_),
    .Y(_10846_),
    .B1(_10845_));
 sg13g2_o21ai_1 _17638_ (.B1(_10846_),
    .Y(_10847_),
    .A1(_10815_),
    .A2(_10844_));
 sg13g2_buf_2 _17639_ (.A(_10847_),
    .X(_10848_));
 sg13g2_nand2_1 _17640_ (.Y(_10849_),
    .A(_10813_),
    .B(_10848_));
 sg13g2_buf_2 _17641_ (.A(_10849_),
    .X(_10850_));
 sg13g2_buf_2 _17642_ (.A(_00307_),
    .X(_10851_));
 sg13g2_buf_1 _17643_ (.A(\cpu.dec.imm[3] ),
    .X(_10852_));
 sg13g2_nor2_1 _17644_ (.A(_09130_),
    .B(net873),
    .Y(_10853_));
 sg13g2_a221oi_1 _17645_ (.B2(_10853_),
    .C1(_10727_),
    .B1(_10094_),
    .A1(_10852_),
    .Y(_10854_),
    .A2(net873));
 sg13g2_nand3_1 _17646_ (.B(net753),
    .C(_10770_),
    .A(\cpu.ex.r_13[3] ),
    .Y(_10855_));
 sg13g2_nor2b_1 _17647_ (.A(net1093),
    .B_N(net1092),
    .Y(_10856_));
 sg13g2_buf_1 _17648_ (.A(_10856_),
    .X(_10857_));
 sg13g2_nand3_1 _17649_ (.B(_10142_),
    .C(_10857_),
    .A(\cpu.ex.r_10[3] ),
    .Y(_10858_));
 sg13g2_buf_2 _17650_ (.A(_10735_),
    .X(_10859_));
 sg13g2_a21oi_1 _17651_ (.A1(_10855_),
    .A2(_10858_),
    .Y(_10860_),
    .B1(net651));
 sg13g2_a22oi_1 _17652_ (.Y(_10861_),
    .B1(_10150_),
    .B2(net1115),
    .A2(net751),
    .A1(\cpu.ex.r_8[3] ));
 sg13g2_nor2b_1 _17653_ (.A(_10861_),
    .B_N(net758),
    .Y(_10862_));
 sg13g2_nand3_1 _17654_ (.B(net758),
    .C(net665),
    .A(\cpu.ex.r_12[3] ),
    .Y(_10863_));
 sg13g2_mux2_1 _17655_ (.A0(\cpu.ex.r_stmp[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net876),
    .X(_10864_));
 sg13g2_nand3_1 _17656_ (.B(net736),
    .C(_10864_),
    .A(_10142_),
    .Y(_10865_));
 sg13g2_mux2_1 _17657_ (.A0(_10246_),
    .A1(\cpu.ex.r_epc[3] ),
    .S(_10131_),
    .X(_10866_));
 sg13g2_nand3_1 _17658_ (.B(net663),
    .C(_10866_),
    .A(net755),
    .Y(_10867_));
 sg13g2_nand3_1 _17659_ (.B(_10865_),
    .C(_10867_),
    .A(_10863_),
    .Y(_10868_));
 sg13g2_nor3_1 _17660_ (.A(_10860_),
    .B(_10862_),
    .C(_10868_),
    .Y(_10869_));
 sg13g2_nand2b_1 _17661_ (.Y(_10870_),
    .B(net880),
    .A_N(_00261_));
 sg13g2_nand2_1 _17662_ (.Y(_10871_),
    .A(\cpu.ex.r_11[3] ),
    .B(net755));
 sg13g2_a21oi_1 _17663_ (.A1(_10870_),
    .A2(_10871_),
    .Y(_10872_),
    .B1(_10827_));
 sg13g2_a22oi_1 _17664_ (.Y(_10873_),
    .B1(net736),
    .B2(\cpu.ex.r_mult[19] ),
    .A2(_10739_),
    .A1(\cpu.ex.r_lr[3] ));
 sg13g2_nand3b_1 _17665_ (.B(_10148_),
    .C(\cpu.ex.r_9[3] ),
    .Y(_10874_),
    .A_N(net875));
 sg13g2_nand3b_1 _17666_ (.B(_10149_),
    .C(_10242_),
    .Y(_10875_),
    .A_N(_10148_));
 sg13g2_a21o_1 _17667_ (.A2(_10875_),
    .A1(_10874_),
    .B1(net881),
    .X(_10876_));
 sg13g2_o21ai_1 _17668_ (.B1(_10876_),
    .Y(_10877_),
    .A1(net756),
    .A2(_10873_));
 sg13g2_o21ai_1 _17669_ (.B1(net664),
    .Y(_10878_),
    .A1(_10872_),
    .A2(_10877_));
 sg13g2_nand3_1 _17670_ (.B(_10869_),
    .C(_10878_),
    .A(_10854_),
    .Y(_10879_));
 sg13g2_nand2_1 _17671_ (.Y(_10880_),
    .A(_10157_),
    .B(_10105_));
 sg13g2_a22oi_1 _17672_ (.Y(_10881_),
    .B1(_10854_),
    .B2(_10880_),
    .A2(net1009),
    .A1(_08149_));
 sg13g2_and2_1 _17673_ (.A(_10879_),
    .B(_10881_),
    .X(_10882_));
 sg13g2_buf_8 _17674_ (.A(_10882_),
    .X(_10883_));
 sg13g2_nor2_1 _17675_ (.A(_10851_),
    .B(net341),
    .Y(_10884_));
 sg13g2_a21oi_1 _17676_ (.A1(_10810_),
    .A2(_10850_),
    .Y(_10885_),
    .B1(_10884_));
 sg13g2_nand2b_1 _17677_ (.Y(_10886_),
    .B(_10885_),
    .A_N(_10808_));
 sg13g2_nor2_2 _17678_ (.A(_00309_),
    .B(_09205_),
    .Y(_10887_));
 sg13g2_buf_1 _17679_ (.A(\cpu.dec.imm[1] ),
    .X(_10888_));
 sg13g2_nor2_1 _17680_ (.A(_09811_),
    .B(net873),
    .Y(_10889_));
 sg13g2_a221oi_1 _17681_ (.B2(_10889_),
    .C1(_10727_),
    .B1(_10094_),
    .A1(_10888_),
    .Y(_10890_),
    .A2(_10159_));
 sg13g2_buf_1 _17682_ (.A(_10890_),
    .X(_10891_));
 sg13g2_a22oi_1 _17683_ (.Y(_10892_),
    .B1(_10136_),
    .B2(\cpu.ex.r_stmp[1] ),
    .A2(_10128_),
    .A1(\cpu.ex.r_12[1] ));
 sg13g2_nor2_1 _17684_ (.A(net753),
    .B(_10892_),
    .Y(_10893_));
 sg13g2_and2_1 _17685_ (.A(\cpu.ex.mmu_read[1] ),
    .B(_10819_),
    .X(_10894_));
 sg13g2_o21ai_1 _17686_ (.B1(net734),
    .Y(_10895_),
    .A1(_10893_),
    .A2(_10894_));
 sg13g2_mux2_1 _17687_ (.A0(\cpu.ex.r_10[1] ),
    .A1(\cpu.ex.r_11[1] ),
    .S(_10098_),
    .X(_10896_));
 sg13g2_nand2_1 _17688_ (.Y(_10897_),
    .A(_10857_),
    .B(_10896_));
 sg13g2_nor2b_1 _17689_ (.A(_00259_),
    .B_N(net1006),
    .Y(_10898_));
 sg13g2_nor2b_1 _17690_ (.A(net1006),
    .B_N(\cpu.ex.r_13[1] ),
    .Y(_10899_));
 sg13g2_and2_1 _17691_ (.A(net1008),
    .B(net1093),
    .X(_10900_));
 sg13g2_buf_2 _17692_ (.A(_10900_),
    .X(_10901_));
 sg13g2_o21ai_1 _17693_ (.B1(_10901_),
    .Y(_10902_),
    .A1(_10898_),
    .A2(_10899_));
 sg13g2_nand3_1 _17694_ (.B(_10897_),
    .C(_10902_),
    .A(net876),
    .Y(_10903_));
 sg13g2_a22oi_1 _17695_ (.Y(_10904_),
    .B1(_10778_),
    .B2(_10288_),
    .A2(net877),
    .A1(\cpu.ex.r_lr[1] ));
 sg13g2_mux2_1 _17696_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(net1005),
    .X(_10905_));
 sg13g2_a21oi_1 _17697_ (.A1(_10108_),
    .A2(_10905_),
    .Y(_10906_),
    .B1(net876));
 sg13g2_o21ai_1 _17698_ (.B1(_10906_),
    .Y(_10907_),
    .A1(net881),
    .A2(_10904_));
 sg13g2_a22oi_1 _17699_ (.Y(_10908_),
    .B1(_10741_),
    .B2(\cpu.ex.r_14[1] ),
    .A2(_10739_),
    .A1(\cpu.ex.r_8[1] ));
 sg13g2_inv_1 _17700_ (.Y(_10909_),
    .A(_10908_));
 sg13g2_nand3_1 _17701_ (.B(net878),
    .C(_10128_),
    .A(\cpu.ex.r_9[1] ),
    .Y(_10910_));
 sg13g2_nand3_1 _17702_ (.B(_10142_),
    .C(_10136_),
    .A(_10318_),
    .Y(_10911_));
 sg13g2_a21oi_1 _17703_ (.A1(_10910_),
    .A2(_10911_),
    .Y(_10912_),
    .B1(net880));
 sg13g2_a221oi_1 _17704_ (.B2(_10745_),
    .C1(_10912_),
    .B1(_10909_),
    .A1(_10903_),
    .Y(_10913_),
    .A2(_10907_));
 sg13g2_a21o_1 _17705_ (.A2(_10913_),
    .A1(_10895_),
    .B1(_10880_),
    .X(_10914_));
 sg13g2_buf_1 _17706_ (.A(_10914_),
    .X(_10915_));
 sg13g2_nor2b_1 _17707_ (.A(net1117),
    .B_N(_10074_),
    .Y(_10916_));
 sg13g2_a21o_1 _17708_ (.A2(net426),
    .A1(net427),
    .B1(_10916_),
    .X(_10917_));
 sg13g2_buf_2 _17709_ (.A(_10917_),
    .X(_10918_));
 sg13g2_nand2b_1 _17710_ (.Y(_10919_),
    .B(net1004),
    .A_N(_10163_));
 sg13g2_a21oi_1 _17711_ (.A1(_08767_),
    .A2(_10094_),
    .Y(_10920_),
    .B1(_10919_));
 sg13g2_buf_1 _17712_ (.A(\cpu.dec.imm[0] ),
    .X(_10921_));
 sg13g2_nor3_1 _17713_ (.A(_10921_),
    .B(_10157_),
    .C(_10163_),
    .Y(_10922_));
 sg13g2_nor2_1 _17714_ (.A(net1095),
    .B(_10922_),
    .Y(_10923_));
 sg13g2_nand2b_1 _17715_ (.Y(_10924_),
    .B(_10923_),
    .A_N(_10920_));
 sg13g2_buf_1 _17716_ (.A(_10924_),
    .X(_10925_));
 sg13g2_nand2_1 _17717_ (.Y(_10926_),
    .A(\cpu.ex.r_9[0] ),
    .B(_10816_));
 sg13g2_mux2_1 _17718_ (.A0(\cpu.ex.r_13[0] ),
    .A1(\cpu.ex.r_15[0] ),
    .S(net874),
    .X(_10927_));
 sg13g2_nand3_1 _17719_ (.B(net756),
    .C(_10927_),
    .A(net753),
    .Y(_10928_));
 sg13g2_mux2_1 _17720_ (.A0(_09073_),
    .A1(\cpu.ex.r_12[0] ),
    .S(net876),
    .X(_10929_));
 sg13g2_nand3_1 _17721_ (.B(_10152_),
    .C(_10929_),
    .A(_10143_),
    .Y(_10930_));
 sg13g2_a21o_1 _17722_ (.A2(_10930_),
    .A1(_10928_),
    .B1(net755),
    .X(_10931_));
 sg13g2_nand3b_1 _17723_ (.B(net880),
    .C(\cpu.ex.r_stmp[0] ),
    .Y(_10932_),
    .A_N(net876));
 sg13g2_nand3b_1 _17724_ (.B(net756),
    .C(\cpu.ex.r_10[0] ),
    .Y(_10933_),
    .A_N(net880));
 sg13g2_a21oi_1 _17725_ (.A1(_10932_),
    .A2(_10933_),
    .Y(_10934_),
    .B1(_10152_));
 sg13g2_and3_1 _17726_ (.X(_10935_),
    .A(\cpu.ex.r_8[0] ),
    .B(_10152_),
    .C(net751));
 sg13g2_o21ai_1 _17727_ (.B1(net752),
    .Y(_10936_),
    .A1(_10934_),
    .A2(_10935_));
 sg13g2_nand3_1 _17728_ (.B(_10931_),
    .C(_10936_),
    .A(_10926_),
    .Y(_10937_));
 sg13g2_mux2_1 _17729_ (.A0(_10343_),
    .A1(\cpu.ex.r_mult[16] ),
    .S(net875),
    .X(_10938_));
 sg13g2_a22oi_1 _17730_ (.Y(_10939_),
    .B1(_10938_),
    .B2(_10735_),
    .A2(net751),
    .A1(\cpu.ex.r_11[0] ));
 sg13g2_nand2_1 _17731_ (.Y(_10940_),
    .A(\cpu.ex.r_14[0] ),
    .B(net665));
 sg13g2_mux2_1 _17732_ (.A0(_10939_),
    .A1(_10940_),
    .S(_10143_),
    .X(_10941_));
 sg13g2_nor2_1 _17733_ (.A(_10153_),
    .B(_10941_),
    .Y(_10942_));
 sg13g2_and2_1 _17734_ (.A(_10106_),
    .B(_10923_),
    .X(_10943_));
 sg13g2_o21ai_1 _17735_ (.B1(_10943_),
    .Y(_10944_),
    .A1(_10937_),
    .A2(_10942_));
 sg13g2_buf_1 _17736_ (.A(_10944_),
    .X(_10945_));
 sg13g2_and2_1 _17737_ (.A(_10925_),
    .B(_10945_),
    .X(_10946_));
 sg13g2_buf_1 _17738_ (.A(_10946_),
    .X(_10947_));
 sg13g2_a221oi_1 _17739_ (.B2(_10918_),
    .C1(_10947_),
    .B1(_10887_),
    .A1(net606),
    .Y(_10948_),
    .A2(_10886_));
 sg13g2_buf_1 _17740_ (.A(_10948_),
    .X(_10949_));
 sg13g2_buf_1 _17741_ (.A(_10161_),
    .X(_10950_));
 sg13g2_mux2_1 _17742_ (.A0(_10416_),
    .A1(\cpu.ex.r_12[7] ),
    .S(net876),
    .X(_10951_));
 sg13g2_a22oi_1 _17743_ (.Y(_10952_),
    .B1(_10951_),
    .B2(_10152_),
    .A2(net663),
    .A1(\cpu.ex.r_stmp[7] ));
 sg13g2_nand3_1 _17744_ (.B(net881),
    .C(net751),
    .A(\cpu.ex.r_10[7] ),
    .Y(_10953_));
 sg13g2_o21ai_1 _17745_ (.B1(_10953_),
    .Y(_10954_),
    .A1(net755),
    .A2(_10952_));
 sg13g2_nor2b_1 _17746_ (.A(_00265_),
    .B_N(net756),
    .Y(_10955_));
 sg13g2_nor2b_1 _17747_ (.A(net756),
    .B_N(\cpu.ex.r_mult[23] ),
    .Y(_10956_));
 sg13g2_o21ai_1 _17748_ (.B1(_10742_),
    .Y(_10957_),
    .A1(_10955_),
    .A2(_10956_));
 sg13g2_nand3_1 _17749_ (.B(net661),
    .C(_10103_),
    .A(\cpu.ex.r_lr[7] ),
    .Y(_10958_));
 sg13g2_nand3_1 _17750_ (.B(_10957_),
    .C(_10958_),
    .A(net753),
    .Y(_10959_));
 sg13g2_o21ai_1 _17751_ (.B1(_10959_),
    .Y(_10960_),
    .A1(_10133_),
    .A2(_10954_));
 sg13g2_a22oi_1 _17752_ (.Y(_10961_),
    .B1(_10137_),
    .B2(\cpu.ex.r_epc[7] ),
    .A2(_10129_),
    .A1(\cpu.ex.r_9[7] ));
 sg13g2_nor2b_1 _17753_ (.A(_10961_),
    .B_N(net877),
    .Y(_10962_));
 sg13g2_and4_1 _17754_ (.A(\cpu.ex.r_14[7] ),
    .B(net752),
    .C(_10826_),
    .D(_10821_),
    .X(_10963_));
 sg13g2_a22oi_1 _17755_ (.Y(_10964_),
    .B1(_10901_),
    .B2(\cpu.ex.r_13[7] ),
    .A2(net735),
    .A1(\cpu.ex.r_8[7] ));
 sg13g2_nor2_1 _17756_ (.A(_10732_),
    .B(_10964_),
    .Y(_10965_));
 sg13g2_a22oi_1 _17757_ (.Y(_10966_),
    .B1(_10771_),
    .B2(_10406_),
    .A2(_10831_),
    .A1(\cpu.ex.r_11[7] ));
 sg13g2_nor2b_1 _17758_ (.A(_10966_),
    .B_N(_10857_),
    .Y(_10967_));
 sg13g2_nor4_1 _17759_ (.A(_10962_),
    .B(_10963_),
    .C(_10965_),
    .D(_10967_),
    .Y(_10968_));
 sg13g2_nand2_1 _17760_ (.Y(_10969_),
    .A(_10960_),
    .B(_10968_));
 sg13g2_a22oi_1 _17761_ (.Y(_10970_),
    .B1(net541),
    .B2(_10969_),
    .A2(net492),
    .A1(_09013_));
 sg13g2_buf_2 _17762_ (.A(_10970_),
    .X(_10971_));
 sg13g2_nor2_1 _17763_ (.A(net1004),
    .B(\cpu.dec.imm[7] ),
    .Y(_10972_));
 sg13g2_a21oi_1 _17764_ (.A1(net868),
    .A2(_10971_),
    .Y(_10973_),
    .B1(_10972_));
 sg13g2_nand2_1 _17765_ (.Y(_10974_),
    .A(_08679_),
    .B(net882));
 sg13g2_o21ai_1 _17766_ (.B1(_10974_),
    .Y(_10975_),
    .A1(_10727_),
    .A2(_10973_));
 sg13g2_buf_2 _17767_ (.A(_10975_),
    .X(_10976_));
 sg13g2_buf_1 _17768_ (.A(_00304_),
    .X(_10977_));
 sg13g2_nor2_1 _17769_ (.A(_10977_),
    .B(net678),
    .Y(_10978_));
 sg13g2_o21ai_1 _17770_ (.B1(_10978_),
    .Y(_10979_),
    .A1(_10501_),
    .A2(_10976_));
 sg13g2_buf_1 _17771_ (.A(_10165_),
    .X(_10980_));
 sg13g2_a22oi_1 _17772_ (.Y(_10981_),
    .B1(_10778_),
    .B2(\cpu.ex.r_14[6] ),
    .A2(net877),
    .A1(\cpu.ex.r_11[6] ));
 sg13g2_nor2_1 _17773_ (.A(_10827_),
    .B(_10981_),
    .Y(_10982_));
 sg13g2_nand2_1 _17774_ (.Y(_10983_),
    .A(_10132_),
    .B(_10122_));
 sg13g2_a22oi_1 _17775_ (.Y(_10984_),
    .B1(net736),
    .B2(_10493_),
    .A2(_10739_),
    .A1(\cpu.ex.r_9[6] ));
 sg13g2_nand3_1 _17776_ (.B(net758),
    .C(net665),
    .A(\cpu.ex.r_12[6] ),
    .Y(_10985_));
 sg13g2_o21ai_1 _17777_ (.B1(_10985_),
    .Y(_10986_),
    .A1(_10983_),
    .A2(_10984_));
 sg13g2_mux4_1 _17778_ (.S0(net878),
    .A0(_10511_),
    .A1(\cpu.ex.r_epc[6] ),
    .A2(\cpu.ex.r_stmp[6] ),
    .A3(_10501_),
    .S1(net875),
    .X(_10987_));
 sg13g2_nor2b_1 _17779_ (.A(_10116_),
    .B_N(\cpu.ex.r_lr[6] ),
    .Y(_10988_));
 sg13g2_a22oi_1 _17780_ (.Y(_10989_),
    .B1(_10988_),
    .B2(_10140_),
    .A2(_10987_),
    .A1(net757));
 sg13g2_nor2_1 _17781_ (.A(_10122_),
    .B(_10989_),
    .Y(_10990_));
 sg13g2_a221oi_1 _17782_ (.B2(\cpu.ex.r_13[6] ),
    .C1(net881),
    .B1(_10901_),
    .A1(\cpu.ex.r_8[6] ),
    .Y(_10991_),
    .A2(_10768_));
 sg13g2_a21oi_1 _17783_ (.A1(\cpu.ex.r_10[6] ),
    .A2(_10768_),
    .Y(_10992_),
    .B1(_10153_));
 sg13g2_nor3_1 _17784_ (.A(net651),
    .B(_10991_),
    .C(_10992_),
    .Y(_10993_));
 sg13g2_or4_1 _17785_ (.A(_10982_),
    .B(_10986_),
    .C(_10990_),
    .D(_10993_),
    .X(_10994_));
 sg13g2_a22oi_1 _17786_ (.Y(_10995_),
    .B1(net541),
    .B2(_10994_),
    .A2(net492),
    .A1(_09010_));
 sg13g2_nor2_1 _17787_ (.A(net1004),
    .B(\cpu.dec.imm[6] ),
    .Y(_10996_));
 sg13g2_a21o_1 _17788_ (.A2(_10995_),
    .A1(net1004),
    .B1(_10996_),
    .X(_10997_));
 sg13g2_nor2b_1 _17789_ (.A(_08669_),
    .B_N(net1009),
    .Y(_10998_));
 sg13g2_a21oi_1 _17790_ (.A1(net733),
    .A2(_10997_),
    .Y(_10999_),
    .B1(_10998_));
 sg13g2_buf_1 _17791_ (.A(_10999_),
    .X(_11000_));
 sg13g2_nand2_1 _17792_ (.Y(_11001_),
    .A(_10501_),
    .B(net606));
 sg13g2_or2_1 _17793_ (.X(_11002_),
    .B(_11001_),
    .A(net323));
 sg13g2_buf_1 _17794_ (.A(_10805_),
    .X(_11003_));
 sg13g2_nand2_1 _17795_ (.Y(_11004_),
    .A(_10801_),
    .B(net322));
 sg13g2_a21oi_1 _17796_ (.A1(_10807_),
    .A2(_10763_),
    .Y(_11005_),
    .B1(net1088));
 sg13g2_nand2_1 _17797_ (.Y(_11006_),
    .A(net606),
    .B(_11005_));
 sg13g2_inv_1 _17798_ (.Y(_11007_),
    .A(_10813_));
 sg13g2_nand4_1 _17799_ (.B(_10829_),
    .C(_10840_),
    .A(_10823_),
    .Y(_11008_),
    .D(_10843_));
 sg13g2_a221oi_1 _17800_ (.B2(_11008_),
    .C1(_10845_),
    .B1(_10106_),
    .A1(_09083_),
    .Y(_11009_),
    .A2(_10095_));
 sg13g2_buf_1 _17801_ (.A(_11009_),
    .X(_11010_));
 sg13g2_nor2_1 _17802_ (.A(_11007_),
    .B(_11010_),
    .Y(_11011_));
 sg13g2_or2_1 _17803_ (.X(_11012_),
    .B(_10916_),
    .A(_10887_));
 sg13g2_a21oi_1 _17804_ (.A1(net427),
    .A2(net426),
    .Y(_11013_),
    .B1(_11012_));
 sg13g2_o21ai_1 _17805_ (.B1(net341),
    .Y(_11014_),
    .A1(_11011_),
    .A2(_11013_));
 sg13g2_nor2_1 _17806_ (.A(_10851_),
    .B(_09205_),
    .Y(_11015_));
 sg13g2_a21oi_1 _17807_ (.A1(_11011_),
    .A2(_11013_),
    .Y(_11016_),
    .B1(net678));
 sg13g2_a21oi_1 _17808_ (.A1(_10851_),
    .A2(net341),
    .Y(_11017_),
    .B1(_10809_));
 sg13g2_a21o_1 _17809_ (.A2(net426),
    .A1(net427),
    .B1(_11012_),
    .X(_11018_));
 sg13g2_buf_1 _17810_ (.A(_11018_),
    .X(_11019_));
 sg13g2_a22oi_1 _17811_ (.Y(_11020_),
    .B1(_10813_),
    .B2(_10848_),
    .A2(_10881_),
    .A1(_10879_));
 sg13g2_buf_2 _17812_ (.A(_11020_),
    .X(_11021_));
 sg13g2_and2_1 _17813_ (.A(_11019_),
    .B(_11021_),
    .X(_11022_));
 sg13g2_a221oi_1 _17814_ (.B2(_11017_),
    .C1(_11022_),
    .B1(_11016_),
    .A1(_11014_),
    .Y(_11023_),
    .A2(_11015_));
 sg13g2_buf_1 _17815_ (.A(_11023_),
    .X(_11024_));
 sg13g2_a21oi_1 _17816_ (.A1(_11004_),
    .A2(_11006_),
    .Y(_11025_),
    .B1(_11024_));
 sg13g2_nor2_1 _17817_ (.A(_10807_),
    .B(net678),
    .Y(_11026_));
 sg13g2_nand2_1 _17818_ (.Y(_11027_),
    .A(net322),
    .B(_11026_));
 sg13g2_nor2_1 _17819_ (.A(net678),
    .B(net373),
    .Y(_11028_));
 sg13g2_a22oi_1 _17820_ (.Y(_11029_),
    .B1(_11028_),
    .B2(_11005_),
    .A2(_11026_),
    .A1(_10801_));
 sg13g2_o21ai_1 _17821_ (.B1(_11029_),
    .Y(_11030_),
    .A1(_11024_),
    .A2(_11027_));
 sg13g2_nor2_1 _17822_ (.A(_11025_),
    .B(_11030_),
    .Y(_11031_));
 sg13g2_a221oi_1 _17823_ (.B2(_11002_),
    .C1(_11031_),
    .B1(_10979_),
    .A1(net122),
    .Y(_11032_),
    .A2(_10949_));
 sg13g2_buf_1 _17824_ (.A(_11032_),
    .X(_11033_));
 sg13g2_a21o_1 _17825_ (.A2(_10971_),
    .A1(net1004),
    .B1(_10972_),
    .X(_11034_));
 sg13g2_nand2_1 _17826_ (.Y(_11035_),
    .A(net733),
    .B(_11034_));
 sg13g2_a21o_1 _17827_ (.A2(_10997_),
    .A1(_10165_),
    .B1(_10998_),
    .X(_11036_));
 sg13g2_buf_1 _17828_ (.A(_11036_),
    .X(_11037_));
 sg13g2_o21ai_1 _17829_ (.B1(net321),
    .Y(_11038_),
    .A1(_11025_),
    .A2(_11030_));
 sg13g2_a221oi_1 _17830_ (.B2(_11035_),
    .C1(_11038_),
    .B1(_10974_),
    .A1(net122),
    .Y(_11039_),
    .A2(_10949_));
 sg13g2_buf_1 _17831_ (.A(_11039_),
    .X(_11040_));
 sg13g2_a22oi_1 _17832_ (.Y(_11041_),
    .B1(net733),
    .B2(_11034_),
    .A2(net1009),
    .A1(_08679_));
 sg13g2_buf_1 _17833_ (.A(_11041_),
    .X(_11042_));
 sg13g2_or2_1 _17834_ (.X(_11043_),
    .B(_11001_),
    .A(_11042_));
 sg13g2_o21ai_1 _17835_ (.B1(_11043_),
    .Y(_11044_),
    .A1(_10979_),
    .A2(net323));
 sg13g2_buf_1 _17836_ (.A(_11044_),
    .X(_11045_));
 sg13g2_nor3_1 _17837_ (.A(_11033_),
    .B(_11040_),
    .C(_11045_),
    .Y(_11046_));
 sg13g2_buf_2 _17838_ (.A(_11046_),
    .X(_11047_));
 sg13g2_inv_1 _17839_ (.Y(_11048_),
    .A(\cpu.dec.imm[9] ));
 sg13g2_buf_1 _17840_ (.A(net541),
    .X(_11049_));
 sg13g2_buf_1 _17841_ (.A(net664),
    .X(_11050_));
 sg13g2_inv_1 _17842_ (.Y(_11051_),
    .A(_00267_));
 sg13g2_buf_1 _17843_ (.A(net755),
    .X(_11052_));
 sg13g2_mux4_1 _17844_ (.S0(net661),
    .A0(_11051_),
    .A1(\cpu.ex.r_13[9] ),
    .A2(\cpu.ex.r_11[9] ),
    .A3(\cpu.ex.r_9[9] ),
    .S1(_11052_),
    .X(_11053_));
 sg13g2_nor2b_1 _17845_ (.A(_11050_),
    .B_N(\cpu.ex.r_14[9] ),
    .Y(_11054_));
 sg13g2_a22oi_1 _17846_ (.Y(_11055_),
    .B1(_11054_),
    .B2(net736),
    .A2(_11053_),
    .A1(_11050_));
 sg13g2_buf_1 _17847_ (.A(net756),
    .X(_11056_));
 sg13g2_nor2b_1 _17848_ (.A(_11056_),
    .B_N(net664),
    .Y(_11057_));
 sg13g2_a22oi_1 _17849_ (.Y(_11058_),
    .B1(net736),
    .B2(\cpu.ex.r_mult[25] ),
    .A2(_10739_),
    .A1(\cpu.ex.r_lr[9] ));
 sg13g2_inv_1 _17850_ (.Y(_11059_),
    .A(_11058_));
 sg13g2_and2_1 _17851_ (.A(\cpu.ex.r_12[9] ),
    .B(_10826_),
    .X(_11060_));
 sg13g2_a21oi_1 _17852_ (.A1(\cpu.ex.r_8[9] ),
    .A2(_11052_),
    .Y(_11061_),
    .B1(_11060_));
 sg13g2_buf_1 _17853_ (.A(net757),
    .X(_11062_));
 sg13g2_nand3_1 _17854_ (.B(_11062_),
    .C(_10150_),
    .A(\cpu.ex.r_stmp[9] ),
    .Y(_11063_));
 sg13g2_o21ai_1 _17855_ (.B1(_11063_),
    .Y(_11064_),
    .A1(_10732_),
    .A2(_11061_));
 sg13g2_mux2_1 _17856_ (.A0(_10629_),
    .A1(\cpu.ex.r_10[9] ),
    .S(_11056_),
    .X(_11065_));
 sg13g2_a22oi_1 _17857_ (.Y(_11066_),
    .B1(_11065_),
    .B2(net662),
    .A2(_11057_),
    .A1(\cpu.ex.r_epc[9] ));
 sg13g2_nor2b_1 _17858_ (.A(_11066_),
    .B_N(_10857_),
    .Y(_11067_));
 sg13g2_a221oi_1 _17859_ (.B2(_10144_),
    .C1(_11067_),
    .B1(_11064_),
    .A1(_11057_),
    .Y(_11068_),
    .A2(_11059_));
 sg13g2_o21ai_1 _17860_ (.B1(_11068_),
    .Y(_11069_),
    .A1(net651),
    .A2(_11055_));
 sg13g2_a22oi_1 _17861_ (.Y(_11070_),
    .B1(net490),
    .B2(_11069_),
    .A2(net492),
    .A1(_10627_));
 sg13g2_mux2_1 _17862_ (.A0(_11048_),
    .A1(_11070_),
    .S(_10950_),
    .X(_11071_));
 sg13g2_a22oi_1 _17863_ (.Y(_11072_),
    .B1(_10980_),
    .B2(_11071_),
    .A2(net882),
    .A1(_08721_));
 sg13g2_buf_1 _17864_ (.A(_11072_),
    .X(_11073_));
 sg13g2_inv_1 _17865_ (.Y(_11074_),
    .A(\cpu.ex.pc[8] ));
 sg13g2_nand2_1 _17866_ (.Y(_11075_),
    .A(_11074_),
    .B(net882));
 sg13g2_mux2_1 _17867_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(\cpu.ex.r_mult[24] ),
    .S(_10120_),
    .X(_11076_));
 sg13g2_a22oi_1 _17868_ (.Y(_11077_),
    .B1(_11076_),
    .B2(_10132_),
    .A2(net735),
    .A1(_10697_));
 sg13g2_nand3_1 _17869_ (.B(net752),
    .C(net751),
    .A(\cpu.ex.r_10[8] ),
    .Y(_11078_));
 sg13g2_o21ai_1 _17870_ (.B1(_11078_),
    .Y(_11079_),
    .A1(net649),
    .A2(_11077_));
 sg13g2_a22oi_1 _17871_ (.Y(_11080_),
    .B1(_10113_),
    .B2(\cpu.ex.r_13[8] ),
    .A2(_10103_),
    .A1(\cpu.ex.r_lr[8] ));
 sg13g2_nand3_1 _17872_ (.B(net752),
    .C(_10147_),
    .A(\cpu.ex.r_8[8] ),
    .Y(_11081_));
 sg13g2_o21ai_1 _17873_ (.B1(_11081_),
    .Y(_11082_),
    .A1(net752),
    .A2(_11080_));
 sg13g2_mux2_1 _17874_ (.A0(_11079_),
    .A1(_11082_),
    .S(net661),
    .X(_11083_));
 sg13g2_mux2_1 _17875_ (.A0(_10704_),
    .A1(\cpu.ex.r_11[8] ),
    .S(net755),
    .X(_11084_));
 sg13g2_a221oi_1 _17876_ (.B2(_10133_),
    .C1(net661),
    .B1(_11084_),
    .A1(\cpu.ex.r_14[8] ),
    .Y(_11085_),
    .A2(_10778_));
 sg13g2_a221oi_1 _17877_ (.B2(\cpu.ex.r_12[8] ),
    .C1(_11062_),
    .B1(_10778_),
    .A1(\cpu.ex.r_9[8] ),
    .Y(_11086_),
    .A2(_10140_));
 sg13g2_nor3_1 _17878_ (.A(net651),
    .B(_11085_),
    .C(_11086_),
    .Y(_11087_));
 sg13g2_and4_1 _17879_ (.A(\cpu.ex.r_stmp[8] ),
    .B(_10144_),
    .C(_10859_),
    .D(net736),
    .X(_11088_));
 sg13g2_or3_1 _17880_ (.A(_11083_),
    .B(_11087_),
    .C(_11088_),
    .X(_11089_));
 sg13g2_a221oi_1 _17881_ (.B2(_11089_),
    .C1(net873),
    .B1(net541),
    .A1(_09011_),
    .Y(_11090_),
    .A2(net492));
 sg13g2_nor2_1 _17882_ (.A(_10161_),
    .B(\cpu.dec.imm[8] ),
    .Y(_11091_));
 sg13g2_o21ai_1 _17883_ (.B1(_10165_),
    .Y(_11092_),
    .A1(_11090_),
    .A2(_11091_));
 sg13g2_buf_1 _17884_ (.A(_11092_),
    .X(_11093_));
 sg13g2_nand2_1 _17885_ (.Y(_11094_),
    .A(_11075_),
    .B(_11093_));
 sg13g2_buf_1 _17886_ (.A(_11094_),
    .X(_11095_));
 sg13g2_nand2b_1 _17887_ (.Y(_11096_),
    .B(net211),
    .A_N(net212));
 sg13g2_buf_1 _17888_ (.A(_11096_),
    .X(_11097_));
 sg13g2_nand2b_1 _17889_ (.Y(_11098_),
    .B(_10076_),
    .A_N(_08710_));
 sg13g2_nand3_1 _17890_ (.B(net650),
    .C(net754),
    .A(\cpu.ex.r_9[10] ),
    .Y(_11099_));
 sg13g2_nand3_1 _17891_ (.B(net734),
    .C(net663),
    .A(_10072_),
    .Y(_11100_));
 sg13g2_a21oi_1 _17892_ (.A1(_11099_),
    .A2(_11100_),
    .Y(_11101_),
    .B1(net662));
 sg13g2_and2_1 _17893_ (.A(\cpu.ex.r_12[10] ),
    .B(_10729_),
    .X(_11102_));
 sg13g2_mux2_1 _17894_ (.A0(\cpu.ex.r_lr[10] ),
    .A1(\cpu.ex.r_epc[10] ),
    .S(net757),
    .X(_11103_));
 sg13g2_mux2_1 _17895_ (.A0(_10662_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net734),
    .X(_11104_));
 sg13g2_a22oi_1 _17896_ (.Y(_11105_),
    .B1(_11104_),
    .B2(_10748_),
    .A2(_11103_),
    .A1(net877));
 sg13g2_nor2_1 _17897_ (.A(net649),
    .B(_11105_),
    .Y(_11106_));
 sg13g2_nor2b_1 _17898_ (.A(_00268_),
    .B_N(net757),
    .Y(_11107_));
 sg13g2_nor2b_1 _17899_ (.A(net757),
    .B_N(\cpu.ex.r_13[10] ),
    .Y(_11108_));
 sg13g2_o21ai_1 _17900_ (.B1(net664),
    .Y(_11109_),
    .A1(_11107_),
    .A2(_11108_));
 sg13g2_a21oi_1 _17901_ (.A1(\cpu.ex.r_14[10] ),
    .A2(_10748_),
    .Y(_11110_),
    .B1(net755));
 sg13g2_mux2_1 _17902_ (.A0(\cpu.ex.r_8[10] ),
    .A1(\cpu.ex.r_10[10] ),
    .S(net757),
    .X(_11111_));
 sg13g2_a22oi_1 _17903_ (.Y(_11112_),
    .B1(_11111_),
    .B2(net752),
    .A2(_10108_),
    .A1(\cpu.ex.r_11[10] ));
 sg13g2_a221oi_1 _17904_ (.B2(net650),
    .C1(net651),
    .B1(_11112_),
    .A1(_11109_),
    .Y(_11113_),
    .A2(_11110_));
 sg13g2_or4_1 _17905_ (.A(_11101_),
    .B(_11102_),
    .C(_11106_),
    .D(_11113_),
    .X(_11114_));
 sg13g2_a221oi_1 _17906_ (.B2(_11114_),
    .C1(net873),
    .B1(net541),
    .A1(net1089),
    .Y(_11115_),
    .A2(_10095_));
 sg13g2_nor2_1 _17907_ (.A(net868),
    .B(\cpu.dec.imm[10] ),
    .Y(_11116_));
 sg13g2_o21ai_1 _17908_ (.B1(_10980_),
    .Y(_11117_),
    .A1(_11115_),
    .A2(_11116_));
 sg13g2_and2_1 _17909_ (.A(_11098_),
    .B(_11117_),
    .X(_11118_));
 sg13g2_buf_1 _17910_ (.A(_11118_),
    .X(_11119_));
 sg13g2_o21ai_1 _17911_ (.B1(net320),
    .Y(_11120_),
    .A1(_11047_),
    .A2(_11097_));
 sg13g2_buf_1 _17912_ (.A(net606),
    .X(_11121_));
 sg13g2_and2_1 _17913_ (.A(net539),
    .B(_10171_),
    .X(_11122_));
 sg13g2_buf_1 _17914_ (.A(_00302_),
    .X(_11123_));
 sg13g2_and2_1 _17915_ (.A(_11075_),
    .B(_11093_),
    .X(_11124_));
 sg13g2_buf_1 _17916_ (.A(_11124_),
    .X(_11125_));
 sg13g2_nand2_1 _17917_ (.Y(_11126_),
    .A(_11123_),
    .B(_11125_));
 sg13g2_nor4_1 _17918_ (.A(_11033_),
    .B(_11040_),
    .C(_11045_),
    .D(_11126_),
    .Y(_11127_));
 sg13g2_buf_1 _17919_ (.A(_00303_),
    .X(_11128_));
 sg13g2_nand2_1 _17920_ (.Y(_11129_),
    .A(net1087),
    .B(net212));
 sg13g2_nor4_1 _17921_ (.A(_11033_),
    .B(_11040_),
    .C(_11045_),
    .D(_11129_),
    .Y(_11130_));
 sg13g2_nand2_1 _17922_ (.Y(_11131_),
    .A(net212),
    .B(_11125_));
 sg13g2_nor4_1 _17923_ (.A(_11033_),
    .B(_11040_),
    .C(_11045_),
    .D(_11131_),
    .Y(_11132_));
 sg13g2_inv_1 _17924_ (.Y(_11133_),
    .A(_11123_));
 sg13g2_a21oi_1 _17925_ (.A1(_11123_),
    .A2(net212),
    .Y(_11134_),
    .B1(net1087));
 sg13g2_a21oi_1 _17926_ (.A1(_11133_),
    .A2(_11131_),
    .Y(_11135_),
    .B1(_11134_));
 sg13g2_nor4_2 _17927_ (.A(_11127_),
    .B(_11130_),
    .C(_11132_),
    .Y(_11136_),
    .D(_11135_));
 sg13g2_a22oi_1 _17928_ (.Y(_11137_),
    .B1(_11122_),
    .B2(_11136_),
    .A2(_11120_),
    .A1(_10171_));
 sg13g2_nand2_1 _17929_ (.Y(_11138_),
    .A(_10077_),
    .B(_10167_));
 sg13g2_buf_1 _17930_ (.A(_11138_),
    .X(_11139_));
 sg13g2_nand2_1 _17931_ (.Y(_11140_),
    .A(_10072_),
    .B(net606));
 sg13g2_nor2_1 _17932_ (.A(net320),
    .B(_11140_),
    .Y(_11141_));
 sg13g2_nor4_1 _17933_ (.A(_10073_),
    .B(_11047_),
    .C(_11097_),
    .D(net320),
    .Y(_11142_));
 sg13g2_a221oi_1 _17934_ (.B2(_11136_),
    .C1(_11142_),
    .B1(_11141_),
    .A1(_10072_),
    .Y(_11143_),
    .A2(net246));
 sg13g2_buf_1 _17935_ (.A(_11143_),
    .X(_11144_));
 sg13g2_nand2b_1 _17936_ (.Y(_11145_),
    .B(net882),
    .A_N(_08361_));
 sg13g2_nand3_1 _17937_ (.B(net650),
    .C(net754),
    .A(\cpu.ex.r_8[12] ),
    .Y(_11146_));
 sg13g2_nand3_1 _17938_ (.B(net734),
    .C(net663),
    .A(\cpu.ex.r_stmp[12] ),
    .Y(_11147_));
 sg13g2_a21oi_1 _17939_ (.A1(_11146_),
    .A2(_11147_),
    .Y(_11148_),
    .B1(net605));
 sg13g2_inv_1 _17940_ (.Y(_11149_),
    .A(net663));
 sg13g2_buf_1 _17941_ (.A(\cpu.ex.r_mult[28] ),
    .X(_11150_));
 sg13g2_a22oi_1 _17942_ (.Y(_11151_),
    .B1(_10901_),
    .B2(_11150_),
    .A2(net735),
    .A1(_10527_));
 sg13g2_nor2_1 _17943_ (.A(_11149_),
    .B(_11151_),
    .Y(_11152_));
 sg13g2_buf_1 _17944_ (.A(net734),
    .X(_11153_));
 sg13g2_mux2_1 _17945_ (.A0(_10541_),
    .A1(\cpu.ex.r_13[12] ),
    .S(net661),
    .X(_11154_));
 sg13g2_and3_1 _17946_ (.X(_11155_),
    .A(net647),
    .B(_11154_),
    .C(_10831_));
 sg13g2_nand3_1 _17947_ (.B(net758),
    .C(net665),
    .A(\cpu.ex.r_12[12] ),
    .Y(_11156_));
 sg13g2_mux2_1 _17948_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(\cpu.ex.r_epc[12] ),
    .S(net757),
    .X(_11157_));
 sg13g2_nand3_1 _17949_ (.B(net877),
    .C(_11157_),
    .A(net651),
    .Y(_11158_));
 sg13g2_nand2_1 _17950_ (.Y(_11159_),
    .A(_11156_),
    .B(_11158_));
 sg13g2_nor4_1 _17951_ (.A(_11148_),
    .B(_11152_),
    .C(_11155_),
    .D(_11159_),
    .Y(_11160_));
 sg13g2_nor2_1 _17952_ (.A(net664),
    .B(_10827_),
    .Y(_11161_));
 sg13g2_a221oi_1 _17953_ (.B2(\cpu.ex.r_14[12] ),
    .C1(net650),
    .B1(_11161_),
    .A1(_10525_),
    .Y(_11162_),
    .A2(_10819_));
 sg13g2_mux2_1 _17954_ (.A0(\cpu.ex.r_9[12] ),
    .A1(\cpu.ex.r_11[12] ),
    .S(net757),
    .X(_11163_));
 sg13g2_a22oi_1 _17955_ (.Y(_11164_),
    .B1(_11163_),
    .B2(net664),
    .A2(_10748_),
    .A1(\cpu.ex.r_10[12] ));
 sg13g2_o21ai_1 _17956_ (.B1(net650),
    .Y(_11165_),
    .A1(net651),
    .A2(_11164_));
 sg13g2_nand2b_1 _17957_ (.Y(_11166_),
    .B(_11165_),
    .A_N(_11162_));
 sg13g2_a21oi_1 _17958_ (.A1(_11160_),
    .A2(_11166_),
    .Y(_11167_),
    .B1(_10815_));
 sg13g2_nor3_1 _17959_ (.A(_08822_),
    .B(_10084_),
    .C(_10092_),
    .Y(_11168_));
 sg13g2_nor3_1 _17960_ (.A(net873),
    .B(_11167_),
    .C(_11168_),
    .Y(_11169_));
 sg13g2_nor2_1 _17961_ (.A(net868),
    .B(\cpu.dec.imm[12] ),
    .Y(_11170_));
 sg13g2_o21ai_1 _17962_ (.B1(net733),
    .Y(_11171_),
    .A1(_11169_),
    .A2(_11170_));
 sg13g2_nand2_1 _17963_ (.Y(_11172_),
    .A(_11145_),
    .B(_11171_));
 sg13g2_buf_2 _17964_ (.A(_11172_),
    .X(_11173_));
 sg13g2_buf_1 _17965_ (.A(_00300_),
    .X(_11174_));
 sg13g2_inv_1 _17966_ (.Y(_11175_),
    .A(_11174_));
 sg13g2_and2_1 _17967_ (.A(_11145_),
    .B(_11171_),
    .X(_11176_));
 sg13g2_buf_2 _17968_ (.A(_11176_),
    .X(_11177_));
 sg13g2_nor2_1 _17969_ (.A(_11174_),
    .B(net678),
    .Y(_11178_));
 sg13g2_nand2_1 _17970_ (.Y(_11179_),
    .A(_11177_),
    .B(_11178_));
 sg13g2_o21ai_1 _17971_ (.B1(_11179_),
    .Y(_11180_),
    .A1(_11175_),
    .A2(_11177_));
 sg13g2_buf_1 _17972_ (.A(_00299_),
    .X(_11181_));
 sg13g2_buf_1 _17973_ (.A(net492),
    .X(_11182_));
 sg13g2_a221oi_1 _17974_ (.B2(_10602_),
    .C1(net647),
    .B1(_10771_),
    .A1(\cpu.ex.r_11[15] ),
    .Y(_11183_),
    .A2(_10831_));
 sg13g2_a221oi_1 _17975_ (.B2(\cpu.ex.r_mult[31] ),
    .C1(net650),
    .B1(_11057_),
    .A1(\cpu.ex.r_14[15] ),
    .Y(_11184_),
    .A2(_10745_));
 sg13g2_nor3_1 _17976_ (.A(net661),
    .B(_11183_),
    .C(_11184_),
    .Y(_11185_));
 sg13g2_a22oi_1 _17977_ (.Y(_11186_),
    .B1(net665),
    .B2(\cpu.ex.r_13[15] ),
    .A2(_10103_),
    .A1(\cpu.ex.r_lr[15] ));
 sg13g2_nor2_1 _17978_ (.A(net662),
    .B(net648),
    .Y(_11187_));
 sg13g2_nor2b_1 _17979_ (.A(_11186_),
    .B_N(_11187_),
    .Y(_11188_));
 sg13g2_nand2_1 _17980_ (.Y(_11189_),
    .A(net649),
    .B(net650));
 sg13g2_a22oi_1 _17981_ (.Y(_11190_),
    .B1(_10748_),
    .B2(\cpu.ex.r_10[15] ),
    .A2(_11187_),
    .A1(\cpu.ex.r_9[15] ));
 sg13g2_nor2_1 _17982_ (.A(net648),
    .B(net649),
    .Y(_11191_));
 sg13g2_a22oi_1 _17983_ (.Y(_11192_),
    .B1(_11191_),
    .B2(_10614_),
    .A2(_10821_),
    .A1(\cpu.ex.r_15[15] ));
 sg13g2_nand2b_1 _17984_ (.Y(_11193_),
    .B(_10901_),
    .A_N(_11192_));
 sg13g2_o21ai_1 _17985_ (.B1(_11193_),
    .Y(_11194_),
    .A1(_11189_),
    .A2(_11190_));
 sg13g2_a22oi_1 _17986_ (.Y(_11195_),
    .B1(_10778_),
    .B2(\cpu.ex.r_stmp[15] ),
    .A2(net877),
    .A1(\cpu.ex.r_epc[15] ));
 sg13g2_mux2_1 _17987_ (.A0(\cpu.ex.r_8[15] ),
    .A1(\cpu.ex.r_12[15] ),
    .S(net647),
    .X(_11196_));
 sg13g2_nand3_1 _17988_ (.B(net758),
    .C(_11196_),
    .A(net649),
    .Y(_11197_));
 sg13g2_o21ai_1 _17989_ (.B1(_11197_),
    .Y(_11198_),
    .A1(_11149_),
    .A2(_11195_));
 sg13g2_or4_1 _17990_ (.A(_11185_),
    .B(_11188_),
    .C(_11194_),
    .D(_11198_),
    .X(_11199_));
 sg13g2_a22oi_1 _17991_ (.Y(_11200_),
    .B1(net490),
    .B2(_11199_),
    .A2(net425),
    .A1(net890));
 sg13g2_nor2_1 _17992_ (.A(net868),
    .B(\cpu.dec.imm[15] ),
    .Y(_11201_));
 sg13g2_a21oi_1 _17993_ (.A1(net868),
    .A2(_11200_),
    .Y(_11202_),
    .B1(_11201_));
 sg13g2_nand2_1 _17994_ (.Y(_11203_),
    .A(_08380_),
    .B(net882));
 sg13g2_o21ai_1 _17995_ (.B1(_11203_),
    .Y(_11204_),
    .A1(_10727_),
    .A2(_11202_));
 sg13g2_buf_1 _17996_ (.A(_11204_),
    .X(_11205_));
 sg13g2_buf_1 _17997_ (.A(_11205_),
    .X(_11206_));
 sg13g2_inv_1 _17998_ (.Y(_11207_),
    .A(net188));
 sg13g2_a221oi_1 _17999_ (.B2(_11181_),
    .C1(_11207_),
    .B1(_11180_),
    .A1(net616),
    .Y(_11208_),
    .A2(_11173_));
 sg13g2_xnor2_1 _18000_ (.Y(_11209_),
    .A(_11174_),
    .B(_11173_));
 sg13g2_nor2_1 _18001_ (.A(_11181_),
    .B(net678),
    .Y(_11210_));
 sg13g2_a21oi_1 _18002_ (.A1(_11209_),
    .A2(_11210_),
    .Y(_11211_),
    .B1(net188));
 sg13g2_nand3b_1 _18003_ (.B(net649),
    .C(\cpu.ex.r_12[14] ),
    .Y(_11212_),
    .A_N(net648));
 sg13g2_nand3b_1 _18004_ (.B(net648),
    .C(\cpu.ex.r_stmp[14] ),
    .Y(_11213_),
    .A_N(net649));
 sg13g2_a21oi_1 _18005_ (.A1(_11212_),
    .A2(_11213_),
    .Y(_11214_),
    .B1(net605));
 sg13g2_and3_1 _18006_ (.X(_11215_),
    .A(\cpu.ex.r_13[14] ),
    .B(net605),
    .C(net754));
 sg13g2_o21ai_1 _18007_ (.B1(net647),
    .Y(_11216_),
    .A1(_11214_),
    .A2(_11215_));
 sg13g2_mux2_1 _18008_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(\cpu.ex.r_mult[30] ),
    .S(net647),
    .X(_11217_));
 sg13g2_a22oi_1 _18009_ (.Y(_11218_),
    .B1(_11217_),
    .B2(net605),
    .A2(net735),
    .A1(_10554_));
 sg13g2_nand2b_1 _18010_ (.Y(_11219_),
    .B(net663),
    .A_N(_11218_));
 sg13g2_nand2b_1 _18011_ (.Y(_11220_),
    .B(net647),
    .A_N(_00272_));
 sg13g2_nand2b_1 _18012_ (.Y(_11221_),
    .B(\cpu.ex.r_11[14] ),
    .A_N(_11153_));
 sg13g2_a21oi_1 _18013_ (.A1(_11220_),
    .A2(_11221_),
    .Y(_11222_),
    .B1(_10827_));
 sg13g2_nand2_1 _18014_ (.Y(_11223_),
    .A(_10566_),
    .B(net647));
 sg13g2_nand2b_1 _18015_ (.Y(_11224_),
    .B(\cpu.ex.r_lr[14] ),
    .A_N(_11153_));
 sg13g2_a21oi_1 _18016_ (.A1(_11223_),
    .A2(_11224_),
    .Y(_11225_),
    .B1(_10818_));
 sg13g2_o21ai_1 _18017_ (.B1(net605),
    .Y(_11226_),
    .A1(_11222_),
    .A2(_11225_));
 sg13g2_nand3b_1 _18018_ (.B(net605),
    .C(\cpu.ex.r_9[14] ),
    .Y(_11227_),
    .A_N(net648));
 sg13g2_nand3b_1 _18019_ (.B(net648),
    .C(\cpu.ex.r_10[14] ),
    .Y(_11228_),
    .A_N(net605));
 sg13g2_nand2_1 _18020_ (.Y(_11229_),
    .A(_11227_),
    .B(_11228_));
 sg13g2_nand3_1 _18021_ (.B(net648),
    .C(net647),
    .A(\cpu.ex.r_14[14] ),
    .Y(_11230_));
 sg13g2_o21ai_1 _18022_ (.B1(_11230_),
    .Y(_11231_),
    .A1(_10560_),
    .A2(_10837_));
 sg13g2_a22oi_1 _18023_ (.Y(_11232_),
    .B1(_10745_),
    .B2(_11231_),
    .A2(_11229_),
    .A1(net751));
 sg13g2_nand4_1 _18024_ (.B(_11219_),
    .C(_11226_),
    .A(_11216_),
    .Y(_11233_),
    .D(_11232_));
 sg13g2_a22oi_1 _18025_ (.Y(_11234_),
    .B1(net490),
    .B2(_11233_),
    .A2(_11182_),
    .A1(net672));
 sg13g2_nand2_1 _18026_ (.Y(_11235_),
    .A(net868),
    .B(_11234_));
 sg13g2_o21ai_1 _18027_ (.B1(_11235_),
    .Y(_11236_),
    .A1(net868),
    .A2(\cpu.dec.imm[14] ));
 sg13g2_nor2b_1 _18028_ (.A(net1050),
    .B_N(net882),
    .Y(_11237_));
 sg13g2_a21o_1 _18029_ (.A2(net733),
    .A1(_11236_),
    .B1(_11237_),
    .X(_11238_));
 sg13g2_buf_2 _18030_ (.A(_11238_),
    .X(_11239_));
 sg13g2_inv_1 _18031_ (.Y(_11240_),
    .A(\cpu.dec.imm[13] ));
 sg13g2_nor2_1 _18032_ (.A(net662),
    .B(_10837_),
    .Y(_11241_));
 sg13g2_mux2_1 _18033_ (.A0(_10579_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net734),
    .X(_11242_));
 sg13g2_a22oi_1 _18034_ (.Y(_11243_),
    .B1(_10857_),
    .B2(\cpu.ex.r_epc[13] ),
    .A2(_10770_),
    .A1(_10594_));
 sg13g2_nor2_1 _18035_ (.A(net662),
    .B(_11243_),
    .Y(_11244_));
 sg13g2_a221oi_1 _18036_ (.B2(_10748_),
    .C1(_11244_),
    .B1(_11242_),
    .A1(\cpu.ex.r_lr[13] ),
    .Y(_11245_),
    .A2(_11241_));
 sg13g2_mux2_1 _18037_ (.A0(\cpu.ex.r_9[13] ),
    .A1(\cpu.ex.r_13[13] ),
    .S(net734),
    .X(_11246_));
 sg13g2_a22oi_1 _18038_ (.Y(_11247_),
    .B1(_11246_),
    .B2(net605),
    .A2(net735),
    .A1(\cpu.ex.r_8[13] ));
 sg13g2_inv_1 _18039_ (.Y(_11248_),
    .A(_11247_));
 sg13g2_inv_2 _18040_ (.Y(_11249_),
    .A(_10585_));
 sg13g2_mux2_1 _18041_ (.A0(_00271_),
    .A1(_11249_),
    .S(net651),
    .X(_11250_));
 sg13g2_nand2_1 _18042_ (.Y(_11251_),
    .A(\cpu.ex.r_14[13] ),
    .B(_10745_));
 sg13g2_o21ai_1 _18043_ (.B1(_11251_),
    .Y(_11252_),
    .A1(net662),
    .A2(_11250_));
 sg13g2_nand3_1 _18044_ (.B(net758),
    .C(net665),
    .A(\cpu.ex.r_12[13] ),
    .Y(_11253_));
 sg13g2_mux2_1 _18045_ (.A0(\cpu.ex.r_10[13] ),
    .A1(\cpu.ex.r_11[13] ),
    .S(net664),
    .X(_11254_));
 sg13g2_nand3_1 _18046_ (.B(net751),
    .C(_11254_),
    .A(net648),
    .Y(_11255_));
 sg13g2_nand2_1 _18047_ (.Y(_11256_),
    .A(_11253_),
    .B(_11255_));
 sg13g2_a221oi_1 _18048_ (.B2(_10742_),
    .C1(_11256_),
    .B1(_11252_),
    .A1(net754),
    .Y(_11257_),
    .A2(_11248_));
 sg13g2_o21ai_1 _18049_ (.B1(_11257_),
    .Y(_11258_),
    .A1(net649),
    .A2(_11245_));
 sg13g2_a22oi_1 _18050_ (.Y(_11259_),
    .B1(_11049_),
    .B2(_11258_),
    .A2(net492),
    .A1(net611));
 sg13g2_mux2_1 _18051_ (.A0(_11240_),
    .A1(_11259_),
    .S(net868),
    .X(_11260_));
 sg13g2_nor2b_1 _18052_ (.A(_08437_),
    .B_N(net882),
    .Y(_11261_));
 sg13g2_a21oi_1 _18053_ (.A1(net733),
    .A2(_11260_),
    .Y(_11262_),
    .B1(_11261_));
 sg13g2_buf_1 _18054_ (.A(_11262_),
    .X(_11263_));
 sg13g2_nor2_1 _18055_ (.A(_11239_),
    .B(_11263_),
    .Y(_11264_));
 sg13g2_nand2_1 _18056_ (.Y(_11265_),
    .A(_10585_),
    .B(_11264_));
 sg13g2_xnor2_1 _18057_ (.Y(_11266_),
    .A(_11249_),
    .B(_11239_));
 sg13g2_nand3_1 _18058_ (.B(_11263_),
    .C(_11266_),
    .A(net1086),
    .Y(_11267_));
 sg13g2_o21ai_1 _18059_ (.B1(_11267_),
    .Y(_11268_),
    .A1(net1086),
    .A2(_11265_));
 sg13g2_a21oi_1 _18060_ (.A1(_11236_),
    .A2(net733),
    .Y(_11269_),
    .B1(_11237_));
 sg13g2_buf_1 _18061_ (.A(_11269_),
    .X(_11270_));
 sg13g2_buf_1 _18062_ (.A(_11263_),
    .X(_11271_));
 sg13g2_nor2_1 _18063_ (.A(_11270_),
    .B(net187),
    .Y(_11272_));
 sg13g2_o21ai_1 _18064_ (.B1(_10725_),
    .Y(_11273_),
    .A1(net1086),
    .A2(_10585_));
 sg13g2_a22oi_1 _18065_ (.Y(_11274_),
    .B1(_11272_),
    .B2(_11273_),
    .A2(_11268_),
    .A1(net606));
 sg13g2_or3_1 _18066_ (.A(_11208_),
    .B(_11211_),
    .C(_11274_),
    .X(_11275_));
 sg13g2_buf_1 _18067_ (.A(_11275_),
    .X(_11276_));
 sg13g2_nand2b_1 _18068_ (.Y(_11277_),
    .B(net539),
    .A_N(_11276_));
 sg13g2_a21oi_1 _18069_ (.A1(_11137_),
    .A2(_11144_),
    .Y(_11278_),
    .B1(_11277_));
 sg13g2_buf_8 _18070_ (.A(_11278_),
    .X(_11279_));
 sg13g2_nand2_1 _18071_ (.Y(_11280_),
    .A(net539),
    .B(_11134_));
 sg13g2_a21o_1 _18072_ (.A2(_11280_),
    .A1(_11097_),
    .B1(_11047_),
    .X(_11281_));
 sg13g2_or3_1 _18073_ (.A(_11033_),
    .B(_11040_),
    .C(_11045_),
    .X(_11282_));
 sg13g2_nor2_1 _18074_ (.A(_11123_),
    .B(_09212_),
    .Y(_11283_));
 sg13g2_inv_1 _18075_ (.Y(_11284_),
    .A(_11283_));
 sg13g2_nor2_1 _18076_ (.A(_11125_),
    .B(_11284_),
    .Y(_11285_));
 sg13g2_buf_1 _18077_ (.A(net212),
    .X(_11286_));
 sg13g2_nand3_1 _18078_ (.B(net211),
    .C(_11134_),
    .A(net606),
    .Y(_11287_));
 sg13g2_o21ai_1 _18079_ (.B1(_11287_),
    .Y(_11288_),
    .A1(net186),
    .A2(_11284_));
 sg13g2_a21oi_1 _18080_ (.A1(_11282_),
    .A2(_11285_),
    .Y(_11289_),
    .B1(_11288_));
 sg13g2_nand2_1 _18081_ (.Y(_11290_),
    .A(_11098_),
    .B(_11117_));
 sg13g2_buf_1 _18082_ (.A(_11290_),
    .X(_11291_));
 sg13g2_nand2_1 _18083_ (.Y(_11292_),
    .A(net246),
    .B(net319));
 sg13g2_a21o_1 _18084_ (.A2(_11289_),
    .A1(_11281_),
    .B1(_11292_),
    .X(_11293_));
 sg13g2_a21o_1 _18085_ (.A2(_11260_),
    .A1(net733),
    .B1(_11261_),
    .X(_11294_));
 sg13g2_buf_2 _18086_ (.A(_11294_),
    .X(_11295_));
 sg13g2_a21oi_1 _18087_ (.A1(_11145_),
    .A2(_11171_),
    .Y(_11296_),
    .B1(_11174_));
 sg13g2_o21ai_1 _18088_ (.B1(net1086),
    .Y(_11297_),
    .A1(net210),
    .A2(_11296_));
 sg13g2_nand2_1 _18089_ (.Y(_11298_),
    .A(net210),
    .B(_11296_));
 sg13g2_a21oi_1 _18090_ (.A1(_11297_),
    .A2(_11298_),
    .Y(_11299_),
    .B1(net678));
 sg13g2_nor2_1 _18091_ (.A(_11239_),
    .B(_11299_),
    .Y(_11300_));
 sg13g2_a21o_1 _18092_ (.A2(_11207_),
    .A1(_11181_),
    .B1(_11249_),
    .X(_11301_));
 sg13g2_nand2_1 _18093_ (.Y(_11302_),
    .A(_11239_),
    .B(_11299_));
 sg13g2_a21o_1 _18094_ (.A2(_11302_),
    .A1(_11207_),
    .B1(_11181_),
    .X(_11303_));
 sg13g2_o21ai_1 _18095_ (.B1(_11303_),
    .Y(_11304_),
    .A1(_11300_),
    .A2(_11301_));
 sg13g2_nor2_1 _18096_ (.A(_11207_),
    .B(_11302_),
    .Y(_11305_));
 sg13g2_a21oi_1 _18097_ (.A1(net539),
    .A2(_11304_),
    .Y(_11306_),
    .B1(_11305_));
 sg13g2_o21ai_1 _18098_ (.B1(_11306_),
    .Y(_11307_),
    .A1(_11276_),
    .A2(_11293_));
 sg13g2_buf_2 _18099_ (.A(_11307_),
    .X(_11308_));
 sg13g2_nor2_1 _18100_ (.A(_09209_),
    .B(net678),
    .Y(_11309_));
 sg13g2_nor2_1 _18101_ (.A(_11004_),
    .B(net323),
    .Y(_11310_));
 sg13g2_nand3_1 _18102_ (.B(net188),
    .C(_11310_),
    .A(_11173_),
    .Y(_11311_));
 sg13g2_nand2_1 _18103_ (.Y(_11312_),
    .A(_10879_),
    .B(_10881_));
 sg13g2_buf_1 _18104_ (.A(_11312_),
    .X(_11313_));
 sg13g2_nand2_1 _18105_ (.Y(_11314_),
    .A(net340),
    .B(_10850_));
 sg13g2_buf_2 _18106_ (.A(_11314_),
    .X(_11315_));
 sg13g2_buf_1 _18107_ (.A(_10947_),
    .X(_11316_));
 sg13g2_nand2_1 _18108_ (.Y(_11317_),
    .A(_10918_),
    .B(net245));
 sg13g2_buf_1 _18109_ (.A(_11317_),
    .X(_11318_));
 sg13g2_nor2_2 _18110_ (.A(_11315_),
    .B(net185),
    .Y(_11319_));
 sg13g2_nand4_1 _18111_ (.B(net210),
    .C(_10976_),
    .A(_11239_),
    .Y(_11320_),
    .D(_11319_));
 sg13g2_nor4_1 _18112_ (.A(_11097_),
    .B(_11292_),
    .C(_11311_),
    .D(_11320_),
    .Y(_11321_));
 sg13g2_nor3_1 _18113_ (.A(_11309_),
    .B(_09221_),
    .C(_11321_),
    .Y(_11322_));
 sg13g2_buf_1 _18114_ (.A(_11322_),
    .X(_11323_));
 sg13g2_buf_1 _18115_ (.A(_11323_),
    .X(_11324_));
 sg13g2_o21ai_1 _18116_ (.B1(net77),
    .Y(_11325_),
    .A1(_11279_),
    .A2(_11308_));
 sg13g2_nor3_1 _18117_ (.A(_10524_),
    .B(_10650_),
    .C(_10720_),
    .Y(_11326_));
 sg13g2_buf_1 _18118_ (.A(_11326_),
    .X(_11327_));
 sg13g2_buf_1 _18119_ (.A(_11327_),
    .X(_11328_));
 sg13g2_buf_1 _18120_ (.A(_11328_),
    .X(_11329_));
 sg13g2_nand2_1 _18121_ (.Y(_11330_),
    .A(_10925_),
    .B(_10945_));
 sg13g2_buf_2 _18122_ (.A(_11330_),
    .X(_11331_));
 sg13g2_buf_1 _18123_ (.A(_11331_),
    .X(_11332_));
 sg13g2_nand3_1 _18124_ (.B(net88),
    .C(net244),
    .A(_09221_),
    .Y(_11333_));
 sg13g2_nand2_1 _18125_ (.Y(_11334_),
    .A(_10061_),
    .B(_10064_));
 sg13g2_buf_1 _18126_ (.A(_11334_),
    .X(_11335_));
 sg13g2_a21oi_1 _18127_ (.A1(_11325_),
    .A2(_11333_),
    .Y(_11336_),
    .B1(net538));
 sg13g2_a21o_1 _18128_ (.A2(net374),
    .A1(_10050_),
    .B1(_11336_),
    .X(\cpu.ex.c_mult[0] ));
 sg13g2_buf_1 _18129_ (.A(\cpu.dec.load ),
    .X(_11337_));
 sg13g2_nand2_1 _18130_ (.Y(_11338_),
    .A(_08734_),
    .B(_09028_));
 sg13g2_nor2_1 _18131_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11339_));
 sg13g2_nand2_1 _18132_ (.Y(_11340_),
    .A(\cpu.dec.iready ),
    .B(_00199_));
 sg13g2_nor2_1 _18133_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11340_),
    .Y(_11341_));
 sg13g2_buf_1 _18134_ (.A(_11341_),
    .X(_11342_));
 sg13g2_nand2_1 _18135_ (.Y(_11343_),
    .A(_09126_),
    .B(_11342_));
 sg13g2_nor2_1 _18136_ (.A(net1111),
    .B(_11343_),
    .Y(_11344_));
 sg13g2_buf_1 _18137_ (.A(_00258_),
    .X(_11345_));
 sg13g2_nand2_1 _18138_ (.Y(_11346_),
    .A(_10176_),
    .B(\cpu.cond[2] ));
 sg13g2_a21o_1 _18139_ (.A2(_11346_),
    .A1(_11345_),
    .B1(net1033),
    .X(_11347_));
 sg13g2_buf_1 _18140_ (.A(_11347_),
    .X(_11348_));
 sg13g2_o21ai_1 _18141_ (.B1(_11348_),
    .Y(_11349_),
    .A1(_10176_),
    .A2(\cpu.dec.jmp ));
 sg13g2_nand2_1 _18142_ (.Y(_11350_),
    .A(_11344_),
    .B(_11349_));
 sg13g2_a21oi_1 _18143_ (.A1(_10343_),
    .A2(\cpu.dec.r_swapsp ),
    .Y(_11351_),
    .B1(_11350_));
 sg13g2_nor2_1 _18144_ (.A(net1030),
    .B(_09211_),
    .Y(_11352_));
 sg13g2_nor2_1 _18145_ (.A(_10067_),
    .B(_11352_),
    .Y(_11353_));
 sg13g2_buf_2 _18146_ (.A(_11353_),
    .X(_11354_));
 sg13g2_a21oi_1 _18147_ (.A1(_11339_),
    .A2(_11351_),
    .Y(_11355_),
    .B1(_11354_));
 sg13g2_a21oi_1 _18148_ (.A1(_11338_),
    .A2(_11355_),
    .Y(_11356_),
    .B1(net1030));
 sg13g2_buf_2 _18149_ (.A(_11356_),
    .X(_11357_));
 sg13g2_nand2_1 _18150_ (.Y(_11358_),
    .A(_00310_),
    .B(_11357_));
 sg13g2_a21o_1 _18151_ (.A2(_11355_),
    .A1(_11338_),
    .B1(net896),
    .X(_11359_));
 sg13g2_buf_1 _18152_ (.A(_11359_),
    .X(_11360_));
 sg13g2_and2_1 _18153_ (.A(net886),
    .B(_09078_),
    .X(_11361_));
 sg13g2_nand2_1 _18154_ (.Y(_11362_),
    .A(_09651_),
    .B(_09653_));
 sg13g2_a21oi_2 _18155_ (.B1(_09103_),
    .Y(_11363_),
    .A2(_11362_),
    .A1(_11361_));
 sg13g2_nand2_1 _18156_ (.Y(_11364_),
    .A(_11360_),
    .B(_11363_));
 sg13g2_a21o_1 _18157_ (.A2(_11364_),
    .A1(_11358_),
    .B1(_08766_),
    .X(_11365_));
 sg13g2_o21ai_1 _18158_ (.B1(_11365_),
    .Y(_00054_),
    .A1(_11337_),
    .A2(_11358_));
 sg13g2_buf_1 _18159_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11366_));
 sg13g2_inv_1 _18160_ (.Y(_11367_),
    .A(_10050_));
 sg13g2_buf_1 _18161_ (.A(_10918_),
    .X(_11368_));
 sg13g2_buf_1 _18162_ (.A(_10722_),
    .X(_11369_));
 sg13g2_nor2_1 _18163_ (.A(net318),
    .B(net99),
    .Y(_11370_));
 sg13g2_buf_1 _18164_ (.A(_09201_),
    .X(_11371_));
 sg13g2_buf_1 _18165_ (.A(net732),
    .X(_11372_));
 sg13g2_buf_1 _18166_ (.A(net646),
    .X(_11373_));
 sg13g2_nor3_1 _18167_ (.A(_11367_),
    .B(_11373_),
    .C(_11370_),
    .Y(_11374_));
 sg13g2_a21oi_1 _18168_ (.A1(_11367_),
    .A2(_11370_),
    .Y(_11375_),
    .B1(_11374_));
 sg13g2_a22oi_1 _18169_ (.Y(_11376_),
    .B1(_11370_),
    .B2(_11373_),
    .A2(net89),
    .A1(_10050_));
 sg13g2_o21ai_1 _18170_ (.B1(_11376_),
    .Y(_11377_),
    .A1(_09216_),
    .A2(_11375_));
 sg13g2_a22oi_1 _18171_ (.Y(_11378_),
    .B1(_11377_),
    .B2(net542),
    .A2(net374),
    .A1(_11366_));
 sg13g2_inv_1 _18172_ (.Y(\cpu.ex.c_mult[1] ),
    .A(_11378_));
 sg13g2_a221oi_1 _18173_ (.B2(net426),
    .C1(_11367_),
    .B1(net427),
    .A1(net1056),
    .Y(_11379_),
    .A2(_10075_));
 sg13g2_buf_1 _18174_ (.A(_11379_),
    .X(_11380_));
 sg13g2_inv_1 _18175_ (.Y(_11381_),
    .A(_11366_));
 sg13g2_o21ai_1 _18176_ (.B1(_11381_),
    .Y(_11382_),
    .A1(_11007_),
    .A2(_11010_));
 sg13g2_buf_1 _18177_ (.A(_11011_),
    .X(_11383_));
 sg13g2_nand2_1 _18178_ (.Y(_11384_),
    .A(_11366_),
    .B(net317));
 sg13g2_o21ai_1 _18179_ (.B1(_11384_),
    .Y(_11385_),
    .A1(net99),
    .A2(_11382_));
 sg13g2_o21ai_1 _18180_ (.B1(net100),
    .Y(_11386_),
    .A1(net317),
    .A2(_11380_));
 sg13g2_a22oi_1 _18181_ (.Y(_11387_),
    .B1(_11386_),
    .B2(_11366_),
    .A2(_11385_),
    .A1(_11380_));
 sg13g2_a21oi_1 _18182_ (.A1(_10891_),
    .A2(_10915_),
    .Y(_11388_),
    .B1(_10916_));
 sg13g2_buf_8 _18183_ (.A(_11388_),
    .X(_11389_));
 sg13g2_nand2_1 _18184_ (.Y(_11390_),
    .A(_10050_),
    .B(net339));
 sg13g2_nand4_1 _18185_ (.B(net317),
    .C(net100),
    .A(_11381_),
    .Y(_11391_),
    .D(_11390_));
 sg13g2_o21ai_1 _18186_ (.B1(_11391_),
    .Y(_11392_),
    .A1(net604),
    .A2(_11387_));
 sg13g2_buf_1 _18187_ (.A(_10850_),
    .X(_11393_));
 sg13g2_buf_1 _18188_ (.A(_11369_),
    .X(_11394_));
 sg13g2_nor3_1 _18189_ (.A(net677),
    .B(net209),
    .C(net87),
    .Y(_11395_));
 sg13g2_a221oi_1 _18190_ (.B2(net1103),
    .C1(_11395_),
    .B1(_11392_),
    .A1(_11366_),
    .Y(_11396_),
    .A2(net89));
 sg13g2_nand2_1 _18191_ (.Y(_11397_),
    .A(\cpu.ex.r_mult[2] ),
    .B(net428));
 sg13g2_o21ai_1 _18192_ (.B1(_11397_),
    .Y(\cpu.ex.c_mult[2] ),
    .A1(net538),
    .A2(_11396_));
 sg13g2_buf_1 _18193_ (.A(_00120_),
    .X(_11398_));
 sg13g2_inv_1 _18194_ (.Y(_11399_),
    .A(_11398_));
 sg13g2_a21oi_1 _18195_ (.A1(_11011_),
    .A2(_11380_),
    .Y(_11400_),
    .B1(_11366_));
 sg13g2_a21oi_1 _18196_ (.A1(net209),
    .A2(_11390_),
    .Y(_11401_),
    .B1(_11400_));
 sg13g2_buf_1 _18197_ (.A(net340),
    .X(_11402_));
 sg13g2_nand2_1 _18198_ (.Y(_11403_),
    .A(_11398_),
    .B(net316));
 sg13g2_nand2_1 _18199_ (.Y(_11404_),
    .A(_11399_),
    .B(net341));
 sg13g2_o21ai_1 _18200_ (.B1(_11404_),
    .Y(_11405_),
    .A1(net122),
    .A2(_11403_));
 sg13g2_nor2_1 _18201_ (.A(_11398_),
    .B(net100),
    .Y(_11406_));
 sg13g2_a21o_1 _18202_ (.A2(_11405_),
    .A1(_11401_),
    .B1(_11406_),
    .X(_11407_));
 sg13g2_nor2_1 _18203_ (.A(_11399_),
    .B(_11402_),
    .Y(_11408_));
 sg13g2_nor2_1 _18204_ (.A(_11398_),
    .B(_09201_),
    .Y(_11409_));
 sg13g2_a22oi_1 _18205_ (.Y(_11410_),
    .B1(_11409_),
    .B2(net316),
    .A2(_11408_),
    .A1(net100));
 sg13g2_nor2_1 _18206_ (.A(_11401_),
    .B(_11410_),
    .Y(_11411_));
 sg13g2_a21o_1 _18207_ (.A2(_11407_),
    .A1(net677),
    .B1(_11411_),
    .X(_11412_));
 sg13g2_nor3_1 _18208_ (.A(net677),
    .B(net316),
    .C(net87),
    .Y(_11413_));
 sg13g2_a221oi_1 _18209_ (.B2(net1103),
    .C1(_11413_),
    .B1(_11412_),
    .A1(_11399_),
    .Y(_11414_),
    .A2(net89));
 sg13g2_nand2_1 _18210_ (.Y(_11415_),
    .A(\cpu.ex.r_mult[3] ),
    .B(net428));
 sg13g2_o21ai_1 _18211_ (.B1(_11415_),
    .Y(\cpu.ex.c_mult[3] ),
    .A1(net538),
    .A2(_11414_));
 sg13g2_buf_1 _18212_ (.A(_00127_),
    .X(_11416_));
 sg13g2_inv_1 _18213_ (.Y(_11417_),
    .A(_11416_));
 sg13g2_nor2_1 _18214_ (.A(_11416_),
    .B(net646),
    .Y(_11418_));
 sg13g2_nor3_1 _18215_ (.A(_11381_),
    .B(_11007_),
    .C(_11010_),
    .Y(_11419_));
 sg13g2_o21ai_1 _18216_ (.B1(_11382_),
    .Y(_11420_),
    .A1(_11380_),
    .A2(_11419_));
 sg13g2_a21oi_1 _18217_ (.A1(net340),
    .A2(_11420_),
    .Y(_11421_),
    .B1(_11398_));
 sg13g2_nor2_1 _18218_ (.A(net340),
    .B(_11420_),
    .Y(_11422_));
 sg13g2_o21ai_1 _18219_ (.B1(net677),
    .Y(_11423_),
    .A1(_11421_),
    .A2(_11422_));
 sg13g2_xnor2_1 _18220_ (.Y(_11424_),
    .A(net373),
    .B(_11423_));
 sg13g2_nand2_1 _18221_ (.Y(_11425_),
    .A(_11327_),
    .B(_11424_));
 sg13g2_mux2_1 _18222_ (.A0(_11416_),
    .A1(_11418_),
    .S(_11425_),
    .X(_11426_));
 sg13g2_nor2_1 _18223_ (.A(net677),
    .B(_11425_),
    .Y(_11427_));
 sg13g2_a221oi_1 _18224_ (.B2(net1103),
    .C1(_11427_),
    .B1(_11426_),
    .A1(_11417_),
    .Y(_11428_),
    .A2(net89));
 sg13g2_nand2_1 _18225_ (.Y(_11429_),
    .A(\cpu.ex.r_mult[4] ),
    .B(net428));
 sg13g2_o21ai_1 _18226_ (.B1(_11429_),
    .Y(\cpu.ex.c_mult[4] ),
    .A1(net538),
    .A2(_11428_));
 sg13g2_nand2_1 _18227_ (.Y(_11430_),
    .A(_11417_),
    .B(net373));
 sg13g2_inv_1 _18228_ (.Y(_11431_),
    .A(_11430_));
 sg13g2_nand2b_1 _18229_ (.Y(_11432_),
    .B(_11416_),
    .A_N(net373));
 sg13g2_nand3_1 _18230_ (.B(net341),
    .C(_11432_),
    .A(_09218_),
    .Y(_11433_));
 sg13g2_nand2_1 _18231_ (.Y(_11434_),
    .A(_11409_),
    .B(_11432_));
 sg13g2_a221oi_1 _18232_ (.B2(_11434_),
    .C1(_11400_),
    .B1(_11433_),
    .A1(_10850_),
    .Y(_11435_),
    .A2(_11390_));
 sg13g2_buf_2 _18233_ (.A(_11435_),
    .X(_11436_));
 sg13g2_nor2b_2 _18234_ (.A(_11404_),
    .B_N(_11432_),
    .Y(_11437_));
 sg13g2_nor3_2 _18235_ (.A(_11431_),
    .B(_11436_),
    .C(_11437_),
    .Y(_11438_));
 sg13g2_buf_1 _18236_ (.A(_00139_),
    .X(_11439_));
 sg13g2_buf_1 _18237_ (.A(_10801_),
    .X(_11440_));
 sg13g2_nand2_1 _18238_ (.Y(_11441_),
    .A(net677),
    .B(net243));
 sg13g2_buf_1 _18239_ (.A(_10763_),
    .X(_11442_));
 sg13g2_nand3_1 _18240_ (.B(net242),
    .C(net100),
    .A(_11439_),
    .Y(_11443_));
 sg13g2_o21ai_1 _18241_ (.B1(_11443_),
    .Y(_11444_),
    .A1(_11439_),
    .A2(_11441_));
 sg13g2_inv_1 _18242_ (.Y(_11445_),
    .A(_11439_));
 sg13g2_nor2_1 _18243_ (.A(_11445_),
    .B(_10763_),
    .Y(_11446_));
 sg13g2_nor2_1 _18244_ (.A(_11439_),
    .B(net243),
    .Y(_11447_));
 sg13g2_a21oi_1 _18245_ (.A1(net100),
    .A2(_11446_),
    .Y(_11448_),
    .B1(_11447_));
 sg13g2_nand2_1 _18246_ (.Y(_11449_),
    .A(_11445_),
    .B(net99));
 sg13g2_o21ai_1 _18247_ (.B1(_11449_),
    .Y(_11450_),
    .A1(_11438_),
    .A2(_11448_));
 sg13g2_a22oi_1 _18248_ (.Y(_11451_),
    .B1(_11450_),
    .B2(_09219_),
    .A2(_11444_),
    .A1(_11438_));
 sg13g2_nor2_1 _18249_ (.A(_09219_),
    .B(net99),
    .Y(_11452_));
 sg13g2_a22oi_1 _18250_ (.Y(_11453_),
    .B1(_11452_),
    .B2(net242),
    .A2(net89),
    .A1(_11445_));
 sg13g2_o21ai_1 _18251_ (.B1(_11453_),
    .Y(_11454_),
    .A1(_09216_),
    .A2(_11451_));
 sg13g2_a22oi_1 _18252_ (.Y(_11455_),
    .B1(_11454_),
    .B2(net542),
    .A2(net374),
    .A1(\cpu.ex.r_mult[5] ));
 sg13g2_inv_1 _18253_ (.Y(\cpu.ex.c_mult[5] ),
    .A(_11455_));
 sg13g2_buf_1 _18254_ (.A(_00151_),
    .X(_11456_));
 sg13g2_inv_1 _18255_ (.Y(_11457_),
    .A(_11456_));
 sg13g2_nand2_1 _18256_ (.Y(_11458_),
    .A(_11457_),
    .B(net77));
 sg13g2_a21o_1 _18257_ (.A2(_11438_),
    .A1(_11440_),
    .B1(_11439_),
    .X(_11459_));
 sg13g2_or2_1 _18258_ (.X(_11460_),
    .B(_11438_),
    .A(_11440_));
 sg13g2_a21o_1 _18259_ (.A2(_11460_),
    .A1(_11459_),
    .B1(net646),
    .X(_11461_));
 sg13g2_xnor2_1 _18260_ (.Y(_11462_),
    .A(net323),
    .B(_11461_));
 sg13g2_nor2_1 _18261_ (.A(_11456_),
    .B(net646),
    .Y(_11463_));
 sg13g2_inv_1 _18262_ (.Y(_11464_),
    .A(_11463_));
 sg13g2_a21oi_1 _18263_ (.A1(net88),
    .A2(_11462_),
    .Y(_11465_),
    .B1(_11464_));
 sg13g2_and3_1 _18264_ (.X(_11466_),
    .A(net88),
    .B(_11462_),
    .C(_11464_));
 sg13g2_o21ai_1 _18265_ (.B1(_09221_),
    .Y(_11467_),
    .A1(_11465_),
    .A2(_11466_));
 sg13g2_a21oi_1 _18266_ (.A1(_11458_),
    .A2(_11467_),
    .Y(_11468_),
    .B1(net538));
 sg13g2_a21o_1 _18267_ (.A2(net374),
    .A1(\cpu.ex.r_mult[6] ),
    .B1(_11468_),
    .X(\cpu.ex.c_mult[6] ));
 sg13g2_inv_1 _18268_ (.Y(_11469_),
    .A(_00163_));
 sg13g2_nor2_1 _18269_ (.A(_11456_),
    .B(net321),
    .Y(_11470_));
 sg13g2_nand2_1 _18270_ (.Y(_11471_),
    .A(_10801_),
    .B(_11430_));
 sg13g2_nor4_2 _18271_ (.A(_11436_),
    .B(_11437_),
    .C(_11470_),
    .Y(_11472_),
    .D(_11471_));
 sg13g2_nand2_1 _18272_ (.Y(_11473_),
    .A(_11439_),
    .B(_11430_));
 sg13g2_nor4_2 _18273_ (.A(_11436_),
    .B(_11437_),
    .C(_11470_),
    .Y(_11474_),
    .D(_11473_));
 sg13g2_o21ai_1 _18274_ (.B1(_11446_),
    .Y(_11475_),
    .A1(_11456_),
    .A2(_11037_));
 sg13g2_o21ai_1 _18275_ (.B1(_11475_),
    .Y(_11476_),
    .A1(_11457_),
    .A2(_10999_));
 sg13g2_buf_1 _18276_ (.A(_11476_),
    .X(_11477_));
 sg13g2_nor4_1 _18277_ (.A(net646),
    .B(_11472_),
    .C(_11474_),
    .D(_11477_),
    .Y(_11478_));
 sg13g2_xnor2_1 _18278_ (.Y(_11479_),
    .A(_10976_),
    .B(_11478_));
 sg13g2_nand2_1 _18279_ (.Y(_11480_),
    .A(net100),
    .B(_11479_));
 sg13g2_nor2_2 _18280_ (.A(_00163_),
    .B(net732),
    .Y(_11481_));
 sg13g2_xnor2_1 _18281_ (.Y(_11482_),
    .A(_11480_),
    .B(_11481_));
 sg13g2_a22oi_1 _18282_ (.Y(_11483_),
    .B1(_11482_),
    .B2(_09221_),
    .A2(net89),
    .A1(_11469_));
 sg13g2_nand2_1 _18283_ (.Y(_11484_),
    .A(\cpu.ex.r_mult[7] ),
    .B(_10070_));
 sg13g2_o21ai_1 _18284_ (.B1(_11484_),
    .Y(\cpu.ex.c_mult[7] ),
    .A1(net538),
    .A2(_11483_));
 sg13g2_nand2b_1 _18285_ (.Y(_11485_),
    .B(_11463_),
    .A_N(_11461_));
 sg13g2_a221oi_1 _18286_ (.B2(_11460_),
    .C1(net122),
    .B1(_11459_),
    .A1(_09197_),
    .Y(_11486_),
    .A2(_10723_));
 sg13g2_o21ai_1 _18287_ (.B1(_11000_),
    .Y(_11487_),
    .A1(_11463_),
    .A2(_11486_));
 sg13g2_buf_1 _18288_ (.A(_11042_),
    .X(_11488_));
 sg13g2_nor2_1 _18289_ (.A(net184),
    .B(_11481_),
    .Y(_11489_));
 sg13g2_a21o_1 _18290_ (.A2(_11487_),
    .A1(_11485_),
    .B1(_11489_),
    .X(_11490_));
 sg13g2_nand2_1 _18291_ (.Y(_11491_),
    .A(net184),
    .B(_11481_));
 sg13g2_and2_1 _18292_ (.A(_09221_),
    .B(net542),
    .X(_11492_));
 sg13g2_buf_1 _18293_ (.A(_11492_),
    .X(_11493_));
 sg13g2_inv_1 _18294_ (.Y(_11494_),
    .A(_00164_));
 sg13g2_nand2_1 _18295_ (.Y(_11495_),
    .A(_11494_),
    .B(_09218_));
 sg13g2_nand4_1 _18296_ (.B(net211),
    .C(_11493_),
    .A(net88),
    .Y(_11496_),
    .D(_11495_));
 sg13g2_nor2_1 _18297_ (.A(_00164_),
    .B(net732),
    .Y(_11497_));
 sg13g2_nand2_1 _18298_ (.Y(_11498_),
    .A(_11493_),
    .B(_11497_));
 sg13g2_buf_1 _18299_ (.A(_11125_),
    .X(_11499_));
 sg13g2_nand2b_1 _18300_ (.Y(_11500_),
    .B(net183),
    .A_N(_11498_));
 sg13g2_a22oi_1 _18301_ (.Y(_11501_),
    .B1(_11496_),
    .B2(_11500_),
    .A2(_11491_),
    .A1(_11490_));
 sg13g2_a21oi_1 _18302_ (.A1(_11485_),
    .A2(_11487_),
    .Y(_11502_),
    .B1(_11489_));
 sg13g2_and2_1 _18303_ (.A(_11042_),
    .B(_11481_),
    .X(_11503_));
 sg13g2_buf_1 _18304_ (.A(_11503_),
    .X(_11504_));
 sg13g2_nand3_1 _18305_ (.B(_11493_),
    .C(_11495_),
    .A(_11499_),
    .Y(_11505_));
 sg13g2_nor4_1 _18306_ (.A(net87),
    .B(_11502_),
    .C(_11504_),
    .D(_11505_),
    .Y(_11506_));
 sg13g2_nor4_1 _18307_ (.A(net183),
    .B(_11502_),
    .C(_11504_),
    .D(_11498_),
    .Y(_11507_));
 sg13g2_and2_1 _18308_ (.A(net542),
    .B(net89),
    .X(_11508_));
 sg13g2_buf_2 _18309_ (.A(_11508_),
    .X(_11509_));
 sg13g2_a22oi_1 _18310_ (.Y(_11510_),
    .B1(_11509_),
    .B2(_11494_),
    .A2(_10070_),
    .A1(\cpu.ex.r_mult[8] ));
 sg13g2_o21ai_1 _18311_ (.B1(_11510_),
    .Y(_11511_),
    .A1(net88),
    .A2(_11498_));
 sg13g2_or4_1 _18312_ (.A(_11501_),
    .B(_11506_),
    .C(_11507_),
    .D(_11511_),
    .X(\cpu.ex.c_mult[8] ));
 sg13g2_nor2_1 _18313_ (.A(net122),
    .B(net186),
    .Y(_11512_));
 sg13g2_inv_1 _18314_ (.Y(_11513_),
    .A(net212));
 sg13g2_nor2_1 _18315_ (.A(net122),
    .B(_11513_),
    .Y(_11514_));
 sg13g2_a21o_1 _18316_ (.A2(_11093_),
    .A1(_11075_),
    .B1(_11497_),
    .X(_11515_));
 sg13g2_buf_1 _18317_ (.A(_11515_),
    .X(_11516_));
 sg13g2_nand2_1 _18318_ (.Y(_11517_),
    .A(_11481_),
    .B(_11516_));
 sg13g2_nor4_2 _18319_ (.A(_11472_),
    .B(_11474_),
    .C(_11477_),
    .Y(_11518_),
    .D(_11517_));
 sg13g2_nand3_1 _18320_ (.B(_11042_),
    .C(_11516_),
    .A(net677),
    .Y(_11519_));
 sg13g2_nor4_2 _18321_ (.A(_11472_),
    .B(_11474_),
    .C(_11477_),
    .Y(_11520_),
    .D(_11519_));
 sg13g2_nor2_1 _18322_ (.A(_11094_),
    .B(_11495_),
    .Y(_11521_));
 sg13g2_a21o_1 _18323_ (.A2(_11516_),
    .A1(_11504_),
    .B1(_11521_),
    .X(_11522_));
 sg13g2_buf_1 _18324_ (.A(_11522_),
    .X(_11523_));
 sg13g2_nor3_1 _18325_ (.A(_11518_),
    .B(_11520_),
    .C(_11523_),
    .Y(_11524_));
 sg13g2_mux2_1 _18326_ (.A0(_11512_),
    .A1(_11514_),
    .S(_11524_),
    .X(_11525_));
 sg13g2_nor2_1 _18327_ (.A(_00165_),
    .B(net732),
    .Y(_11526_));
 sg13g2_buf_1 _18328_ (.A(_11526_),
    .X(_11527_));
 sg13g2_mux2_1 _18329_ (.A0(_11527_),
    .A1(_00165_),
    .S(_11525_),
    .X(_11528_));
 sg13g2_nor2b_1 _18330_ (.A(_00165_),
    .B_N(_11323_),
    .Y(_11529_));
 sg13g2_a221oi_1 _18331_ (.B2(_09215_),
    .C1(_11529_),
    .B1(_11528_),
    .A1(net604),
    .Y(_11530_),
    .A2(_11525_));
 sg13g2_nand2_1 _18332_ (.Y(_11531_),
    .A(\cpu.ex.r_mult[9] ),
    .B(net428));
 sg13g2_o21ai_1 _18333_ (.B1(_11531_),
    .Y(\cpu.ex.c_mult[9] ),
    .A1(_11335_),
    .A2(_11530_));
 sg13g2_nand2_1 _18334_ (.Y(_11532_),
    .A(net542),
    .B(net89));
 sg13g2_buf_1 _18335_ (.A(_11532_),
    .X(_11533_));
 sg13g2_nor2_1 _18336_ (.A(_11073_),
    .B(_11527_),
    .Y(_11534_));
 sg13g2_and2_1 _18337_ (.A(net212),
    .B(_11527_),
    .X(_11535_));
 sg13g2_buf_1 _18338_ (.A(_11535_),
    .X(_11536_));
 sg13g2_nor4_2 _18339_ (.A(_11518_),
    .B(_11520_),
    .C(_11523_),
    .Y(_11537_),
    .D(_11536_));
 sg13g2_nor2_1 _18340_ (.A(_11534_),
    .B(_11537_),
    .Y(_11538_));
 sg13g2_xnor2_1 _18341_ (.Y(_11539_),
    .A(net320),
    .B(_11538_));
 sg13g2_nand2_1 _18342_ (.Y(_11540_),
    .A(_09221_),
    .B(_10066_));
 sg13g2_buf_1 _18343_ (.A(_11540_),
    .X(_11541_));
 sg13g2_nor2_1 _18344_ (.A(net604),
    .B(_11541_),
    .Y(_11542_));
 sg13g2_buf_1 _18345_ (.A(_11542_),
    .X(_11543_));
 sg13g2_o21ai_1 _18346_ (.B1(_11543_),
    .Y(_11544_),
    .A1(net87),
    .A2(_11539_));
 sg13g2_a21oi_1 _18347_ (.A1(_11533_),
    .A2(_11544_),
    .Y(_11545_),
    .B1(_00166_));
 sg13g2_nor2_1 _18348_ (.A(_11394_),
    .B(_11539_),
    .Y(_11546_));
 sg13g2_nor2_1 _18349_ (.A(_00166_),
    .B(_09201_),
    .Y(_11547_));
 sg13g2_buf_2 _18350_ (.A(_11547_),
    .X(_11548_));
 sg13g2_nor2_1 _18351_ (.A(_11541_),
    .B(_11548_),
    .Y(_11549_));
 sg13g2_a22oi_1 _18352_ (.Y(_11550_),
    .B1(_11546_),
    .B2(_11549_),
    .A2(net428),
    .A1(\cpu.ex.r_mult[10] ));
 sg13g2_nor2b_1 _18353_ (.A(_11545_),
    .B_N(_11550_),
    .Y(_11551_));
 sg13g2_inv_1 _18354_ (.Y(\cpu.ex.c_mult[10] ),
    .A(_11551_));
 sg13g2_a21oi_1 _18355_ (.A1(net212),
    .A2(_11527_),
    .Y(_11552_),
    .B1(_11548_));
 sg13g2_nor2_1 _18356_ (.A(net319),
    .B(_11552_),
    .Y(_11553_));
 sg13g2_a21oi_1 _18357_ (.A1(_11536_),
    .A2(_11548_),
    .Y(_11554_),
    .B1(_11553_));
 sg13g2_o21ai_1 _18358_ (.B1(_11286_),
    .Y(_11555_),
    .A1(_11119_),
    .A2(_11548_));
 sg13g2_inv_1 _18359_ (.Y(_11556_),
    .A(_11555_));
 sg13g2_a221oi_1 _18360_ (.B2(_11327_),
    .C1(_11553_),
    .B1(_11556_),
    .A1(_11536_),
    .Y(_11557_),
    .A2(_11548_));
 sg13g2_nor4_1 _18361_ (.A(_10524_),
    .B(_10650_),
    .C(_10720_),
    .D(net319),
    .Y(_11558_));
 sg13g2_o21ai_1 _18362_ (.B1(_11527_),
    .Y(_11559_),
    .A1(_11548_),
    .A2(_11558_));
 sg13g2_a221oi_1 _18363_ (.B2(_11559_),
    .C1(net122),
    .B1(_11557_),
    .A1(_11524_),
    .Y(_11560_),
    .A2(_11554_));
 sg13g2_buf_1 _18364_ (.A(_11560_),
    .X(_11561_));
 sg13g2_buf_2 _18365_ (.A(_00167_),
    .X(_11562_));
 sg13g2_nor2_2 _18366_ (.A(_11562_),
    .B(net732),
    .Y(_11563_));
 sg13g2_buf_1 _18367_ (.A(_10169_),
    .X(_11564_));
 sg13g2_nand2_1 _18368_ (.Y(_11565_),
    .A(_11329_),
    .B(net208));
 sg13g2_xnor2_1 _18369_ (.Y(_11566_),
    .A(_11563_),
    .B(_11565_));
 sg13g2_xnor2_1 _18370_ (.Y(_11567_),
    .A(_11561_),
    .B(_11566_));
 sg13g2_inv_1 _18371_ (.Y(_11568_),
    .A(_11562_));
 sg13g2_a22oi_1 _18372_ (.Y(_11569_),
    .B1(_11509_),
    .B2(_11568_),
    .A2(net374),
    .A1(\cpu.ex.r_mult[11] ));
 sg13g2_o21ai_1 _18373_ (.B1(_11569_),
    .Y(\cpu.ex.c_mult[11] ),
    .A1(_11541_),
    .A2(_11567_));
 sg13g2_nand2_1 _18374_ (.Y(_11570_),
    .A(\cpu.ex.r_mult[12] ),
    .B(net428));
 sg13g2_inv_1 _18375_ (.Y(_11571_),
    .A(_11570_));
 sg13g2_buf_1 _18376_ (.A(_11173_),
    .X(_11572_));
 sg13g2_or3_1 _18377_ (.A(_11518_),
    .B(_11520_),
    .C(_11523_),
    .X(_11573_));
 sg13g2_mux2_1 _18378_ (.A0(_11562_),
    .A1(_11563_),
    .S(_11138_),
    .X(_11574_));
 sg13g2_a22oi_1 _18379_ (.Y(_11575_),
    .B1(_11574_),
    .B2(_00166_),
    .A2(_10169_),
    .A1(net732));
 sg13g2_xnor2_1 _18380_ (.Y(_11576_),
    .A(_11568_),
    .B(_11138_));
 sg13g2_nand2_1 _18381_ (.Y(_11577_),
    .A(_11548_),
    .B(_11576_));
 sg13g2_mux2_1 _18382_ (.A0(_11575_),
    .A1(_11577_),
    .S(_11291_),
    .X(_11578_));
 sg13g2_buf_1 _18383_ (.A(_11578_),
    .X(_11579_));
 sg13g2_nor2_1 _18384_ (.A(_11534_),
    .B(_11579_),
    .Y(_11580_));
 sg13g2_nand2_1 _18385_ (.Y(_11581_),
    .A(_11286_),
    .B(_11527_));
 sg13g2_nand3_1 _18386_ (.B(_11117_),
    .C(_11548_),
    .A(_11098_),
    .Y(_11582_));
 sg13g2_nand3_1 _18387_ (.B(_10167_),
    .C(_11563_),
    .A(_10077_),
    .Y(_11583_));
 sg13g2_a21oi_1 _18388_ (.A1(_10077_),
    .A2(_10167_),
    .Y(_11584_),
    .B1(_11563_));
 sg13g2_a21o_1 _18389_ (.A2(_11583_),
    .A1(_11582_),
    .B1(_11584_),
    .X(_11585_));
 sg13g2_buf_1 _18390_ (.A(_11585_),
    .X(_11586_));
 sg13g2_o21ai_1 _18391_ (.B1(_11586_),
    .Y(_11587_),
    .A1(_11581_),
    .A2(_11579_));
 sg13g2_a21oi_1 _18392_ (.A1(_11573_),
    .A2(_11580_),
    .Y(_11588_),
    .B1(_11587_));
 sg13g2_xnor2_1 _18393_ (.Y(_11589_),
    .A(_11572_),
    .B(_11588_));
 sg13g2_buf_1 _18394_ (.A(_00168_),
    .X(_11590_));
 sg13g2_nor2_1 _18395_ (.A(_11590_),
    .B(net732),
    .Y(_11591_));
 sg13g2_nor4_1 _18396_ (.A(net87),
    .B(_11541_),
    .C(_11589_),
    .D(_11591_),
    .Y(_11592_));
 sg13g2_o21ai_1 _18397_ (.B1(_11543_),
    .Y(_11593_),
    .A1(net87),
    .A2(_11589_));
 sg13g2_a21oi_1 _18398_ (.A1(_11533_),
    .A2(_11593_),
    .Y(_11594_),
    .B1(_11590_));
 sg13g2_or3_1 _18399_ (.A(_11571_),
    .B(_11592_),
    .C(_11594_),
    .X(\cpu.ex.c_mult[12] ));
 sg13g2_or2_1 _18400_ (.X(_11595_),
    .B(_11371_),
    .A(_11590_));
 sg13g2_nor3_1 _18401_ (.A(net99),
    .B(net246),
    .C(_11595_),
    .Y(_11596_));
 sg13g2_nor4_1 _18402_ (.A(_11562_),
    .B(net646),
    .C(net182),
    .D(net99),
    .Y(_11597_));
 sg13g2_o21ai_1 _18403_ (.B1(_11561_),
    .Y(_11598_),
    .A1(_11596_),
    .A2(_11597_));
 sg13g2_nor3_1 _18404_ (.A(_11562_),
    .B(_11590_),
    .C(net646),
    .Y(_11599_));
 sg13g2_nor3_1 _18405_ (.A(net182),
    .B(_11369_),
    .C(net246),
    .Y(_11600_));
 sg13g2_o21ai_1 _18406_ (.B1(_11561_),
    .Y(_11601_),
    .A1(_11599_),
    .A2(_11600_));
 sg13g2_nor4_1 _18407_ (.A(_11562_),
    .B(_11372_),
    .C(net182),
    .D(net246),
    .Y(_11602_));
 sg13g2_nand2_1 _18408_ (.Y(_11603_),
    .A(_10169_),
    .B(_11599_));
 sg13g2_nand2_1 _18409_ (.Y(_11604_),
    .A(_11177_),
    .B(_11591_));
 sg13g2_a21oi_1 _18410_ (.A1(_11603_),
    .A2(_11604_),
    .Y(_11605_),
    .B1(net99));
 sg13g2_a21oi_1 _18411_ (.A1(_11328_),
    .A2(_11602_),
    .Y(_11606_),
    .B1(_11605_));
 sg13g2_nand3_1 _18412_ (.B(_11601_),
    .C(_11606_),
    .A(_11598_),
    .Y(_11607_));
 sg13g2_buf_1 _18413_ (.A(_00169_),
    .X(_11608_));
 sg13g2_nor2_2 _18414_ (.A(_11608_),
    .B(_11371_),
    .Y(_11609_));
 sg13g2_nand2_1 _18415_ (.Y(_11610_),
    .A(net187),
    .B(net100));
 sg13g2_xnor2_1 _18416_ (.Y(_11611_),
    .A(_11609_),
    .B(_11610_));
 sg13g2_xnor2_1 _18417_ (.Y(_11612_),
    .A(_11607_),
    .B(_11611_));
 sg13g2_inv_1 _18418_ (.Y(_11613_),
    .A(_11608_));
 sg13g2_a22oi_1 _18419_ (.Y(_11614_),
    .B1(_11509_),
    .B2(_11613_),
    .A2(net428),
    .A1(\cpu.ex.r_mult[13] ));
 sg13g2_o21ai_1 _18420_ (.B1(_11614_),
    .Y(_11615_),
    .A1(_11541_),
    .A2(_11612_));
 sg13g2_buf_1 _18421_ (.A(_11615_),
    .X(\cpu.ex.c_mult[13] ));
 sg13g2_nand2_1 _18422_ (.Y(_11616_),
    .A(_11263_),
    .B(_11609_));
 sg13g2_nand2b_1 _18423_ (.Y(_11617_),
    .B(net210),
    .A_N(_11609_));
 sg13g2_buf_1 _18424_ (.A(_11617_),
    .X(_11618_));
 sg13g2_xnor2_1 _18425_ (.Y(_11619_),
    .A(_11173_),
    .B(_11591_));
 sg13g2_nand4_1 _18426_ (.B(_11616_),
    .C(_11618_),
    .A(_11327_),
    .Y(_11620_),
    .D(_11619_));
 sg13g2_nor4_2 _18427_ (.A(_11534_),
    .B(_11537_),
    .C(_11579_),
    .Y(_11621_),
    .D(_11620_));
 sg13g2_nand2_1 _18428_ (.Y(_11622_),
    .A(_11270_),
    .B(_11327_));
 sg13g2_buf_1 _18429_ (.A(_11270_),
    .X(_11623_));
 sg13g2_o21ai_1 _18430_ (.B1(_11595_),
    .Y(_11624_),
    .A1(_11173_),
    .A2(_11586_));
 sg13g2_nand2_1 _18431_ (.Y(_11625_),
    .A(_11173_),
    .B(_11586_));
 sg13g2_nand3_1 _18432_ (.B(_11624_),
    .C(_11625_),
    .A(_11618_),
    .Y(_11626_));
 sg13g2_nand3_1 _18433_ (.B(_11616_),
    .C(_11626_),
    .A(net163),
    .Y(_11627_));
 sg13g2_buf_1 _18434_ (.A(_11239_),
    .X(_11628_));
 sg13g2_and2_1 _18435_ (.A(_11263_),
    .B(_11609_),
    .X(_11629_));
 sg13g2_a21o_1 _18436_ (.A2(_11625_),
    .A1(_11624_),
    .B1(_11629_),
    .X(_11630_));
 sg13g2_nand3_1 _18437_ (.B(_11618_),
    .C(_11630_),
    .A(net162),
    .Y(_11631_));
 sg13g2_o21ai_1 _18438_ (.B1(_11631_),
    .Y(_11632_),
    .A1(_11621_),
    .A2(_11627_));
 sg13g2_a22oi_1 _18439_ (.Y(_11633_),
    .B1(_11632_),
    .B2(net88),
    .A2(_11622_),
    .A1(_11621_));
 sg13g2_buf_2 _18440_ (.A(_00170_),
    .X(_11634_));
 sg13g2_nor2_1 _18441_ (.A(_11634_),
    .B(net732),
    .Y(_11635_));
 sg13g2_xnor2_1 _18442_ (.Y(_11636_),
    .A(_11633_),
    .B(_11635_));
 sg13g2_nor2_1 _18443_ (.A(_11634_),
    .B(_11533_),
    .Y(_11637_));
 sg13g2_a221oi_1 _18444_ (.B2(_11636_),
    .C1(_11637_),
    .B1(_11493_),
    .A1(\cpu.ex.r_mult[14] ),
    .Y(_11638_),
    .A2(net374));
 sg13g2_inv_1 _18445_ (.Y(\cpu.ex.c_mult[14] ),
    .A(_11638_));
 sg13g2_or4_1 _18446_ (.A(_11205_),
    .B(_10524_),
    .C(_10650_),
    .D(_10720_),
    .X(_11639_));
 sg13g2_buf_1 _18447_ (.A(_11639_),
    .X(_11640_));
 sg13g2_buf_1 _18448_ (.A(_00171_),
    .X(_11641_));
 sg13g2_nor2_1 _18449_ (.A(_11641_),
    .B(net604),
    .Y(_11642_));
 sg13g2_xor2_1 _18450_ (.B(_11642_),
    .A(_11640_),
    .X(_11643_));
 sg13g2_nand2_1 _18451_ (.Y(_11644_),
    .A(_11493_),
    .B(_11643_));
 sg13g2_or2_1 _18452_ (.X(_11645_),
    .B(_11643_),
    .A(_11541_));
 sg13g2_o21ai_1 _18453_ (.B1(_11635_),
    .Y(_11646_),
    .A1(net163),
    .A2(_11629_));
 sg13g2_o21ai_1 _18454_ (.B1(_11646_),
    .Y(_11647_),
    .A1(net162),
    .A2(_11616_));
 sg13g2_nor2_1 _18455_ (.A(_11272_),
    .B(net99),
    .Y(_11648_));
 sg13g2_nor4_1 _18456_ (.A(_11608_),
    .B(_11634_),
    .C(net604),
    .D(_11648_),
    .Y(_11649_));
 sg13g2_mux2_1 _18457_ (.A0(_11634_),
    .A1(_11635_),
    .S(_11239_),
    .X(_11650_));
 sg13g2_a22oi_1 _18458_ (.Y(_11651_),
    .B1(_11650_),
    .B2(_11608_),
    .A2(net163),
    .A1(net646));
 sg13g2_or2_1 _18459_ (.X(_11652_),
    .B(_11651_),
    .A(net210));
 sg13g2_nand3_1 _18460_ (.B(_11264_),
    .C(_11609_),
    .A(_11634_),
    .Y(_11653_));
 sg13g2_a21oi_1 _18461_ (.A1(_11652_),
    .A2(_11653_),
    .Y(_11654_),
    .B1(_11394_));
 sg13g2_nor2_1 _18462_ (.A(_11649_),
    .B(_11654_),
    .Y(_11655_));
 sg13g2_inv_1 _18463_ (.Y(_11656_),
    .A(_11655_));
 sg13g2_a22oi_1 _18464_ (.Y(_11657_),
    .B1(_11656_),
    .B2(_11607_),
    .A2(_11647_),
    .A1(_11329_));
 sg13g2_mux2_1 _18465_ (.A0(_11644_),
    .A1(_11645_),
    .S(_11657_),
    .X(_11658_));
 sg13g2_buf_1 _18466_ (.A(_11509_),
    .X(_11659_));
 sg13g2_inv_1 _18467_ (.Y(_11660_),
    .A(_11641_));
 sg13g2_a22oi_1 _18468_ (.Y(_11661_),
    .B1(net61),
    .B2(_11660_),
    .A2(_10071_),
    .A1(\cpu.ex.r_mult[15] ));
 sg13g2_nand2_1 _18469_ (.Y(\cpu.ex.c_mult[15] ),
    .A(_11658_),
    .B(_11661_));
 sg13g2_inv_1 _18470_ (.Y(_00000_),
    .A(net2));
 sg13g2_nand2_1 _18471_ (.Y(_11662_),
    .A(_09703_),
    .B(_09705_));
 sg13g2_nor2_1 _18472_ (.A(net617),
    .B(_11662_),
    .Y(_00007_));
 sg13g2_buf_1 _18473_ (.A(net781),
    .X(_11663_));
 sg13g2_and3_1 _18474_ (.X(_00008_),
    .A(_09677_),
    .B(net645),
    .C(net107));
 sg13g2_buf_1 _18475_ (.A(\cpu.qspi.r_state[11] ),
    .X(_11664_));
 sg13g2_and2_1 _18476_ (.A(_11664_),
    .B(net645),
    .X(_00004_));
 sg13g2_buf_2 _18477_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11665_));
 sg13g2_and2_1 _18478_ (.A(_11665_),
    .B(net645),
    .X(_00009_));
 sg13g2_buf_2 _18479_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11666_));
 sg13g2_and2_1 _18480_ (.A(_11666_),
    .B(net645),
    .X(_00003_));
 sg13g2_buf_1 _18481_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11667_));
 sg13g2_and2_1 _18482_ (.A(_11667_),
    .B(_11663_),
    .X(_00002_));
 sg13g2_and3_1 _18483_ (.X(_00001_),
    .A(_09673_),
    .B(net645),
    .C(_09670_));
 sg13g2_nor2_1 _18484_ (.A(_10222_),
    .B(_10285_),
    .Y(_11668_));
 sg13g2_nand2_1 _18485_ (.Y(_11669_),
    .A(_10354_),
    .B(_10392_));
 sg13g2_and4_1 _18486_ (.A(_11669_),
    .B(_10430_),
    .C(_10573_),
    .D(_10645_),
    .X(_11670_));
 sg13g2_nand4_1 _18487_ (.B(_10547_),
    .C(_10693_),
    .A(_10600_),
    .Y(_11671_),
    .D(_11670_));
 sg13g2_or2_1 _18488_ (.X(_11672_),
    .B(_10347_),
    .A(_10327_));
 sg13g2_a221oi_1 _18489_ (.B2(_10714_),
    .C1(_10456_),
    .B1(_10696_),
    .A1(_10461_),
    .Y(_11673_),
    .A2(_10484_));
 sg13g2_nand4_1 _18490_ (.B(_10516_),
    .C(_10675_),
    .A(_11672_),
    .Y(_11674_),
    .D(_11673_));
 sg13g2_nor4_1 _18491_ (.A(_10325_),
    .B(_11668_),
    .C(_11671_),
    .D(_11674_),
    .Y(_11675_));
 sg13g2_o21ai_1 _18492_ (.B1(_10619_),
    .Y(_11676_),
    .A1(\cpu.cond[1] ),
    .A2(_11675_));
 sg13g2_xnor2_1 _18493_ (.Y(_11677_),
    .A(net1033),
    .B(_11676_));
 sg13g2_a21o_1 _18494_ (.A2(_11677_),
    .A1(_00273_),
    .B1(_10203_),
    .X(_11678_));
 sg13g2_nor2b_1 _18495_ (.A(\cpu.dec.jmp ),
    .B_N(_11678_),
    .Y(_11679_));
 sg13g2_nor2_1 _18496_ (.A(_11343_),
    .B(_11679_),
    .Y(_00053_));
 sg13g2_and3_1 _18497_ (.X(_00005_),
    .A(net1102),
    .B(net781),
    .C(_09670_));
 sg13g2_buf_2 _18498_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11680_));
 sg13g2_and2_1 _18499_ (.A(_11680_),
    .B(net645),
    .X(_00006_));
 sg13g2_buf_2 _18500_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11681_));
 sg13g2_and2_1 _18501_ (.A(_11681_),
    .B(net645),
    .X(_00010_));
 sg13g2_nor2_1 _18502_ (.A(net91),
    .B(net617),
    .Y(_00052_));
 sg13g2_or2_1 _18503_ (.X(_11682_),
    .B(net1105),
    .A(_09136_));
 sg13g2_buf_1 _18504_ (.A(_11682_),
    .X(_11683_));
 sg13g2_nor3_1 _18505_ (.A(_09116_),
    .B(net1104),
    .C(_11683_),
    .Y(_11684_));
 sg13g2_a21oi_1 _18506_ (.A1(_09009_),
    .A2(_11683_),
    .Y(_11685_),
    .B1(_11684_));
 sg13g2_nand2_1 _18507_ (.Y(_11686_),
    .A(_09124_),
    .B(_11685_));
 sg13g2_inv_1 _18508_ (.Y(_11687_),
    .A(_00226_));
 sg13g2_nor3_2 _18509_ (.A(net1105),
    .B(net1104),
    .C(_11687_),
    .Y(_11688_));
 sg13g2_buf_1 _18510_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11689_));
 sg13g2_buf_1 _18511_ (.A(_11689_),
    .X(_11690_));
 sg13g2_buf_1 _18512_ (.A(\cpu.spi.r_src[2] ),
    .X(_11691_));
 sg13g2_inv_1 _18513_ (.Y(_11692_),
    .A(_00282_));
 sg13g2_buf_2 _18514_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11693_));
 sg13g2_buf_1 _18515_ (.A(_11693_),
    .X(_11694_));
 sg13g2_mux2_1 _18516_ (.A0(_11691_),
    .A1(_11692_),
    .S(_11694_),
    .X(_11695_));
 sg13g2_buf_1 _18517_ (.A(_11689_),
    .X(_11696_));
 sg13g2_buf_1 _18518_ (.A(_11693_),
    .X(_11697_));
 sg13g2_nand2_1 _18519_ (.Y(_11698_),
    .A(_11697_),
    .B(_00283_));
 sg13g2_o21ai_1 _18520_ (.B1(_11698_),
    .Y(_11699_),
    .A1(net998),
    .A2(_11692_));
 sg13g2_nor2_1 _18521_ (.A(_11696_),
    .B(_11699_),
    .Y(_11700_));
 sg13g2_a21oi_2 _18522_ (.B1(_11700_),
    .Y(_11701_),
    .A2(_11695_),
    .A1(net999));
 sg13g2_nor2_1 _18523_ (.A(_11688_),
    .B(_11701_),
    .Y(_11702_));
 sg13g2_nor2_1 _18524_ (.A(net1029),
    .B(net1104),
    .Y(_11703_));
 sg13g2_inv_1 _18525_ (.Y(_11704_),
    .A(_11689_));
 sg13g2_buf_1 _18526_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11705_));
 sg13g2_buf_1 _18527_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11706_));
 sg13g2_buf_1 _18528_ (.A(net996),
    .X(_11707_));
 sg13g2_mux2_1 _18529_ (.A0(_11705_),
    .A1(_11706_),
    .S(net867),
    .X(_11708_));
 sg13g2_nor2_1 _18530_ (.A(_11704_),
    .B(_11693_),
    .Y(_11709_));
 sg13g2_buf_1 _18531_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11710_));
 sg13g2_a22oi_1 _18532_ (.Y(_11711_),
    .B1(_11709_),
    .B2(_11710_),
    .A2(_11708_),
    .A1(_11704_));
 sg13g2_xnor2_1 _18533_ (.Y(_11712_),
    .A(_11703_),
    .B(_11711_));
 sg13g2_or3_1 _18534_ (.A(net1105),
    .B(net1104),
    .C(_11687_),
    .X(_11713_));
 sg13g2_buf_1 _18535_ (.A(_11713_),
    .X(_11714_));
 sg13g2_buf_1 _18536_ (.A(_10431_),
    .X(_11715_));
 sg13g2_inv_1 _18537_ (.Y(_11716_),
    .A(_00283_));
 sg13g2_buf_1 _18538_ (.A(net670),
    .X(_11717_));
 sg13g2_buf_1 _18539_ (.A(net603),
    .X(_11718_));
 sg13g2_buf_2 _18540_ (.A(net537),
    .X(_11719_));
 sg13g2_mux2_1 _18541_ (.A0(_11692_),
    .A1(_11716_),
    .S(net489),
    .X(_11720_));
 sg13g2_nor2_2 _18542_ (.A(_10431_),
    .B(_11719_),
    .Y(_11721_));
 sg13g2_a22oi_1 _18543_ (.Y(_11722_),
    .B1(_11721_),
    .B2(_11691_),
    .A2(_11720_),
    .A1(net865));
 sg13g2_nor2_1 _18544_ (.A(net866),
    .B(_11722_),
    .Y(_11723_));
 sg13g2_buf_1 _18545_ (.A(_09818_),
    .X(_11724_));
 sg13g2_buf_1 _18546_ (.A(net995),
    .X(_11725_));
 sg13g2_buf_1 _18547_ (.A(_11725_),
    .X(_11726_));
 sg13g2_buf_1 _18548_ (.A(net731),
    .X(_11727_));
 sg13g2_buf_1 _18549_ (.A(net489),
    .X(_11728_));
 sg13g2_nand2b_1 _18550_ (.Y(_11729_),
    .B(net489),
    .A_N(_11705_));
 sg13g2_o21ai_1 _18551_ (.B1(_11729_),
    .Y(_11730_),
    .A1(_11728_),
    .A2(_11710_));
 sg13g2_mux2_1 _18552_ (.A0(_11705_),
    .A1(_11706_),
    .S(net489),
    .X(_11731_));
 sg13g2_nor2_1 _18553_ (.A(net731),
    .B(_11731_),
    .Y(_11732_));
 sg13g2_a21oi_1 _18554_ (.A1(_11727_),
    .A2(_11730_),
    .Y(_11733_),
    .B1(_11732_));
 sg13g2_a22oi_1 _18555_ (.Y(_11734_),
    .B1(_11723_),
    .B2(_11733_),
    .A2(_11712_),
    .A1(_11702_));
 sg13g2_nor2_1 _18556_ (.A(_11702_),
    .B(_11723_),
    .Y(_11735_));
 sg13g2_buf_1 _18557_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_11736_));
 sg13g2_o21ai_1 _18558_ (.B1(_11736_),
    .Y(_11737_),
    .A1(_11686_),
    .A2(_11735_));
 sg13g2_o21ai_1 _18559_ (.B1(_11737_),
    .Y(_00318_),
    .A1(_11686_),
    .A2(_11734_));
 sg13g2_mux2_1 _18560_ (.A0(_11712_),
    .A1(_11733_),
    .S(_11688_),
    .X(_11738_));
 sg13g2_buf_1 _18561_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_11739_));
 sg13g2_nand3_1 _18562_ (.B(_11685_),
    .C(_11735_),
    .A(_09124_),
    .Y(_11740_));
 sg13g2_mux2_1 _18563_ (.A0(_11738_),
    .A1(_11739_),
    .S(_11740_),
    .X(_00319_));
 sg13g2_buf_1 _18564_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_11741_));
 sg13g2_mux2_1 _18565_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_09940_),
    .S(net1028),
    .X(_11742_));
 sg13g2_inv_1 _18566_ (.Y(_11743_),
    .A(_00224_));
 sg13g2_mux2_1 _18567_ (.A0(_11743_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_11693_),
    .X(_11744_));
 sg13g2_a22oi_1 _18568_ (.Y(_11745_),
    .B1(_11744_),
    .B2(_11704_),
    .A2(_11709_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18569_ (.A(_11745_),
    .X(_11746_));
 sg13g2_nand2_1 _18570_ (.Y(_11747_),
    .A(_09139_),
    .B(_11746_));
 sg13g2_a21oi_1 _18571_ (.A1(_00221_),
    .A2(_09144_),
    .Y(_11748_),
    .B1(_09176_));
 sg13g2_nor2b_1 _18572_ (.A(_11747_),
    .B_N(_11748_),
    .Y(_11749_));
 sg13g2_o21ai_1 _18573_ (.B1(net1105),
    .Y(_11750_),
    .A1(_09009_),
    .A2(_11746_));
 sg13g2_nor2b_1 _18574_ (.A(net1029),
    .B_N(_11750_),
    .Y(_11751_));
 sg13g2_o21ai_1 _18575_ (.B1(net897),
    .Y(_11752_),
    .A1(_11749_),
    .A2(_11751_));
 sg13g2_buf_1 _18576_ (.A(_11746_),
    .X(_11753_));
 sg13g2_a21oi_1 _18577_ (.A1(net70),
    .A2(net602),
    .Y(_11754_),
    .B1(_09106_));
 sg13g2_nor3_1 _18578_ (.A(_09105_),
    .B(net1104),
    .C(_11683_),
    .Y(_11755_));
 sg13g2_nor3_1 _18579_ (.A(_11752_),
    .B(_11754_),
    .C(_11755_),
    .Y(_11756_));
 sg13g2_nor2b_1 _18580_ (.A(_11701_),
    .B_N(_11756_),
    .Y(_11757_));
 sg13g2_mux2_1 _18581_ (.A0(net1083),
    .A1(_11742_),
    .S(_11757_),
    .X(_00320_));
 sg13g2_buf_1 _18582_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_11758_));
 sg13g2_nand2_1 _18583_ (.Y(_11759_),
    .A(_11701_),
    .B(_11756_));
 sg13g2_mux2_1 _18584_ (.A0(_11742_),
    .A1(net1082),
    .S(_11759_),
    .X(_00321_));
 sg13g2_buf_1 _18585_ (.A(uio_in[0]),
    .X(_11760_));
 sg13g2_buf_2 _18586_ (.A(_11760_),
    .X(_11761_));
 sg13g2_buf_1 _18587_ (.A(net673),
    .X(_11762_));
 sg13g2_nand2_1 _18588_ (.Y(_11763_),
    .A(net1025),
    .B(net601));
 sg13g2_buf_1 _18589_ (.A(_11763_),
    .X(_11764_));
 sg13g2_buf_1 _18590_ (.A(\cpu.d_wstrobe_d ),
    .X(_11765_));
 sg13g2_buf_1 _18591_ (.A(_11765_),
    .X(_11766_));
 sg13g2_buf_1 _18592_ (.A(_00276_),
    .X(_11767_));
 sg13g2_buf_1 _18593_ (.A(_11767_),
    .X(_11768_));
 sg13g2_buf_1 _18594_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_11769_));
 sg13g2_buf_1 _18595_ (.A(_11769_),
    .X(_11770_));
 sg13g2_buf_2 _18596_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_11771_));
 sg13g2_nor2b_1 _18597_ (.A(_11770_),
    .B_N(_11771_),
    .Y(_11772_));
 sg13g2_nand3_1 _18598_ (.B(net993),
    .C(_11772_),
    .A(net994),
    .Y(_11773_));
 sg13g2_buf_2 _18599_ (.A(_11773_),
    .X(_11774_));
 sg13g2_or2_1 _18600_ (.X(_11775_),
    .B(_11774_),
    .A(net488));
 sg13g2_buf_1 _18601_ (.A(_11775_),
    .X(_11776_));
 sg13g2_mux2_1 _18602_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][0] ),
    .S(_11776_),
    .X(_11777_));
 sg13g2_buf_1 _18603_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_11778_));
 sg13g2_and2_1 _18604_ (.A(_11769_),
    .B(_11771_),
    .X(_11779_));
 sg13g2_buf_1 _18605_ (.A(_11779_),
    .X(_11780_));
 sg13g2_and3_1 _18606_ (.X(_11781_),
    .A(net1080),
    .B(_11765_),
    .C(net863));
 sg13g2_buf_1 _18607_ (.A(_11781_),
    .X(_11782_));
 sg13g2_nor3_1 _18608_ (.A(_09223_),
    .B(_08764_),
    .C(_09657_),
    .Y(_11783_));
 sg13g2_o21ai_1 _18609_ (.B1(_11783_),
    .Y(_11784_),
    .A1(_09653_),
    .A2(_11782_));
 sg13g2_buf_1 _18610_ (.A(_11784_),
    .X(_11785_));
 sg13g2_or2_1 _18611_ (.X(_11786_),
    .B(_11785_),
    .A(_11763_));
 sg13g2_buf_1 _18612_ (.A(_11786_),
    .X(_11787_));
 sg13g2_nand2_1 _18613_ (.Y(_11788_),
    .A(_08762_),
    .B(net886));
 sg13g2_buf_1 _18614_ (.A(_11788_),
    .X(_11789_));
 sg13g2_buf_2 _18615_ (.A(_00275_),
    .X(_11790_));
 sg13g2_o21ai_1 _18616_ (.B1(_11790_),
    .Y(_11791_),
    .A1(net1107),
    .A2(_11789_));
 sg13g2_nor2_1 _18617_ (.A(_11787_),
    .B(_11791_),
    .Y(_11792_));
 sg13g2_buf_4 _18618_ (.X(_11793_),
    .A(_11792_));
 sg13g2_mux2_1 _18619_ (.A0(_11777_),
    .A1(net884),
    .S(_11793_),
    .X(_00322_));
 sg13g2_buf_1 _18620_ (.A(uio_in[2]),
    .X(_11794_));
 sg13g2_buf_2 _18621_ (.A(_11794_),
    .X(_11795_));
 sg13g2_nand3_1 _18622_ (.B(net993),
    .C(net863),
    .A(net994),
    .Y(_11796_));
 sg13g2_buf_2 _18623_ (.A(_11796_),
    .X(_11797_));
 sg13g2_or2_1 _18624_ (.X(_11798_),
    .B(_11797_),
    .A(net488));
 sg13g2_buf_1 _18625_ (.A(_11798_),
    .X(_11799_));
 sg13g2_mux2_1 _18626_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][10] ),
    .S(_11799_),
    .X(_11800_));
 sg13g2_nor2b_1 _18627_ (.A(net1031),
    .B_N(_08762_),
    .Y(_11801_));
 sg13g2_and2_1 _18628_ (.A(net1107),
    .B(_11801_),
    .X(_11802_));
 sg13g2_buf_2 _18629_ (.A(_11802_),
    .X(_11803_));
 sg13g2_mux2_1 _18630_ (.A0(_09909_),
    .A1(_10018_),
    .S(_11803_),
    .X(_11804_));
 sg13g2_buf_2 _18631_ (.A(_11804_),
    .X(_11805_));
 sg13g2_buf_1 _18632_ (.A(_11805_),
    .X(_11806_));
 sg13g2_inv_1 _18633_ (.Y(_11807_),
    .A(_11790_));
 sg13g2_mux2_1 _18634_ (.A0(net991),
    .A1(_09118_),
    .S(net1107),
    .X(_11808_));
 sg13g2_nor3_1 _18635_ (.A(_11787_),
    .B(_11789_),
    .C(_11808_),
    .Y(_11809_));
 sg13g2_buf_1 _18636_ (.A(_11809_),
    .X(_11810_));
 sg13g2_mux2_1 _18637_ (.A0(_11800_),
    .A1(net487),
    .S(net65),
    .X(_00323_));
 sg13g2_buf_1 _18638_ (.A(uio_in[3]),
    .X(_11811_));
 sg13g2_buf_2 _18639_ (.A(_11811_),
    .X(_11812_));
 sg13g2_mux2_1 _18640_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][11] ),
    .S(_11799_),
    .X(_11813_));
 sg13g2_mux2_1 _18641_ (.A0(net1098),
    .A1(_10025_),
    .S(_11803_),
    .X(_11814_));
 sg13g2_buf_2 _18642_ (.A(_11814_),
    .X(_11815_));
 sg13g2_buf_1 _18643_ (.A(_11815_),
    .X(_11816_));
 sg13g2_mux2_1 _18644_ (.A0(_11813_),
    .A1(net486),
    .S(net65),
    .X(_00324_));
 sg13g2_nand2_1 _18645_ (.Y(_11817_),
    .A(net1107),
    .B(_11801_));
 sg13g2_and2_1 _18646_ (.A(_10030_),
    .B(_11803_),
    .X(_11818_));
 sg13g2_a21oi_1 _18647_ (.A1(_09921_),
    .A2(_11817_),
    .Y(_11819_),
    .B1(_11818_));
 sg13g2_buf_2 _18648_ (.A(_11819_),
    .X(_11820_));
 sg13g2_nor2b_1 _18649_ (.A(_11771_),
    .B_N(_11769_),
    .Y(_11821_));
 sg13g2_nand3_1 _18650_ (.B(_11767_),
    .C(_11821_),
    .A(net994),
    .Y(_11822_));
 sg13g2_buf_4 _18651_ (.X(_11823_),
    .A(_11822_));
 sg13g2_or2_1 _18652_ (.X(_11824_),
    .B(_11823_),
    .A(net488));
 sg13g2_buf_1 _18653_ (.A(_11824_),
    .X(_11825_));
 sg13g2_mux2_1 _18654_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][12] ),
    .S(_11825_),
    .X(_11826_));
 sg13g2_nor2_1 _18655_ (.A(net65),
    .B(_11826_),
    .Y(_11827_));
 sg13g2_a21oi_1 _18656_ (.A1(net65),
    .A2(_11820_),
    .Y(_00325_),
    .B1(_11827_));
 sg13g2_and2_1 _18657_ (.A(_10036_),
    .B(_11803_),
    .X(_11828_));
 sg13g2_a21oi_1 _18658_ (.A1(_09927_),
    .A2(_11817_),
    .Y(_11829_),
    .B1(_11828_));
 sg13g2_buf_2 _18659_ (.A(_11829_),
    .X(_11830_));
 sg13g2_buf_1 _18660_ (.A(uio_in[1]),
    .X(_11831_));
 sg13g2_buf_2 _18661_ (.A(_11831_),
    .X(_11832_));
 sg13g2_mux2_1 _18662_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][13] ),
    .S(_11825_),
    .X(_11833_));
 sg13g2_nor2_1 _18663_ (.A(net65),
    .B(_11833_),
    .Y(_11834_));
 sg13g2_a21oi_1 _18664_ (.A1(_11810_),
    .A2(_11830_),
    .Y(_00326_),
    .B1(_11834_));
 sg13g2_and2_1 _18665_ (.A(_10043_),
    .B(_11803_),
    .X(_11835_));
 sg13g2_a21oi_1 _18666_ (.A1(_09933_),
    .A2(_11817_),
    .Y(_11836_),
    .B1(_11835_));
 sg13g2_buf_2 _18667_ (.A(_11836_),
    .X(_11837_));
 sg13g2_mux2_1 _18668_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][14] ),
    .S(_11825_),
    .X(_11838_));
 sg13g2_nor2_1 _18669_ (.A(_11809_),
    .B(_11838_),
    .Y(_11839_));
 sg13g2_a21oi_1 _18670_ (.A1(_11810_),
    .A2(_11837_),
    .Y(_00327_),
    .B1(_11839_));
 sg13g2_and2_1 _18671_ (.A(_10048_),
    .B(_11803_),
    .X(_11840_));
 sg13g2_a21oi_1 _18672_ (.A1(_09940_),
    .A2(_11817_),
    .Y(_11841_),
    .B1(_11840_));
 sg13g2_buf_2 _18673_ (.A(_11841_),
    .X(_11842_));
 sg13g2_mux2_1 _18674_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][15] ),
    .S(_11825_),
    .X(_11843_));
 sg13g2_nor2_1 _18675_ (.A(_11809_),
    .B(_11843_),
    .Y(_11844_));
 sg13g2_a21oi_1 _18676_ (.A1(net65),
    .A2(_11842_),
    .Y(_00328_),
    .B1(_11844_));
 sg13g2_nand3_1 _18677_ (.B(net994),
    .C(_11772_),
    .A(net1080),
    .Y(_11845_));
 sg13g2_buf_2 _18678_ (.A(_11845_),
    .X(_11846_));
 sg13g2_or2_1 _18679_ (.X(_11847_),
    .B(_11846_),
    .A(net488));
 sg13g2_buf_1 _18680_ (.A(_11847_),
    .X(_11848_));
 sg13g2_mux2_1 _18681_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][16] ),
    .S(_11848_),
    .X(_11849_));
 sg13g2_buf_1 _18682_ (.A(_09117_),
    .X(_11850_));
 sg13g2_o21ai_1 _18683_ (.B1(net730),
    .Y(_11851_),
    .A1(net1107),
    .A2(_11789_));
 sg13g2_nor2_1 _18684_ (.A(_11787_),
    .B(_11851_),
    .Y(_11852_));
 sg13g2_buf_4 _18685_ (.X(_11853_),
    .A(_11852_));
 sg13g2_mux2_1 _18686_ (.A0(_11849_),
    .A1(net884),
    .S(_11853_),
    .X(_00329_));
 sg13g2_mux2_1 _18687_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][17] ),
    .S(_11848_),
    .X(_11854_));
 sg13g2_mux2_1 _18688_ (.A0(_11854_),
    .A1(net883),
    .S(_11853_),
    .X(_00330_));
 sg13g2_mux2_1 _18689_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][18] ),
    .S(_11848_),
    .X(_11855_));
 sg13g2_buf_1 _18690_ (.A(net1018),
    .X(_11856_));
 sg13g2_mux2_1 _18691_ (.A0(_11855_),
    .A1(net862),
    .S(_11853_),
    .X(_00331_));
 sg13g2_mux2_1 _18692_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][19] ),
    .S(_11848_),
    .X(_11857_));
 sg13g2_buf_1 _18693_ (.A(net1098),
    .X(_11858_));
 sg13g2_mux2_1 _18694_ (.A0(_11857_),
    .A1(net990),
    .S(_11853_),
    .X(_00332_));
 sg13g2_mux2_1 _18695_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][1] ),
    .S(_11776_),
    .X(_11859_));
 sg13g2_mux2_1 _18696_ (.A0(_11859_),
    .A1(net883),
    .S(_11793_),
    .X(_00333_));
 sg13g2_nor2_1 _18697_ (.A(_11769_),
    .B(_11771_),
    .Y(_11860_));
 sg13g2_nand3_1 _18698_ (.B(net994),
    .C(_11860_),
    .A(net1080),
    .Y(_11861_));
 sg13g2_buf_2 _18699_ (.A(_11861_),
    .X(_11862_));
 sg13g2_or2_1 _18700_ (.X(_11863_),
    .B(_11862_),
    .A(net488));
 sg13g2_buf_1 _18701_ (.A(_11863_),
    .X(_11864_));
 sg13g2_mux2_1 _18702_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][20] ),
    .S(_11864_),
    .X(_11865_));
 sg13g2_buf_1 _18703_ (.A(_09921_),
    .X(_11866_));
 sg13g2_mux2_1 _18704_ (.A0(_11865_),
    .A1(_11866_),
    .S(_11853_),
    .X(_00334_));
 sg13g2_mux2_1 _18705_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][21] ),
    .S(_11864_),
    .X(_11867_));
 sg13g2_buf_1 _18706_ (.A(_09927_),
    .X(_11868_));
 sg13g2_mux2_1 _18707_ (.A0(_11867_),
    .A1(_11868_),
    .S(_11853_),
    .X(_00335_));
 sg13g2_mux2_1 _18708_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][22] ),
    .S(_11864_),
    .X(_11869_));
 sg13g2_buf_1 _18709_ (.A(_09933_),
    .X(_11870_));
 sg13g2_mux2_1 _18710_ (.A0(_11869_),
    .A1(_11870_),
    .S(_11853_),
    .X(_00336_));
 sg13g2_mux2_1 _18711_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][23] ),
    .S(_11864_),
    .X(_11871_));
 sg13g2_mux2_1 _18712_ (.A0(_11871_),
    .A1(_09941_),
    .S(_11853_),
    .X(_00337_));
 sg13g2_nand2b_1 _18713_ (.Y(_11872_),
    .B(_11782_),
    .A_N(net488));
 sg13g2_buf_2 _18714_ (.A(_11872_),
    .X(_11873_));
 sg13g2_mux2_1 _18715_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(_11873_),
    .X(_11874_));
 sg13g2_mux2_1 _18716_ (.A0(_09895_),
    .A1(_10008_),
    .S(_11803_),
    .X(_11875_));
 sg13g2_buf_2 _18717_ (.A(_11875_),
    .X(_11876_));
 sg13g2_buf_1 _18718_ (.A(_11876_),
    .X(_11877_));
 sg13g2_nand2_1 _18719_ (.Y(_11878_),
    .A(net1107),
    .B(_11790_));
 sg13g2_o21ai_1 _18720_ (.B1(_11878_),
    .Y(_11879_),
    .A1(net1107),
    .A2(net782));
 sg13g2_nor3_1 _18721_ (.A(_11787_),
    .B(_11789_),
    .C(_11879_),
    .Y(_11880_));
 sg13g2_buf_1 _18722_ (.A(_11880_),
    .X(_11881_));
 sg13g2_mux2_1 _18723_ (.A0(_11874_),
    .A1(net485),
    .S(net64),
    .X(_00338_));
 sg13g2_mux2_1 _18724_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(_11873_),
    .X(_11882_));
 sg13g2_mux2_1 _18725_ (.A0(_09904_),
    .A1(_10013_),
    .S(_11803_),
    .X(_11883_));
 sg13g2_buf_2 _18726_ (.A(_11883_),
    .X(_11884_));
 sg13g2_buf_1 _18727_ (.A(_11884_),
    .X(_11885_));
 sg13g2_mux2_1 _18728_ (.A0(_11882_),
    .A1(net484),
    .S(_11881_),
    .X(_00339_));
 sg13g2_mux2_1 _18729_ (.A0(_11795_),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(_11873_),
    .X(_11886_));
 sg13g2_mux2_1 _18730_ (.A0(_11886_),
    .A1(net487),
    .S(net64),
    .X(_00340_));
 sg13g2_mux2_1 _18731_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(_11873_),
    .X(_11887_));
 sg13g2_mux2_1 _18732_ (.A0(_11887_),
    .A1(net486),
    .S(net64),
    .X(_00341_));
 sg13g2_buf_1 _18733_ (.A(_11820_),
    .X(_11888_));
 sg13g2_nand3_1 _18734_ (.B(_11765_),
    .C(_11821_),
    .A(_11778_),
    .Y(_11889_));
 sg13g2_buf_4 _18735_ (.X(_11890_),
    .A(_11889_));
 sg13g2_or2_1 _18736_ (.X(_11891_),
    .B(_11890_),
    .A(_11764_));
 sg13g2_buf_1 _18737_ (.A(_11891_),
    .X(_11892_));
 sg13g2_mux2_1 _18738_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][28] ),
    .S(_11892_),
    .X(_11893_));
 sg13g2_nor2_1 _18739_ (.A(net64),
    .B(_11893_),
    .Y(_11894_));
 sg13g2_a21oi_1 _18740_ (.A1(net423),
    .A2(net64),
    .Y(_00342_),
    .B1(_11894_));
 sg13g2_buf_1 _18741_ (.A(_11830_),
    .X(_11895_));
 sg13g2_mux2_1 _18742_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][29] ),
    .S(_11892_),
    .X(_11896_));
 sg13g2_nor2_1 _18743_ (.A(net64),
    .B(_11896_),
    .Y(_11897_));
 sg13g2_a21oi_1 _18744_ (.A1(net422),
    .A2(net64),
    .Y(_00343_),
    .B1(_11897_));
 sg13g2_mux2_1 _18745_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][2] ),
    .S(_11776_),
    .X(_11898_));
 sg13g2_mux2_1 _18746_ (.A0(_11898_),
    .A1(net862),
    .S(_11793_),
    .X(_00344_));
 sg13g2_buf_1 _18747_ (.A(_11837_),
    .X(_11899_));
 sg13g2_mux2_1 _18748_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][30] ),
    .S(_11892_),
    .X(_11900_));
 sg13g2_nor2_1 _18749_ (.A(_11880_),
    .B(_11900_),
    .Y(_11901_));
 sg13g2_a21oi_1 _18750_ (.A1(net421),
    .A2(net64),
    .Y(_00345_),
    .B1(_11901_));
 sg13g2_buf_1 _18751_ (.A(_11842_),
    .X(_11902_));
 sg13g2_mux2_1 _18752_ (.A0(_11812_),
    .A1(\cpu.dcache.r_data[0][31] ),
    .S(_11892_),
    .X(_11903_));
 sg13g2_nor2_1 _18753_ (.A(_11880_),
    .B(_11903_),
    .Y(_11904_));
 sg13g2_a21oi_1 _18754_ (.A1(_11902_),
    .A2(_11881_),
    .Y(_00346_),
    .B1(_11904_));
 sg13g2_mux2_1 _18755_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][3] ),
    .S(_11776_),
    .X(_11905_));
 sg13g2_mux2_1 _18756_ (.A0(_11905_),
    .A1(net990),
    .S(_11793_),
    .X(_00347_));
 sg13g2_nand3_1 _18757_ (.B(net993),
    .C(_11860_),
    .A(net994),
    .Y(_11906_));
 sg13g2_buf_2 _18758_ (.A(_11906_),
    .X(_11907_));
 sg13g2_or2_1 _18759_ (.X(_11908_),
    .B(_11907_),
    .A(net488));
 sg13g2_buf_1 _18760_ (.A(_11908_),
    .X(_11909_));
 sg13g2_mux2_1 _18761_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][4] ),
    .S(_11909_),
    .X(_11910_));
 sg13g2_mux2_1 _18762_ (.A0(_11910_),
    .A1(net989),
    .S(_11793_),
    .X(_00348_));
 sg13g2_mux2_1 _18763_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][5] ),
    .S(_11909_),
    .X(_11911_));
 sg13g2_mux2_1 _18764_ (.A0(_11911_),
    .A1(_11868_),
    .S(_11793_),
    .X(_00349_));
 sg13g2_mux2_1 _18765_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[0][6] ),
    .S(_11909_),
    .X(_11912_));
 sg13g2_mux2_1 _18766_ (.A0(_11912_),
    .A1(_11870_),
    .S(_11793_),
    .X(_00350_));
 sg13g2_mux2_1 _18767_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[0][7] ),
    .S(_11909_),
    .X(_11913_));
 sg13g2_mux2_1 _18768_ (.A0(_11913_),
    .A1(_09941_),
    .S(_11793_),
    .X(_00351_));
 sg13g2_mux2_1 _18769_ (.A0(net1081),
    .A1(\cpu.dcache.r_data[0][8] ),
    .S(_11799_),
    .X(_11914_));
 sg13g2_mux2_1 _18770_ (.A0(_11914_),
    .A1(net485),
    .S(net65),
    .X(_00352_));
 sg13g2_mux2_1 _18771_ (.A0(net1077),
    .A1(\cpu.dcache.r_data[0][9] ),
    .S(_11799_),
    .X(_11915_));
 sg13g2_mux2_1 _18772_ (.A0(_11915_),
    .A1(net484),
    .S(net65),
    .X(_00353_));
 sg13g2_nand2_1 _18773_ (.Y(_11916_),
    .A(_09251_),
    .B(_09270_));
 sg13g2_buf_1 _18774_ (.A(_11916_),
    .X(_11917_));
 sg13g2_buf_1 _18775_ (.A(_11917_),
    .X(_11918_));
 sg13g2_or2_1 _18776_ (.X(_11919_),
    .B(_11791_),
    .A(_11785_));
 sg13g2_buf_2 _18777_ (.A(_11919_),
    .X(_11920_));
 sg13g2_nor2_1 _18778_ (.A(net536),
    .B(_11920_),
    .Y(_11921_));
 sg13g2_buf_2 _18779_ (.A(_11921_),
    .X(_11922_));
 sg13g2_buf_1 _18780_ (.A(_11922_),
    .X(_11923_));
 sg13g2_buf_1 _18781_ (.A(_11760_),
    .X(_11924_));
 sg13g2_buf_2 _18782_ (.A(net1076),
    .X(_11925_));
 sg13g2_nor2_1 _18783_ (.A(net536),
    .B(_11774_),
    .Y(_11926_));
 sg13g2_buf_2 _18784_ (.A(_11926_),
    .X(_11927_));
 sg13g2_nor2b_1 _18785_ (.A(_11927_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_11928_));
 sg13g2_a21oi_1 _18786_ (.A1(net986),
    .A2(_11927_),
    .Y(_11929_),
    .B1(_11928_));
 sg13g2_buf_1 _18787_ (.A(net1020),
    .X(_11930_));
 sg13g2_nand2_1 _18788_ (.Y(_11931_),
    .A(_11930_),
    .B(net60));
 sg13g2_o21ai_1 _18789_ (.B1(_11931_),
    .Y(_00354_),
    .A1(net60),
    .A2(_11929_));
 sg13g2_or3_1 _18790_ (.A(_11785_),
    .B(_11789_),
    .C(_11808_),
    .X(_11932_));
 sg13g2_buf_2 _18791_ (.A(_11932_),
    .X(_11933_));
 sg13g2_nor2_1 _18792_ (.A(net536),
    .B(_11933_),
    .Y(_11934_));
 sg13g2_buf_1 _18793_ (.A(_11934_),
    .X(_11935_));
 sg13g2_buf_1 _18794_ (.A(_11935_),
    .X(_11936_));
 sg13g2_buf_1 _18795_ (.A(_11794_),
    .X(_11937_));
 sg13g2_buf_2 _18796_ (.A(net1075),
    .X(_11938_));
 sg13g2_nor2_1 _18797_ (.A(net536),
    .B(_11797_),
    .Y(_11939_));
 sg13g2_buf_2 _18798_ (.A(_11939_),
    .X(_11940_));
 sg13g2_nor2b_1 _18799_ (.A(_11940_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_11941_));
 sg13g2_a21oi_1 _18800_ (.A1(net985),
    .A2(_11940_),
    .Y(_11942_),
    .B1(_11941_));
 sg13g2_nand2_1 _18801_ (.Y(_11943_),
    .A(net487),
    .B(net59));
 sg13g2_o21ai_1 _18802_ (.B1(_11943_),
    .Y(_00355_),
    .A1(net59),
    .A2(_11942_));
 sg13g2_buf_1 _18803_ (.A(_11811_),
    .X(_11944_));
 sg13g2_buf_2 _18804_ (.A(net1074),
    .X(_11945_));
 sg13g2_nor2b_1 _18805_ (.A(_11940_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_11946_));
 sg13g2_a21oi_1 _18806_ (.A1(net984),
    .A2(_11940_),
    .Y(_11947_),
    .B1(_11946_));
 sg13g2_nand2_1 _18807_ (.Y(_11948_),
    .A(net486),
    .B(net59));
 sg13g2_o21ai_1 _18808_ (.B1(_11948_),
    .Y(_00356_),
    .A1(net59),
    .A2(_11947_));
 sg13g2_buf_1 _18809_ (.A(_11760_),
    .X(_11949_));
 sg13g2_nor2_2 _18810_ (.A(net536),
    .B(_11823_),
    .Y(_11950_));
 sg13g2_mux2_1 _18811_ (.A0(\cpu.dcache.r_data[1][12] ),
    .A1(net1073),
    .S(_11950_),
    .X(_11951_));
 sg13g2_nor2_1 _18812_ (.A(_11935_),
    .B(_11951_),
    .Y(_11952_));
 sg13g2_a21oi_1 _18813_ (.A1(net423),
    .A2(net59),
    .Y(_00357_),
    .B1(_11952_));
 sg13g2_buf_1 _18814_ (.A(_11831_),
    .X(_11953_));
 sg13g2_mux2_1 _18815_ (.A0(\cpu.dcache.r_data[1][13] ),
    .A1(net1072),
    .S(_11950_),
    .X(_11954_));
 sg13g2_nor2_1 _18816_ (.A(_11935_),
    .B(_11954_),
    .Y(_11955_));
 sg13g2_a21oi_1 _18817_ (.A1(_11895_),
    .A2(net59),
    .Y(_00358_),
    .B1(_11955_));
 sg13g2_buf_1 _18818_ (.A(_11794_),
    .X(_11956_));
 sg13g2_mux2_1 _18819_ (.A0(\cpu.dcache.r_data[1][14] ),
    .A1(net1071),
    .S(_11950_),
    .X(_11957_));
 sg13g2_nor2_1 _18820_ (.A(_11935_),
    .B(_11957_),
    .Y(_11958_));
 sg13g2_a21oi_1 _18821_ (.A1(net421),
    .A2(_11936_),
    .Y(_00359_),
    .B1(_11958_));
 sg13g2_buf_1 _18822_ (.A(_11811_),
    .X(_11959_));
 sg13g2_mux2_1 _18823_ (.A0(\cpu.dcache.r_data[1][15] ),
    .A1(net1070),
    .S(_11950_),
    .X(_11960_));
 sg13g2_nor2_1 _18824_ (.A(_11935_),
    .B(_11960_),
    .Y(_11961_));
 sg13g2_a21oi_1 _18825_ (.A1(net420),
    .A2(_11936_),
    .Y(_00360_),
    .B1(_11961_));
 sg13g2_or2_1 _18826_ (.X(_11962_),
    .B(_11851_),
    .A(_11785_));
 sg13g2_buf_2 _18827_ (.A(_11962_),
    .X(_11963_));
 sg13g2_nor2_1 _18828_ (.A(net536),
    .B(_11963_),
    .Y(_11964_));
 sg13g2_buf_2 _18829_ (.A(_11964_),
    .X(_11965_));
 sg13g2_buf_1 _18830_ (.A(_11965_),
    .X(_11966_));
 sg13g2_nor2_1 _18831_ (.A(net536),
    .B(_11846_),
    .Y(_11967_));
 sg13g2_buf_2 _18832_ (.A(_11967_),
    .X(_11968_));
 sg13g2_nor2b_1 _18833_ (.A(_11968_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_11969_));
 sg13g2_a21oi_1 _18834_ (.A1(net986),
    .A2(_11968_),
    .Y(_11970_),
    .B1(_11969_));
 sg13g2_buf_1 _18835_ (.A(net1020),
    .X(_11971_));
 sg13g2_nand2_1 _18836_ (.Y(_11972_),
    .A(net860),
    .B(net58));
 sg13g2_o21ai_1 _18837_ (.B1(_11972_),
    .Y(_00361_),
    .A1(net58),
    .A2(_11970_));
 sg13g2_buf_1 _18838_ (.A(_11831_),
    .X(_11973_));
 sg13g2_buf_2 _18839_ (.A(net1069),
    .X(_11974_));
 sg13g2_nor2b_1 _18840_ (.A(_11968_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_11975_));
 sg13g2_a21oi_1 _18841_ (.A1(net983),
    .A2(_11968_),
    .Y(_11976_),
    .B1(_11975_));
 sg13g2_buf_1 _18842_ (.A(net1019),
    .X(_11977_));
 sg13g2_nand2_1 _18843_ (.Y(_11978_),
    .A(net859),
    .B(net58));
 sg13g2_o21ai_1 _18844_ (.B1(_11978_),
    .Y(_00362_),
    .A1(net58),
    .A2(_11976_));
 sg13g2_nor2b_1 _18845_ (.A(_11968_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_11979_));
 sg13g2_a21oi_1 _18846_ (.A1(net985),
    .A2(_11968_),
    .Y(_11980_),
    .B1(_11979_));
 sg13g2_buf_1 _18847_ (.A(net1018),
    .X(_11981_));
 sg13g2_nand2_1 _18848_ (.Y(_11982_),
    .A(_11981_),
    .B(_11965_));
 sg13g2_o21ai_1 _18849_ (.B1(_11982_),
    .Y(_00363_),
    .A1(net58),
    .A2(_11980_));
 sg13g2_nor2b_1 _18850_ (.A(_11968_),
    .B_N(\cpu.dcache.r_data[1][19] ),
    .Y(_11983_));
 sg13g2_a21oi_1 _18851_ (.A1(net984),
    .A2(_11968_),
    .Y(_11984_),
    .B1(_11983_));
 sg13g2_buf_1 _18852_ (.A(net1098),
    .X(_11985_));
 sg13g2_nand2_1 _18853_ (.Y(_11986_),
    .A(net982),
    .B(_11965_));
 sg13g2_o21ai_1 _18854_ (.B1(_11986_),
    .Y(_00364_),
    .A1(net58),
    .A2(_11984_));
 sg13g2_nor2b_1 _18855_ (.A(_11927_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_11987_));
 sg13g2_a21oi_1 _18856_ (.A1(net983),
    .A2(_11927_),
    .Y(_11988_),
    .B1(_11987_));
 sg13g2_nand2_1 _18857_ (.Y(_11989_),
    .A(_11977_),
    .B(net60));
 sg13g2_o21ai_1 _18858_ (.B1(_11989_),
    .Y(_00365_),
    .A1(net60),
    .A2(_11988_));
 sg13g2_nor2_1 _18859_ (.A(_11917_),
    .B(_11862_),
    .Y(_11990_));
 sg13g2_buf_2 _18860_ (.A(_11990_),
    .X(_11991_));
 sg13g2_nor2b_1 _18861_ (.A(_11991_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_11992_));
 sg13g2_a21oi_1 _18862_ (.A1(net986),
    .A2(_11991_),
    .Y(_11993_),
    .B1(_11992_));
 sg13g2_buf_1 _18863_ (.A(_09921_),
    .X(_11994_));
 sg13g2_nand2_1 _18864_ (.Y(_11995_),
    .A(_11994_),
    .B(_11965_));
 sg13g2_o21ai_1 _18865_ (.B1(_11995_),
    .Y(_00366_),
    .A1(net58),
    .A2(_11993_));
 sg13g2_nor2b_1 _18866_ (.A(_11991_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_11996_));
 sg13g2_a21oi_1 _18867_ (.A1(net983),
    .A2(_11991_),
    .Y(_11997_),
    .B1(_11996_));
 sg13g2_buf_1 _18868_ (.A(_09927_),
    .X(_11998_));
 sg13g2_nand2_1 _18869_ (.Y(_11999_),
    .A(net980),
    .B(_11965_));
 sg13g2_o21ai_1 _18870_ (.B1(_11999_),
    .Y(_00367_),
    .A1(net58),
    .A2(_11997_));
 sg13g2_nor2b_1 _18871_ (.A(_11991_),
    .B_N(\cpu.dcache.r_data[1][22] ),
    .Y(_12000_));
 sg13g2_a21oi_1 _18872_ (.A1(net985),
    .A2(_11991_),
    .Y(_12001_),
    .B1(_12000_));
 sg13g2_buf_1 _18873_ (.A(_09933_),
    .X(_12002_));
 sg13g2_nand2_1 _18874_ (.Y(_12003_),
    .A(net979),
    .B(_11965_));
 sg13g2_o21ai_1 _18875_ (.B1(_12003_),
    .Y(_00368_),
    .A1(_11966_),
    .A2(_12001_));
 sg13g2_nor2b_1 _18876_ (.A(_11991_),
    .B_N(\cpu.dcache.r_data[1][23] ),
    .Y(_12004_));
 sg13g2_a21oi_1 _18877_ (.A1(net984),
    .A2(_11991_),
    .Y(_12005_),
    .B1(_12004_));
 sg13g2_buf_1 _18878_ (.A(_09940_),
    .X(_12006_));
 sg13g2_nand2_1 _18879_ (.Y(_12007_),
    .A(_12006_),
    .B(_11965_));
 sg13g2_o21ai_1 _18880_ (.B1(_12007_),
    .Y(_00369_),
    .A1(_11966_),
    .A2(_12005_));
 sg13g2_or3_1 _18881_ (.A(_11785_),
    .B(_11789_),
    .C(_11879_),
    .X(_12008_));
 sg13g2_buf_2 _18882_ (.A(_12008_),
    .X(_12009_));
 sg13g2_nor2_1 _18883_ (.A(_11918_),
    .B(_12009_),
    .Y(_12010_));
 sg13g2_buf_1 _18884_ (.A(_12010_),
    .X(_12011_));
 sg13g2_buf_1 _18885_ (.A(_12011_),
    .X(_12012_));
 sg13g2_buf_1 _18886_ (.A(net1080),
    .X(_12013_));
 sg13g2_nand3_1 _18887_ (.B(_11766_),
    .C(net863),
    .A(net977),
    .Y(_12014_));
 sg13g2_buf_1 _18888_ (.A(_12014_),
    .X(_12015_));
 sg13g2_nor2_1 _18889_ (.A(_11917_),
    .B(_12015_),
    .Y(_12016_));
 sg13g2_buf_1 _18890_ (.A(_12016_),
    .X(_12017_));
 sg13g2_nor2b_1 _18891_ (.A(net483),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12018_));
 sg13g2_a21oi_1 _18892_ (.A1(net986),
    .A2(net483),
    .Y(_12019_),
    .B1(_12018_));
 sg13g2_nand2_1 _18893_ (.Y(_12020_),
    .A(net485),
    .B(_12012_));
 sg13g2_o21ai_1 _18894_ (.B1(_12020_),
    .Y(_00370_),
    .A1(net57),
    .A2(_12019_));
 sg13g2_nor2b_1 _18895_ (.A(net483),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12021_));
 sg13g2_a21oi_1 _18896_ (.A1(net983),
    .A2(net483),
    .Y(_12022_),
    .B1(_12021_));
 sg13g2_nand2_1 _18897_ (.Y(_12023_),
    .A(_11885_),
    .B(net57));
 sg13g2_o21ai_1 _18898_ (.B1(_12023_),
    .Y(_00371_),
    .A1(net57),
    .A2(_12022_));
 sg13g2_nor2b_1 _18899_ (.A(net483),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12024_));
 sg13g2_a21oi_1 _18900_ (.A1(net985),
    .A2(net483),
    .Y(_12025_),
    .B1(_12024_));
 sg13g2_nand2_1 _18901_ (.Y(_12026_),
    .A(net487),
    .B(_12011_));
 sg13g2_o21ai_1 _18902_ (.B1(_12026_),
    .Y(_00372_),
    .A1(net57),
    .A2(_12025_));
 sg13g2_nor2b_1 _18903_ (.A(net483),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12027_));
 sg13g2_a21oi_1 _18904_ (.A1(net984),
    .A2(_12017_),
    .Y(_12028_),
    .B1(_12027_));
 sg13g2_nand2_1 _18905_ (.Y(_12029_),
    .A(net486),
    .B(_12011_));
 sg13g2_o21ai_1 _18906_ (.B1(_12029_),
    .Y(_00373_),
    .A1(_12012_),
    .A2(_12028_));
 sg13g2_nor2_2 _18907_ (.A(_11918_),
    .B(_11890_),
    .Y(_12030_));
 sg13g2_mux2_1 _18908_ (.A0(\cpu.dcache.r_data[1][28] ),
    .A1(net1073),
    .S(_12030_),
    .X(_12031_));
 sg13g2_nor2_1 _18909_ (.A(_12011_),
    .B(_12031_),
    .Y(_12032_));
 sg13g2_a21oi_1 _18910_ (.A1(net423),
    .A2(net57),
    .Y(_00374_),
    .B1(_12032_));
 sg13g2_mux2_1 _18911_ (.A0(\cpu.dcache.r_data[1][29] ),
    .A1(_11953_),
    .S(_12030_),
    .X(_12033_));
 sg13g2_nor2_1 _18912_ (.A(_12011_),
    .B(_12033_),
    .Y(_12034_));
 sg13g2_a21oi_1 _18913_ (.A1(net422),
    .A2(net57),
    .Y(_00375_),
    .B1(_12034_));
 sg13g2_nor2b_1 _18914_ (.A(_11927_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_12035_));
 sg13g2_a21oi_1 _18915_ (.A1(net985),
    .A2(_11927_),
    .Y(_12036_),
    .B1(_12035_));
 sg13g2_nand2_1 _18916_ (.Y(_12037_),
    .A(_11981_),
    .B(_11922_));
 sg13g2_o21ai_1 _18917_ (.B1(_12037_),
    .Y(_00376_),
    .A1(net60),
    .A2(_12036_));
 sg13g2_mux2_1 _18918_ (.A0(\cpu.dcache.r_data[1][30] ),
    .A1(net1071),
    .S(_12030_),
    .X(_12038_));
 sg13g2_nor2_1 _18919_ (.A(_12011_),
    .B(_12038_),
    .Y(_12039_));
 sg13g2_a21oi_1 _18920_ (.A1(net421),
    .A2(net57),
    .Y(_00377_),
    .B1(_12039_));
 sg13g2_mux2_1 _18921_ (.A0(\cpu.dcache.r_data[1][31] ),
    .A1(net1070),
    .S(_12030_),
    .X(_12040_));
 sg13g2_nor2_1 _18922_ (.A(_12011_),
    .B(_12040_),
    .Y(_12041_));
 sg13g2_a21oi_1 _18923_ (.A1(net420),
    .A2(net57),
    .Y(_00378_),
    .B1(_12041_));
 sg13g2_nor2b_1 _18924_ (.A(_11927_),
    .B_N(\cpu.dcache.r_data[1][3] ),
    .Y(_12042_));
 sg13g2_a21oi_1 _18925_ (.A1(net984),
    .A2(_11927_),
    .Y(_12043_),
    .B1(_12042_));
 sg13g2_nand2_1 _18926_ (.Y(_12044_),
    .A(net982),
    .B(_11922_));
 sg13g2_o21ai_1 _18927_ (.B1(_12044_),
    .Y(_00379_),
    .A1(_11923_),
    .A2(_12043_));
 sg13g2_nor2_1 _18928_ (.A(_11917_),
    .B(_11907_),
    .Y(_12045_));
 sg13g2_buf_2 _18929_ (.A(_12045_),
    .X(_12046_));
 sg13g2_nor2b_1 _18930_ (.A(_12046_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_12047_));
 sg13g2_a21oi_1 _18931_ (.A1(net986),
    .A2(_12046_),
    .Y(_12048_),
    .B1(_12047_));
 sg13g2_nand2_1 _18932_ (.Y(_12049_),
    .A(net981),
    .B(_11922_));
 sg13g2_o21ai_1 _18933_ (.B1(_12049_),
    .Y(_00380_),
    .A1(net60),
    .A2(_12048_));
 sg13g2_nor2b_1 _18934_ (.A(_12046_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_12050_));
 sg13g2_a21oi_1 _18935_ (.A1(net983),
    .A2(_12046_),
    .Y(_12051_),
    .B1(_12050_));
 sg13g2_nand2_1 _18936_ (.Y(_12052_),
    .A(_11998_),
    .B(_11922_));
 sg13g2_o21ai_1 _18937_ (.B1(_12052_),
    .Y(_00381_),
    .A1(net60),
    .A2(_12051_));
 sg13g2_nor2b_1 _18938_ (.A(_12046_),
    .B_N(\cpu.dcache.r_data[1][6] ),
    .Y(_12053_));
 sg13g2_a21oi_1 _18939_ (.A1(net985),
    .A2(_12046_),
    .Y(_12054_),
    .B1(_12053_));
 sg13g2_nand2_1 _18940_ (.Y(_12055_),
    .A(_12002_),
    .B(_11922_));
 sg13g2_o21ai_1 _18941_ (.B1(_12055_),
    .Y(_00382_),
    .A1(net60),
    .A2(_12054_));
 sg13g2_nor2b_1 _18942_ (.A(_12046_),
    .B_N(\cpu.dcache.r_data[1][7] ),
    .Y(_12056_));
 sg13g2_a21oi_1 _18943_ (.A1(net984),
    .A2(_12046_),
    .Y(_12057_),
    .B1(_12056_));
 sg13g2_buf_1 _18944_ (.A(_09940_),
    .X(_12058_));
 sg13g2_nand2_1 _18945_ (.Y(_12059_),
    .A(net976),
    .B(_11922_));
 sg13g2_o21ai_1 _18946_ (.B1(_12059_),
    .Y(_00383_),
    .A1(_11923_),
    .A2(_12057_));
 sg13g2_nor2b_1 _18947_ (.A(_11940_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12060_));
 sg13g2_a21oi_1 _18948_ (.A1(net986),
    .A2(_11940_),
    .Y(_12061_),
    .B1(_12060_));
 sg13g2_nand2_1 _18949_ (.Y(_12062_),
    .A(net485),
    .B(_11935_));
 sg13g2_o21ai_1 _18950_ (.B1(_12062_),
    .Y(_00384_),
    .A1(net59),
    .A2(_12061_));
 sg13g2_nor2b_1 _18951_ (.A(_11940_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12063_));
 sg13g2_a21oi_1 _18952_ (.A1(net983),
    .A2(_11940_),
    .Y(_12064_),
    .B1(_12063_));
 sg13g2_nand2_1 _18953_ (.Y(_12065_),
    .A(net484),
    .B(_11935_));
 sg13g2_o21ai_1 _18954_ (.B1(_12065_),
    .Y(_00385_),
    .A1(net59),
    .A2(_12064_));
 sg13g2_nand2_1 _18955_ (.Y(_12066_),
    .A(net1025),
    .B(net894));
 sg13g2_buf_1 _18956_ (.A(_12066_),
    .X(_12067_));
 sg13g2_buf_1 _18957_ (.A(_12067_),
    .X(_12068_));
 sg13g2_nor2_1 _18958_ (.A(net600),
    .B(_11920_),
    .Y(_12069_));
 sg13g2_buf_2 _18959_ (.A(_12069_),
    .X(_12070_));
 sg13g2_buf_1 _18960_ (.A(_12070_),
    .X(_12071_));
 sg13g2_buf_1 _18961_ (.A(net1076),
    .X(_12072_));
 sg13g2_nor2_1 _18962_ (.A(net600),
    .B(_11774_),
    .Y(_12073_));
 sg13g2_buf_2 _18963_ (.A(_12073_),
    .X(_12074_));
 sg13g2_nor2b_1 _18964_ (.A(_12074_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12075_));
 sg13g2_a21oi_1 _18965_ (.A1(net975),
    .A2(_12074_),
    .Y(_12076_),
    .B1(_12075_));
 sg13g2_nand2_1 _18966_ (.Y(_12077_),
    .A(_11971_),
    .B(net56));
 sg13g2_o21ai_1 _18967_ (.B1(_12077_),
    .Y(_00386_),
    .A1(net56),
    .A2(_12076_));
 sg13g2_nor2_1 _18968_ (.A(net600),
    .B(_11933_),
    .Y(_12078_));
 sg13g2_buf_1 _18969_ (.A(_12078_),
    .X(_12079_));
 sg13g2_buf_1 _18970_ (.A(_12079_),
    .X(_12080_));
 sg13g2_buf_1 _18971_ (.A(net1075),
    .X(_12081_));
 sg13g2_nor2_1 _18972_ (.A(net600),
    .B(_11797_),
    .Y(_12082_));
 sg13g2_buf_2 _18973_ (.A(_12082_),
    .X(_12083_));
 sg13g2_nor2b_1 _18974_ (.A(_12083_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12084_));
 sg13g2_a21oi_1 _18975_ (.A1(net974),
    .A2(_12083_),
    .Y(_12085_),
    .B1(_12084_));
 sg13g2_nand2_1 _18976_ (.Y(_12086_),
    .A(net487),
    .B(net55));
 sg13g2_o21ai_1 _18977_ (.B1(_12086_),
    .Y(_00387_),
    .A1(net55),
    .A2(_12085_));
 sg13g2_buf_1 _18978_ (.A(net1074),
    .X(_12087_));
 sg13g2_nor2b_1 _18979_ (.A(_12083_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12088_));
 sg13g2_a21oi_1 _18980_ (.A1(net973),
    .A2(_12083_),
    .Y(_12089_),
    .B1(_12088_));
 sg13g2_nand2_1 _18981_ (.Y(_12090_),
    .A(net486),
    .B(net55));
 sg13g2_o21ai_1 _18982_ (.B1(_12090_),
    .Y(_00388_),
    .A1(net55),
    .A2(_12089_));
 sg13g2_nor2_2 _18983_ (.A(net600),
    .B(_11823_),
    .Y(_12091_));
 sg13g2_mux2_1 _18984_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(net1073),
    .S(_12091_),
    .X(_12092_));
 sg13g2_nor2_1 _18985_ (.A(_12079_),
    .B(_12092_),
    .Y(_12093_));
 sg13g2_a21oi_1 _18986_ (.A1(net423),
    .A2(net55),
    .Y(_00389_),
    .B1(_12093_));
 sg13g2_mux2_1 _18987_ (.A0(\cpu.dcache.r_data[2][13] ),
    .A1(net1072),
    .S(_12091_),
    .X(_12094_));
 sg13g2_nor2_1 _18988_ (.A(_12079_),
    .B(_12094_),
    .Y(_12095_));
 sg13g2_a21oi_1 _18989_ (.A1(net422),
    .A2(net55),
    .Y(_00390_),
    .B1(_12095_));
 sg13g2_mux2_1 _18990_ (.A0(\cpu.dcache.r_data[2][14] ),
    .A1(net1071),
    .S(_12091_),
    .X(_12096_));
 sg13g2_nor2_1 _18991_ (.A(_12079_),
    .B(_12096_),
    .Y(_12097_));
 sg13g2_a21oi_1 _18992_ (.A1(net421),
    .A2(_12080_),
    .Y(_00391_),
    .B1(_12097_));
 sg13g2_mux2_1 _18993_ (.A0(\cpu.dcache.r_data[2][15] ),
    .A1(net1070),
    .S(_12091_),
    .X(_12098_));
 sg13g2_nor2_1 _18994_ (.A(_12079_),
    .B(_12098_),
    .Y(_12099_));
 sg13g2_a21oi_1 _18995_ (.A1(net420),
    .A2(net55),
    .Y(_00392_),
    .B1(_12099_));
 sg13g2_nor2_1 _18996_ (.A(net600),
    .B(_11963_),
    .Y(_12100_));
 sg13g2_buf_2 _18997_ (.A(_12100_),
    .X(_12101_));
 sg13g2_buf_1 _18998_ (.A(_12101_),
    .X(_12102_));
 sg13g2_nor2_1 _18999_ (.A(net600),
    .B(_11846_),
    .Y(_12103_));
 sg13g2_buf_2 _19000_ (.A(_12103_),
    .X(_12104_));
 sg13g2_nor2b_1 _19001_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12105_));
 sg13g2_a21oi_1 _19002_ (.A1(net975),
    .A2(_12104_),
    .Y(_12106_),
    .B1(_12105_));
 sg13g2_nand2_1 _19003_ (.Y(_12107_),
    .A(net860),
    .B(_12102_));
 sg13g2_o21ai_1 _19004_ (.B1(_12107_),
    .Y(_00393_),
    .A1(_12102_),
    .A2(_12106_));
 sg13g2_buf_1 _19005_ (.A(net1069),
    .X(_12108_));
 sg13g2_nor2b_1 _19006_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12109_));
 sg13g2_a21oi_1 _19007_ (.A1(net972),
    .A2(_12104_),
    .Y(_12110_),
    .B1(_12109_));
 sg13g2_nand2_1 _19008_ (.Y(_12111_),
    .A(_11977_),
    .B(net54));
 sg13g2_o21ai_1 _19009_ (.B1(_12111_),
    .Y(_00394_),
    .A1(net54),
    .A2(_12110_));
 sg13g2_nor2b_1 _19010_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12112_));
 sg13g2_a21oi_1 _19011_ (.A1(net974),
    .A2(_12104_),
    .Y(_12113_),
    .B1(_12112_));
 sg13g2_nand2_1 _19012_ (.Y(_12114_),
    .A(net858),
    .B(_12101_));
 sg13g2_o21ai_1 _19013_ (.B1(_12114_),
    .Y(_00395_),
    .A1(net54),
    .A2(_12113_));
 sg13g2_nor2b_1 _19014_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[2][19] ),
    .Y(_12115_));
 sg13g2_a21oi_1 _19015_ (.A1(net973),
    .A2(_12104_),
    .Y(_12116_),
    .B1(_12115_));
 sg13g2_nand2_1 _19016_ (.Y(_12117_),
    .A(net982),
    .B(_12101_));
 sg13g2_o21ai_1 _19017_ (.B1(_12117_),
    .Y(_00396_),
    .A1(net54),
    .A2(_12116_));
 sg13g2_nor2b_1 _19018_ (.A(_12074_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12118_));
 sg13g2_a21oi_1 _19019_ (.A1(net972),
    .A2(_12074_),
    .Y(_12119_),
    .B1(_12118_));
 sg13g2_buf_1 _19020_ (.A(net1019),
    .X(_12120_));
 sg13g2_nand2_1 _19021_ (.Y(_12121_),
    .A(net857),
    .B(_12071_));
 sg13g2_o21ai_1 _19022_ (.B1(_12121_),
    .Y(_00397_),
    .A1(_12071_),
    .A2(_12119_));
 sg13g2_nor2_1 _19023_ (.A(_12067_),
    .B(_11862_),
    .Y(_12122_));
 sg13g2_buf_2 _19024_ (.A(_12122_),
    .X(_12123_));
 sg13g2_nor2b_1 _19025_ (.A(_12123_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12124_));
 sg13g2_a21oi_1 _19026_ (.A1(net975),
    .A2(_12123_),
    .Y(_12125_),
    .B1(_12124_));
 sg13g2_nand2_1 _19027_ (.Y(_12126_),
    .A(_11994_),
    .B(_12101_));
 sg13g2_o21ai_1 _19028_ (.B1(_12126_),
    .Y(_00398_),
    .A1(net54),
    .A2(_12125_));
 sg13g2_nor2b_1 _19029_ (.A(_12123_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12127_));
 sg13g2_a21oi_1 _19030_ (.A1(net972),
    .A2(_12123_),
    .Y(_12128_),
    .B1(_12127_));
 sg13g2_nand2_1 _19031_ (.Y(_12129_),
    .A(_11998_),
    .B(_12101_));
 sg13g2_o21ai_1 _19032_ (.B1(_12129_),
    .Y(_00399_),
    .A1(net54),
    .A2(_12128_));
 sg13g2_nor2b_1 _19033_ (.A(_12123_),
    .B_N(\cpu.dcache.r_data[2][22] ),
    .Y(_12130_));
 sg13g2_a21oi_1 _19034_ (.A1(net974),
    .A2(_12123_),
    .Y(_12131_),
    .B1(_12130_));
 sg13g2_nand2_1 _19035_ (.Y(_12132_),
    .A(net979),
    .B(_12101_));
 sg13g2_o21ai_1 _19036_ (.B1(_12132_),
    .Y(_00400_),
    .A1(net54),
    .A2(_12131_));
 sg13g2_nor2b_1 _19037_ (.A(_12123_),
    .B_N(\cpu.dcache.r_data[2][23] ),
    .Y(_12133_));
 sg13g2_a21oi_1 _19038_ (.A1(net973),
    .A2(_12123_),
    .Y(_12134_),
    .B1(_12133_));
 sg13g2_nand2_1 _19039_ (.Y(_12135_),
    .A(net976),
    .B(_12101_));
 sg13g2_o21ai_1 _19040_ (.B1(_12135_),
    .Y(_00401_),
    .A1(net54),
    .A2(_12134_));
 sg13g2_nor2_1 _19041_ (.A(_12068_),
    .B(_12009_),
    .Y(_12136_));
 sg13g2_buf_1 _19042_ (.A(_12136_),
    .X(_12137_));
 sg13g2_buf_1 _19043_ (.A(_12137_),
    .X(_12138_));
 sg13g2_nor2_1 _19044_ (.A(_12067_),
    .B(_12015_),
    .Y(_12139_));
 sg13g2_buf_1 _19045_ (.A(_12139_),
    .X(_12140_));
 sg13g2_nor2b_1 _19046_ (.A(_12140_),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12141_));
 sg13g2_a21oi_1 _19047_ (.A1(_12072_),
    .A2(_12140_),
    .Y(_12142_),
    .B1(_12141_));
 sg13g2_nand2_1 _19048_ (.Y(_12143_),
    .A(_11877_),
    .B(net53));
 sg13g2_o21ai_1 _19049_ (.B1(_12143_),
    .Y(_00402_),
    .A1(_12138_),
    .A2(_12142_));
 sg13g2_nor2b_1 _19050_ (.A(net535),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12144_));
 sg13g2_a21oi_1 _19051_ (.A1(net972),
    .A2(net535),
    .Y(_12145_),
    .B1(_12144_));
 sg13g2_nand2_1 _19052_ (.Y(_12146_),
    .A(net484),
    .B(net53));
 sg13g2_o21ai_1 _19053_ (.B1(_12146_),
    .Y(_00403_),
    .A1(net53),
    .A2(_12145_));
 sg13g2_nor2b_1 _19054_ (.A(net535),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12147_));
 sg13g2_a21oi_1 _19055_ (.A1(_12081_),
    .A2(net535),
    .Y(_12148_),
    .B1(_12147_));
 sg13g2_nand2_1 _19056_ (.Y(_12149_),
    .A(_11806_),
    .B(_12137_));
 sg13g2_o21ai_1 _19057_ (.B1(_12149_),
    .Y(_00404_),
    .A1(net53),
    .A2(_12148_));
 sg13g2_nor2b_1 _19058_ (.A(net535),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12150_));
 sg13g2_a21oi_1 _19059_ (.A1(_12087_),
    .A2(net535),
    .Y(_12151_),
    .B1(_12150_));
 sg13g2_nand2_1 _19060_ (.Y(_12152_),
    .A(_11816_),
    .B(_12137_));
 sg13g2_o21ai_1 _19061_ (.B1(_12152_),
    .Y(_00405_),
    .A1(_12138_),
    .A2(_12151_));
 sg13g2_nor2_2 _19062_ (.A(_12068_),
    .B(_11890_),
    .Y(_12153_));
 sg13g2_mux2_1 _19063_ (.A0(\cpu.dcache.r_data[2][28] ),
    .A1(net1073),
    .S(_12153_),
    .X(_12154_));
 sg13g2_nor2_1 _19064_ (.A(_12137_),
    .B(_12154_),
    .Y(_12155_));
 sg13g2_a21oi_1 _19065_ (.A1(net423),
    .A2(net53),
    .Y(_00406_),
    .B1(_12155_));
 sg13g2_mux2_1 _19066_ (.A0(\cpu.dcache.r_data[2][29] ),
    .A1(_11953_),
    .S(_12153_),
    .X(_12156_));
 sg13g2_nor2_1 _19067_ (.A(_12137_),
    .B(_12156_),
    .Y(_12157_));
 sg13g2_a21oi_1 _19068_ (.A1(net422),
    .A2(net53),
    .Y(_00407_),
    .B1(_12157_));
 sg13g2_nor2b_1 _19069_ (.A(_12074_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12158_));
 sg13g2_a21oi_1 _19070_ (.A1(net974),
    .A2(_12074_),
    .Y(_12159_),
    .B1(_12158_));
 sg13g2_buf_1 _19071_ (.A(net1018),
    .X(_12160_));
 sg13g2_nand2_1 _19072_ (.Y(_12161_),
    .A(net856),
    .B(_12070_));
 sg13g2_o21ai_1 _19073_ (.B1(_12161_),
    .Y(_00408_),
    .A1(net56),
    .A2(_12159_));
 sg13g2_mux2_1 _19074_ (.A0(\cpu.dcache.r_data[2][30] ),
    .A1(net1071),
    .S(_12153_),
    .X(_12162_));
 sg13g2_nor2_1 _19075_ (.A(_12137_),
    .B(_12162_),
    .Y(_12163_));
 sg13g2_a21oi_1 _19076_ (.A1(net421),
    .A2(net53),
    .Y(_00409_),
    .B1(_12163_));
 sg13g2_mux2_1 _19077_ (.A0(\cpu.dcache.r_data[2][31] ),
    .A1(net1070),
    .S(_12153_),
    .X(_12164_));
 sg13g2_nor2_1 _19078_ (.A(_12137_),
    .B(_12164_),
    .Y(_12165_));
 sg13g2_a21oi_1 _19079_ (.A1(_11902_),
    .A2(net53),
    .Y(_00410_),
    .B1(_12165_));
 sg13g2_nor2b_1 _19080_ (.A(_12074_),
    .B_N(\cpu.dcache.r_data[2][3] ),
    .Y(_12166_));
 sg13g2_a21oi_1 _19081_ (.A1(net973),
    .A2(_12074_),
    .Y(_12167_),
    .B1(_12166_));
 sg13g2_nand2_1 _19082_ (.Y(_12168_),
    .A(net982),
    .B(_12070_));
 sg13g2_o21ai_1 _19083_ (.B1(_12168_),
    .Y(_00411_),
    .A1(net56),
    .A2(_12167_));
 sg13g2_nor2_1 _19084_ (.A(_12067_),
    .B(_11907_),
    .Y(_12169_));
 sg13g2_buf_2 _19085_ (.A(_12169_),
    .X(_12170_));
 sg13g2_nor2b_1 _19086_ (.A(_12170_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12171_));
 sg13g2_a21oi_1 _19087_ (.A1(net975),
    .A2(_12170_),
    .Y(_12172_),
    .B1(_12171_));
 sg13g2_buf_1 _19088_ (.A(_09921_),
    .X(_12173_));
 sg13g2_nand2_1 _19089_ (.Y(_12174_),
    .A(net971),
    .B(_12070_));
 sg13g2_o21ai_1 _19090_ (.B1(_12174_),
    .Y(_00412_),
    .A1(net56),
    .A2(_12172_));
 sg13g2_nor2b_1 _19091_ (.A(_12170_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12175_));
 sg13g2_a21oi_1 _19092_ (.A1(net972),
    .A2(_12170_),
    .Y(_12176_),
    .B1(_12175_));
 sg13g2_buf_1 _19093_ (.A(_09927_),
    .X(_12177_));
 sg13g2_nand2_1 _19094_ (.Y(_12178_),
    .A(net970),
    .B(_12070_));
 sg13g2_o21ai_1 _19095_ (.B1(_12178_),
    .Y(_00413_),
    .A1(net56),
    .A2(_12176_));
 sg13g2_nor2b_1 _19096_ (.A(_12170_),
    .B_N(\cpu.dcache.r_data[2][6] ),
    .Y(_12179_));
 sg13g2_a21oi_1 _19097_ (.A1(net974),
    .A2(_12170_),
    .Y(_12180_),
    .B1(_12179_));
 sg13g2_buf_1 _19098_ (.A(_09933_),
    .X(_12181_));
 sg13g2_nand2_1 _19099_ (.Y(_12182_),
    .A(net969),
    .B(_12070_));
 sg13g2_o21ai_1 _19100_ (.B1(_12182_),
    .Y(_00414_),
    .A1(net56),
    .A2(_12180_));
 sg13g2_nor2b_1 _19101_ (.A(_12170_),
    .B_N(\cpu.dcache.r_data[2][7] ),
    .Y(_12183_));
 sg13g2_a21oi_1 _19102_ (.A1(net973),
    .A2(_12170_),
    .Y(_12184_),
    .B1(_12183_));
 sg13g2_nand2_1 _19103_ (.Y(_12185_),
    .A(net976),
    .B(_12070_));
 sg13g2_o21ai_1 _19104_ (.B1(_12185_),
    .Y(_00415_),
    .A1(net56),
    .A2(_12184_));
 sg13g2_nor2b_1 _19105_ (.A(_12083_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12186_));
 sg13g2_a21oi_1 _19106_ (.A1(net975),
    .A2(_12083_),
    .Y(_12187_),
    .B1(_12186_));
 sg13g2_nand2_1 _19107_ (.Y(_12188_),
    .A(net485),
    .B(_12079_));
 sg13g2_o21ai_1 _19108_ (.B1(_12188_),
    .Y(_00416_),
    .A1(_12080_),
    .A2(_12187_));
 sg13g2_nor2b_1 _19109_ (.A(_12083_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12189_));
 sg13g2_a21oi_1 _19110_ (.A1(_12108_),
    .A2(_12083_),
    .Y(_12190_),
    .B1(_12189_));
 sg13g2_nand2_1 _19111_ (.Y(_12191_),
    .A(net484),
    .B(_12079_));
 sg13g2_o21ai_1 _19112_ (.B1(_12191_),
    .Y(_00417_),
    .A1(net55),
    .A2(_12190_));
 sg13g2_nand2_1 _19113_ (.Y(_12192_),
    .A(net1025),
    .B(net669));
 sg13g2_buf_1 _19114_ (.A(_12192_),
    .X(_12193_));
 sg13g2_buf_1 _19115_ (.A(_12193_),
    .X(_12194_));
 sg13g2_nor2_1 _19116_ (.A(net482),
    .B(_11920_),
    .Y(_12195_));
 sg13g2_buf_2 _19117_ (.A(_12195_),
    .X(_12196_));
 sg13g2_buf_1 _19118_ (.A(_12196_),
    .X(_12197_));
 sg13g2_nor2_1 _19119_ (.A(net482),
    .B(_11774_),
    .Y(_12198_));
 sg13g2_buf_2 _19120_ (.A(_12198_),
    .X(_12199_));
 sg13g2_nor2b_1 _19121_ (.A(_12199_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12200_));
 sg13g2_a21oi_1 _19122_ (.A1(net975),
    .A2(_12199_),
    .Y(_12201_),
    .B1(_12200_));
 sg13g2_nand2_1 _19123_ (.Y(_12202_),
    .A(net860),
    .B(_12197_));
 sg13g2_o21ai_1 _19124_ (.B1(_12202_),
    .Y(_00418_),
    .A1(net52),
    .A2(_12201_));
 sg13g2_nor2_1 _19125_ (.A(net482),
    .B(_11933_),
    .Y(_12203_));
 sg13g2_buf_2 _19126_ (.A(_12203_),
    .X(_12204_));
 sg13g2_buf_1 _19127_ (.A(_12204_),
    .X(_12205_));
 sg13g2_nor2_1 _19128_ (.A(net482),
    .B(_11797_),
    .Y(_12206_));
 sg13g2_buf_2 _19129_ (.A(_12206_),
    .X(_12207_));
 sg13g2_nor2b_1 _19130_ (.A(_12207_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12208_));
 sg13g2_a21oi_1 _19131_ (.A1(net974),
    .A2(_12207_),
    .Y(_12209_),
    .B1(_12208_));
 sg13g2_nand2_1 _19132_ (.Y(_12210_),
    .A(net487),
    .B(net51));
 sg13g2_o21ai_1 _19133_ (.B1(_12210_),
    .Y(_00419_),
    .A1(net51),
    .A2(_12209_));
 sg13g2_nor2b_1 _19134_ (.A(_12207_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12211_));
 sg13g2_a21oi_1 _19135_ (.A1(net973),
    .A2(_12207_),
    .Y(_12212_),
    .B1(_12211_));
 sg13g2_nand2_1 _19136_ (.Y(_12213_),
    .A(net486),
    .B(net51));
 sg13g2_o21ai_1 _19137_ (.B1(_12213_),
    .Y(_00420_),
    .A1(net51),
    .A2(_12212_));
 sg13g2_nor2_2 _19138_ (.A(net482),
    .B(_11823_),
    .Y(_12214_));
 sg13g2_mux2_1 _19139_ (.A0(\cpu.dcache.r_data[3][12] ),
    .A1(net1073),
    .S(_12214_),
    .X(_12215_));
 sg13g2_nor2_1 _19140_ (.A(_12204_),
    .B(_12215_),
    .Y(_12216_));
 sg13g2_a21oi_1 _19141_ (.A1(net423),
    .A2(net51),
    .Y(_00421_),
    .B1(_12216_));
 sg13g2_mux2_1 _19142_ (.A0(\cpu.dcache.r_data[3][13] ),
    .A1(net1072),
    .S(_12214_),
    .X(_12217_));
 sg13g2_nor2_1 _19143_ (.A(_12204_),
    .B(_12217_),
    .Y(_12218_));
 sg13g2_a21oi_1 _19144_ (.A1(net422),
    .A2(net51),
    .Y(_00422_),
    .B1(_12218_));
 sg13g2_mux2_1 _19145_ (.A0(\cpu.dcache.r_data[3][14] ),
    .A1(net1071),
    .S(_12214_),
    .X(_12219_));
 sg13g2_nor2_1 _19146_ (.A(_12204_),
    .B(_12219_),
    .Y(_12220_));
 sg13g2_a21oi_1 _19147_ (.A1(net421),
    .A2(_12205_),
    .Y(_00423_),
    .B1(_12220_));
 sg13g2_mux2_1 _19148_ (.A0(\cpu.dcache.r_data[3][15] ),
    .A1(net1070),
    .S(_12214_),
    .X(_12221_));
 sg13g2_nor2_1 _19149_ (.A(_12204_),
    .B(_12221_),
    .Y(_12222_));
 sg13g2_a21oi_1 _19150_ (.A1(net420),
    .A2(_12205_),
    .Y(_00424_),
    .B1(_12222_));
 sg13g2_nor2_1 _19151_ (.A(net482),
    .B(_11963_),
    .Y(_12223_));
 sg13g2_buf_2 _19152_ (.A(_12223_),
    .X(_12224_));
 sg13g2_buf_1 _19153_ (.A(_12224_),
    .X(_12225_));
 sg13g2_nor2_1 _19154_ (.A(net482),
    .B(_11846_),
    .Y(_12226_));
 sg13g2_buf_2 _19155_ (.A(_12226_),
    .X(_12227_));
 sg13g2_nor2b_1 _19156_ (.A(_12227_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12228_));
 sg13g2_a21oi_1 _19157_ (.A1(net975),
    .A2(_12227_),
    .Y(_12229_),
    .B1(_12228_));
 sg13g2_nand2_1 _19158_ (.Y(_12230_),
    .A(net860),
    .B(net50));
 sg13g2_o21ai_1 _19159_ (.B1(_12230_),
    .Y(_00425_),
    .A1(net50),
    .A2(_12229_));
 sg13g2_nor2b_1 _19160_ (.A(_12227_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12231_));
 sg13g2_a21oi_1 _19161_ (.A1(net972),
    .A2(_12227_),
    .Y(_12232_),
    .B1(_12231_));
 sg13g2_nand2_1 _19162_ (.Y(_12233_),
    .A(net857),
    .B(net50));
 sg13g2_o21ai_1 _19163_ (.B1(_12233_),
    .Y(_00426_),
    .A1(net50),
    .A2(_12232_));
 sg13g2_nor2b_1 _19164_ (.A(_12227_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12234_));
 sg13g2_a21oi_1 _19165_ (.A1(net974),
    .A2(_12227_),
    .Y(_12235_),
    .B1(_12234_));
 sg13g2_nand2_1 _19166_ (.Y(_12236_),
    .A(net856),
    .B(_12224_));
 sg13g2_o21ai_1 _19167_ (.B1(_12236_),
    .Y(_00427_),
    .A1(net50),
    .A2(_12235_));
 sg13g2_nor2b_1 _19168_ (.A(_12227_),
    .B_N(\cpu.dcache.r_data[3][19] ),
    .Y(_12237_));
 sg13g2_a21oi_1 _19169_ (.A1(net973),
    .A2(_12227_),
    .Y(_12238_),
    .B1(_12237_));
 sg13g2_nand2_1 _19170_ (.Y(_12239_),
    .A(_11985_),
    .B(_12224_));
 sg13g2_o21ai_1 _19171_ (.B1(_12239_),
    .Y(_00428_),
    .A1(net50),
    .A2(_12238_));
 sg13g2_nor2b_1 _19172_ (.A(_12199_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12240_));
 sg13g2_a21oi_1 _19173_ (.A1(net972),
    .A2(_12199_),
    .Y(_12241_),
    .B1(_12240_));
 sg13g2_nand2_1 _19174_ (.Y(_12242_),
    .A(net857),
    .B(net52));
 sg13g2_o21ai_1 _19175_ (.B1(_12242_),
    .Y(_00429_),
    .A1(net52),
    .A2(_12241_));
 sg13g2_nor2_1 _19176_ (.A(_12193_),
    .B(_11862_),
    .Y(_12243_));
 sg13g2_buf_2 _19177_ (.A(_12243_),
    .X(_12244_));
 sg13g2_nor2b_1 _19178_ (.A(_12244_),
    .B_N(\cpu.dcache.r_data[3][20] ),
    .Y(_12245_));
 sg13g2_a21oi_1 _19179_ (.A1(net975),
    .A2(_12244_),
    .Y(_12246_),
    .B1(_12245_));
 sg13g2_nand2_1 _19180_ (.Y(_12247_),
    .A(net971),
    .B(_12224_));
 sg13g2_o21ai_1 _19181_ (.B1(_12247_),
    .Y(_00430_),
    .A1(net50),
    .A2(_12246_));
 sg13g2_nor2b_1 _19182_ (.A(_12244_),
    .B_N(\cpu.dcache.r_data[3][21] ),
    .Y(_12248_));
 sg13g2_a21oi_1 _19183_ (.A1(net972),
    .A2(_12244_),
    .Y(_12249_),
    .B1(_12248_));
 sg13g2_nand2_1 _19184_ (.Y(_12250_),
    .A(net970),
    .B(_12224_));
 sg13g2_o21ai_1 _19185_ (.B1(_12250_),
    .Y(_00431_),
    .A1(_12225_),
    .A2(_12249_));
 sg13g2_nor2b_1 _19186_ (.A(_12244_),
    .B_N(\cpu.dcache.r_data[3][22] ),
    .Y(_12251_));
 sg13g2_a21oi_1 _19187_ (.A1(net974),
    .A2(_12244_),
    .Y(_12252_),
    .B1(_12251_));
 sg13g2_nand2_1 _19188_ (.Y(_12253_),
    .A(net969),
    .B(_12224_));
 sg13g2_o21ai_1 _19189_ (.B1(_12253_),
    .Y(_00432_),
    .A1(_12225_),
    .A2(_12252_));
 sg13g2_nor2b_1 _19190_ (.A(_12244_),
    .B_N(\cpu.dcache.r_data[3][23] ),
    .Y(_12254_));
 sg13g2_a21oi_1 _19191_ (.A1(net973),
    .A2(_12244_),
    .Y(_12255_),
    .B1(_12254_));
 sg13g2_nand2_1 _19192_ (.Y(_12256_),
    .A(net976),
    .B(_12224_));
 sg13g2_o21ai_1 _19193_ (.B1(_12256_),
    .Y(_00433_),
    .A1(net50),
    .A2(_12255_));
 sg13g2_nor2_1 _19194_ (.A(_12194_),
    .B(_12009_),
    .Y(_12257_));
 sg13g2_buf_1 _19195_ (.A(_12257_),
    .X(_12258_));
 sg13g2_buf_1 _19196_ (.A(_12258_),
    .X(_12259_));
 sg13g2_nor2_1 _19197_ (.A(_12193_),
    .B(_12015_),
    .Y(_12260_));
 sg13g2_buf_1 _19198_ (.A(_12260_),
    .X(_12261_));
 sg13g2_nor2b_1 _19199_ (.A(net419),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12262_));
 sg13g2_a21oi_1 _19200_ (.A1(_12072_),
    .A2(net419),
    .Y(_12263_),
    .B1(_12262_));
 sg13g2_nand2_1 _19201_ (.Y(_12264_),
    .A(net485),
    .B(net49));
 sg13g2_o21ai_1 _19202_ (.B1(_12264_),
    .Y(_00434_),
    .A1(net49),
    .A2(_12263_));
 sg13g2_nor2b_1 _19203_ (.A(net419),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12265_));
 sg13g2_a21oi_1 _19204_ (.A1(_12108_),
    .A2(net419),
    .Y(_12266_),
    .B1(_12265_));
 sg13g2_nand2_1 _19205_ (.Y(_12267_),
    .A(net484),
    .B(net49));
 sg13g2_o21ai_1 _19206_ (.B1(_12267_),
    .Y(_00435_),
    .A1(net49),
    .A2(_12266_));
 sg13g2_nor2b_1 _19207_ (.A(net419),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12268_));
 sg13g2_a21oi_1 _19208_ (.A1(_12081_),
    .A2(net419),
    .Y(_12269_),
    .B1(_12268_));
 sg13g2_nand2_1 _19209_ (.Y(_12270_),
    .A(_11806_),
    .B(_12258_));
 sg13g2_o21ai_1 _19210_ (.B1(_12270_),
    .Y(_00436_),
    .A1(net49),
    .A2(_12269_));
 sg13g2_nor2b_1 _19211_ (.A(net419),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12271_));
 sg13g2_a21oi_1 _19212_ (.A1(_12087_),
    .A2(net419),
    .Y(_12272_),
    .B1(_12271_));
 sg13g2_nand2_1 _19213_ (.Y(_12273_),
    .A(_11816_),
    .B(_12258_));
 sg13g2_o21ai_1 _19214_ (.B1(_12273_),
    .Y(_00437_),
    .A1(net49),
    .A2(_12272_));
 sg13g2_nor2_2 _19215_ (.A(_12194_),
    .B(_11890_),
    .Y(_12274_));
 sg13g2_mux2_1 _19216_ (.A0(\cpu.dcache.r_data[3][28] ),
    .A1(_11949_),
    .S(_12274_),
    .X(_12275_));
 sg13g2_nor2_1 _19217_ (.A(_12258_),
    .B(_12275_),
    .Y(_12276_));
 sg13g2_a21oi_1 _19218_ (.A1(_11888_),
    .A2(_12259_),
    .Y(_00438_),
    .B1(_12276_));
 sg13g2_mux2_1 _19219_ (.A0(\cpu.dcache.r_data[3][29] ),
    .A1(net1072),
    .S(_12274_),
    .X(_12277_));
 sg13g2_nor2_1 _19220_ (.A(_12258_),
    .B(_12277_),
    .Y(_12278_));
 sg13g2_a21oi_1 _19221_ (.A1(net422),
    .A2(net49),
    .Y(_00439_),
    .B1(_12278_));
 sg13g2_buf_1 _19222_ (.A(net1075),
    .X(_12279_));
 sg13g2_nor2b_1 _19223_ (.A(_12199_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12280_));
 sg13g2_a21oi_1 _19224_ (.A1(net968),
    .A2(_12199_),
    .Y(_12281_),
    .B1(_12280_));
 sg13g2_nand2_1 _19225_ (.Y(_12282_),
    .A(net856),
    .B(_12196_));
 sg13g2_o21ai_1 _19226_ (.B1(_12282_),
    .Y(_00440_),
    .A1(net52),
    .A2(_12281_));
 sg13g2_mux2_1 _19227_ (.A0(\cpu.dcache.r_data[3][30] ),
    .A1(net1071),
    .S(_12274_),
    .X(_12283_));
 sg13g2_nor2_1 _19228_ (.A(_12258_),
    .B(_12283_),
    .Y(_12284_));
 sg13g2_a21oi_1 _19229_ (.A1(net421),
    .A2(net49),
    .Y(_00441_),
    .B1(_12284_));
 sg13g2_mux2_1 _19230_ (.A0(\cpu.dcache.r_data[3][31] ),
    .A1(_11959_),
    .S(_12274_),
    .X(_12285_));
 sg13g2_nor2_1 _19231_ (.A(_12258_),
    .B(_12285_),
    .Y(_12286_));
 sg13g2_a21oi_1 _19232_ (.A1(net420),
    .A2(_12259_),
    .Y(_00442_),
    .B1(_12286_));
 sg13g2_buf_1 _19233_ (.A(net1074),
    .X(_12287_));
 sg13g2_nor2b_1 _19234_ (.A(_12199_),
    .B_N(\cpu.dcache.r_data[3][3] ),
    .Y(_12288_));
 sg13g2_a21oi_1 _19235_ (.A1(net967),
    .A2(_12199_),
    .Y(_12289_),
    .B1(_12288_));
 sg13g2_nand2_1 _19236_ (.Y(_12290_),
    .A(_11985_),
    .B(_12196_));
 sg13g2_o21ai_1 _19237_ (.B1(_12290_),
    .Y(_00443_),
    .A1(net52),
    .A2(_12289_));
 sg13g2_buf_1 _19238_ (.A(net1076),
    .X(_12291_));
 sg13g2_nor2_1 _19239_ (.A(_12193_),
    .B(_11907_),
    .Y(_12292_));
 sg13g2_buf_2 _19240_ (.A(_12292_),
    .X(_12293_));
 sg13g2_nor2b_1 _19241_ (.A(_12293_),
    .B_N(\cpu.dcache.r_data[3][4] ),
    .Y(_12294_));
 sg13g2_a21oi_1 _19242_ (.A1(net966),
    .A2(_12293_),
    .Y(_12295_),
    .B1(_12294_));
 sg13g2_nand2_1 _19243_ (.Y(_12296_),
    .A(net971),
    .B(_12196_));
 sg13g2_o21ai_1 _19244_ (.B1(_12296_),
    .Y(_00444_),
    .A1(net52),
    .A2(_12295_));
 sg13g2_buf_1 _19245_ (.A(net1069),
    .X(_12297_));
 sg13g2_nor2b_1 _19246_ (.A(_12293_),
    .B_N(\cpu.dcache.r_data[3][5] ),
    .Y(_12298_));
 sg13g2_a21oi_1 _19247_ (.A1(net965),
    .A2(_12293_),
    .Y(_12299_),
    .B1(_12298_));
 sg13g2_nand2_1 _19248_ (.Y(_12300_),
    .A(net970),
    .B(_12196_));
 sg13g2_o21ai_1 _19249_ (.B1(_12300_),
    .Y(_00445_),
    .A1(net52),
    .A2(_12299_));
 sg13g2_nor2b_1 _19250_ (.A(_12293_),
    .B_N(\cpu.dcache.r_data[3][6] ),
    .Y(_12301_));
 sg13g2_a21oi_1 _19251_ (.A1(net968),
    .A2(_12293_),
    .Y(_12302_),
    .B1(_12301_));
 sg13g2_nand2_1 _19252_ (.Y(_12303_),
    .A(net969),
    .B(_12196_));
 sg13g2_o21ai_1 _19253_ (.B1(_12303_),
    .Y(_00446_),
    .A1(net52),
    .A2(_12302_));
 sg13g2_nor2b_1 _19254_ (.A(_12293_),
    .B_N(\cpu.dcache.r_data[3][7] ),
    .Y(_12304_));
 sg13g2_a21oi_1 _19255_ (.A1(net967),
    .A2(_12293_),
    .Y(_12305_),
    .B1(_12304_));
 sg13g2_nand2_1 _19256_ (.Y(_12306_),
    .A(net976),
    .B(_12196_));
 sg13g2_o21ai_1 _19257_ (.B1(_12306_),
    .Y(_00447_),
    .A1(_12197_),
    .A2(_12305_));
 sg13g2_nor2b_1 _19258_ (.A(_12207_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12307_));
 sg13g2_a21oi_1 _19259_ (.A1(net966),
    .A2(_12207_),
    .Y(_12308_),
    .B1(_12307_));
 sg13g2_nand2_1 _19260_ (.Y(_12309_),
    .A(net485),
    .B(_12204_));
 sg13g2_o21ai_1 _19261_ (.B1(_12309_),
    .Y(_00448_),
    .A1(net51),
    .A2(_12308_));
 sg13g2_nor2b_1 _19262_ (.A(_12207_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12310_));
 sg13g2_a21oi_1 _19263_ (.A1(_12297_),
    .A2(_12207_),
    .Y(_12311_),
    .B1(_12310_));
 sg13g2_nand2_1 _19264_ (.Y(_12312_),
    .A(net484),
    .B(_12204_));
 sg13g2_o21ai_1 _19265_ (.B1(_12312_),
    .Y(_00449_),
    .A1(net51),
    .A2(_12311_));
 sg13g2_buf_1 _19266_ (.A(_09947_),
    .X(_12313_));
 sg13g2_nor2_1 _19267_ (.A(net599),
    .B(_11920_),
    .Y(_12314_));
 sg13g2_buf_2 _19268_ (.A(_12314_),
    .X(_12315_));
 sg13g2_buf_1 _19269_ (.A(_12315_),
    .X(_12316_));
 sg13g2_nor2_1 _19270_ (.A(net599),
    .B(_11774_),
    .Y(_12317_));
 sg13g2_buf_2 _19271_ (.A(_12317_),
    .X(_12318_));
 sg13g2_nor2b_1 _19272_ (.A(_12318_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12319_));
 sg13g2_a21oi_1 _19273_ (.A1(net966),
    .A2(_12318_),
    .Y(_12320_),
    .B1(_12319_));
 sg13g2_nand2_1 _19274_ (.Y(_12321_),
    .A(net860),
    .B(net48));
 sg13g2_o21ai_1 _19275_ (.B1(_12321_),
    .Y(_00450_),
    .A1(net48),
    .A2(_12320_));
 sg13g2_nor2_1 _19276_ (.A(net599),
    .B(_11933_),
    .Y(_12322_));
 sg13g2_buf_1 _19277_ (.A(_12322_),
    .X(_12323_));
 sg13g2_buf_1 _19278_ (.A(_12323_),
    .X(_12324_));
 sg13g2_nor2_1 _19279_ (.A(_12313_),
    .B(_11797_),
    .Y(_12325_));
 sg13g2_buf_2 _19280_ (.A(_12325_),
    .X(_12326_));
 sg13g2_nor2b_1 _19281_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12327_));
 sg13g2_a21oi_1 _19282_ (.A1(net968),
    .A2(_12326_),
    .Y(_12328_),
    .B1(_12327_));
 sg13g2_nand2_1 _19283_ (.Y(_12329_),
    .A(net487),
    .B(net47));
 sg13g2_o21ai_1 _19284_ (.B1(_12329_),
    .Y(_00451_),
    .A1(net47),
    .A2(_12328_));
 sg13g2_nor2b_1 _19285_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12330_));
 sg13g2_a21oi_1 _19286_ (.A1(net967),
    .A2(_12326_),
    .Y(_12331_),
    .B1(_12330_));
 sg13g2_nand2_1 _19287_ (.Y(_12332_),
    .A(net486),
    .B(net47));
 sg13g2_o21ai_1 _19288_ (.B1(_12332_),
    .Y(_00452_),
    .A1(net47),
    .A2(_12331_));
 sg13g2_nor2_2 _19289_ (.A(net599),
    .B(_11823_),
    .Y(_12333_));
 sg13g2_mux2_1 _19290_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(net1073),
    .S(_12333_),
    .X(_12334_));
 sg13g2_nor2_1 _19291_ (.A(_12323_),
    .B(_12334_),
    .Y(_12335_));
 sg13g2_a21oi_1 _19292_ (.A1(net423),
    .A2(_12324_),
    .Y(_00453_),
    .B1(_12335_));
 sg13g2_mux2_1 _19293_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(net1072),
    .S(_12333_),
    .X(_12336_));
 sg13g2_nor2_1 _19294_ (.A(_12323_),
    .B(_12336_),
    .Y(_12337_));
 sg13g2_a21oi_1 _19295_ (.A1(net422),
    .A2(net47),
    .Y(_00454_),
    .B1(_12337_));
 sg13g2_mux2_1 _19296_ (.A0(\cpu.dcache.r_data[4][14] ),
    .A1(net1071),
    .S(_12333_),
    .X(_12338_));
 sg13g2_nor2_1 _19297_ (.A(_12323_),
    .B(_12338_),
    .Y(_12339_));
 sg13g2_a21oi_1 _19298_ (.A1(_11899_),
    .A2(net47),
    .Y(_00455_),
    .B1(_12339_));
 sg13g2_mux2_1 _19299_ (.A0(\cpu.dcache.r_data[4][15] ),
    .A1(net1070),
    .S(_12333_),
    .X(_12340_));
 sg13g2_nor2_1 _19300_ (.A(_12323_),
    .B(_12340_),
    .Y(_12341_));
 sg13g2_a21oi_1 _19301_ (.A1(net420),
    .A2(_12324_),
    .Y(_00456_),
    .B1(_12341_));
 sg13g2_nor2_1 _19302_ (.A(net599),
    .B(_11963_),
    .Y(_12342_));
 sg13g2_buf_2 _19303_ (.A(_12342_),
    .X(_12343_));
 sg13g2_buf_1 _19304_ (.A(_12343_),
    .X(_12344_));
 sg13g2_nor2_1 _19305_ (.A(net599),
    .B(_11846_),
    .Y(_12345_));
 sg13g2_buf_2 _19306_ (.A(_12345_),
    .X(_12346_));
 sg13g2_nor2b_1 _19307_ (.A(_12346_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12347_));
 sg13g2_a21oi_1 _19308_ (.A1(net966),
    .A2(_12346_),
    .Y(_12348_),
    .B1(_12347_));
 sg13g2_nand2_1 _19309_ (.Y(_12349_),
    .A(net860),
    .B(net46));
 sg13g2_o21ai_1 _19310_ (.B1(_12349_),
    .Y(_00457_),
    .A1(net46),
    .A2(_12348_));
 sg13g2_nor2b_1 _19311_ (.A(_12346_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12350_));
 sg13g2_a21oi_1 _19312_ (.A1(net965),
    .A2(_12346_),
    .Y(_12351_),
    .B1(_12350_));
 sg13g2_nand2_1 _19313_ (.Y(_12352_),
    .A(_12120_),
    .B(_12344_));
 sg13g2_o21ai_1 _19314_ (.B1(_12352_),
    .Y(_00458_),
    .A1(_12344_),
    .A2(_12351_));
 sg13g2_nor2b_1 _19315_ (.A(_12346_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12353_));
 sg13g2_a21oi_1 _19316_ (.A1(_12279_),
    .A2(_12346_),
    .Y(_12354_),
    .B1(_12353_));
 sg13g2_nand2_1 _19317_ (.Y(_12355_),
    .A(_12160_),
    .B(_12343_));
 sg13g2_o21ai_1 _19318_ (.B1(_12355_),
    .Y(_00459_),
    .A1(net46),
    .A2(_12354_));
 sg13g2_nor2b_1 _19319_ (.A(_12346_),
    .B_N(\cpu.dcache.r_data[4][19] ),
    .Y(_12356_));
 sg13g2_a21oi_1 _19320_ (.A1(_12287_),
    .A2(_12346_),
    .Y(_12357_),
    .B1(_12356_));
 sg13g2_buf_1 _19321_ (.A(net1098),
    .X(_12358_));
 sg13g2_nand2_1 _19322_ (.Y(_12359_),
    .A(net964),
    .B(_12343_));
 sg13g2_o21ai_1 _19323_ (.B1(_12359_),
    .Y(_00460_),
    .A1(net46),
    .A2(_12357_));
 sg13g2_inv_1 _19324_ (.Y(_12360_),
    .A(\cpu.dcache.r_data[4][1] ));
 sg13g2_nor2_1 _19325_ (.A(_12360_),
    .B(_12318_),
    .Y(_12361_));
 sg13g2_a21oi_1 _19326_ (.A1(net965),
    .A2(_12318_),
    .Y(_12362_),
    .B1(_12361_));
 sg13g2_nand2_1 _19327_ (.Y(_12363_),
    .A(net857),
    .B(net48));
 sg13g2_o21ai_1 _19328_ (.B1(_12363_),
    .Y(_00461_),
    .A1(net48),
    .A2(_12362_));
 sg13g2_nor2_1 _19329_ (.A(_09947_),
    .B(_11862_),
    .Y(_12364_));
 sg13g2_buf_2 _19330_ (.A(_12364_),
    .X(_12365_));
 sg13g2_nor2b_1 _19331_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12366_));
 sg13g2_a21oi_1 _19332_ (.A1(net966),
    .A2(_12365_),
    .Y(_12367_),
    .B1(_12366_));
 sg13g2_nand2_1 _19333_ (.Y(_12368_),
    .A(_12173_),
    .B(_12343_));
 sg13g2_o21ai_1 _19334_ (.B1(_12368_),
    .Y(_00462_),
    .A1(net46),
    .A2(_12367_));
 sg13g2_nor2b_1 _19335_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12369_));
 sg13g2_a21oi_1 _19336_ (.A1(net965),
    .A2(_12365_),
    .Y(_12370_),
    .B1(_12369_));
 sg13g2_nand2_1 _19337_ (.Y(_12371_),
    .A(net970),
    .B(_12343_));
 sg13g2_o21ai_1 _19338_ (.B1(_12371_),
    .Y(_00463_),
    .A1(net46),
    .A2(_12370_));
 sg13g2_nor2b_1 _19339_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[4][22] ),
    .Y(_12372_));
 sg13g2_a21oi_1 _19340_ (.A1(_12279_),
    .A2(_12365_),
    .Y(_12373_),
    .B1(_12372_));
 sg13g2_nand2_1 _19341_ (.Y(_12374_),
    .A(net969),
    .B(_12343_));
 sg13g2_o21ai_1 _19342_ (.B1(_12374_),
    .Y(_00464_),
    .A1(net46),
    .A2(_12373_));
 sg13g2_nor2b_1 _19343_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[4][23] ),
    .Y(_12375_));
 sg13g2_a21oi_1 _19344_ (.A1(_12287_),
    .A2(_12365_),
    .Y(_12376_),
    .B1(_12375_));
 sg13g2_nand2_1 _19345_ (.Y(_12377_),
    .A(net976),
    .B(_12343_));
 sg13g2_o21ai_1 _19346_ (.B1(_12377_),
    .Y(_00465_),
    .A1(net46),
    .A2(_12376_));
 sg13g2_buf_1 _19347_ (.A(_09394_),
    .X(_12378_));
 sg13g2_nand2_1 _19348_ (.Y(_12379_),
    .A(_12378_),
    .B(_11782_));
 sg13g2_buf_2 _19349_ (.A(_12379_),
    .X(_12380_));
 sg13g2_mux2_1 _19350_ (.A0(_11761_),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(_12380_),
    .X(_12381_));
 sg13g2_nor2_1 _19351_ (.A(net599),
    .B(_12009_),
    .Y(_12382_));
 sg13g2_buf_1 _19352_ (.A(_12382_),
    .X(_12383_));
 sg13g2_mux2_1 _19353_ (.A0(_12381_),
    .A1(_11877_),
    .S(net63),
    .X(_00466_));
 sg13g2_mux2_1 _19354_ (.A0(_11832_),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(_12380_),
    .X(_12384_));
 sg13g2_mux2_1 _19355_ (.A0(_12384_),
    .A1(_11885_),
    .S(net63),
    .X(_00467_));
 sg13g2_mux2_1 _19356_ (.A0(net1079),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(_12380_),
    .X(_12385_));
 sg13g2_mux2_1 _19357_ (.A0(_12385_),
    .A1(net487),
    .S(net63),
    .X(_00468_));
 sg13g2_mux2_1 _19358_ (.A0(net1078),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(_12380_),
    .X(_12386_));
 sg13g2_mux2_1 _19359_ (.A0(_12386_),
    .A1(net486),
    .S(net63),
    .X(_00469_));
 sg13g2_nor2_2 _19360_ (.A(_12313_),
    .B(_11890_),
    .Y(_12387_));
 sg13g2_mux2_1 _19361_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(net1073),
    .S(_12387_),
    .X(_12388_));
 sg13g2_nor2_1 _19362_ (.A(net63),
    .B(_12388_),
    .Y(_12389_));
 sg13g2_a21oi_1 _19363_ (.A1(_11888_),
    .A2(net63),
    .Y(_00470_),
    .B1(_12389_));
 sg13g2_mux2_1 _19364_ (.A0(\cpu.dcache.r_data[4][29] ),
    .A1(net1072),
    .S(_12387_),
    .X(_12390_));
 sg13g2_nor2_1 _19365_ (.A(_12383_),
    .B(_12390_),
    .Y(_12391_));
 sg13g2_a21oi_1 _19366_ (.A1(_11895_),
    .A2(_12383_),
    .Y(_00471_),
    .B1(_12391_));
 sg13g2_nor2b_1 _19367_ (.A(_12318_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12392_));
 sg13g2_a21oi_1 _19368_ (.A1(net968),
    .A2(_12318_),
    .Y(_12393_),
    .B1(_12392_));
 sg13g2_nand2_1 _19369_ (.Y(_12394_),
    .A(net856),
    .B(_12315_));
 sg13g2_o21ai_1 _19370_ (.B1(_12394_),
    .Y(_00472_),
    .A1(_12316_),
    .A2(_12393_));
 sg13g2_mux2_1 _19371_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(_11956_),
    .S(_12387_),
    .X(_12395_));
 sg13g2_nor2_1 _19372_ (.A(_12382_),
    .B(_12395_),
    .Y(_12396_));
 sg13g2_a21oi_1 _19373_ (.A1(net421),
    .A2(net63),
    .Y(_00473_),
    .B1(_12396_));
 sg13g2_mux2_1 _19374_ (.A0(\cpu.dcache.r_data[4][31] ),
    .A1(net1070),
    .S(_12387_),
    .X(_12397_));
 sg13g2_nor2_1 _19375_ (.A(_12382_),
    .B(_12397_),
    .Y(_12398_));
 sg13g2_a21oi_1 _19376_ (.A1(net420),
    .A2(net63),
    .Y(_00474_),
    .B1(_12398_));
 sg13g2_nor2b_1 _19377_ (.A(_12318_),
    .B_N(\cpu.dcache.r_data[4][3] ),
    .Y(_12399_));
 sg13g2_a21oi_1 _19378_ (.A1(net967),
    .A2(_12318_),
    .Y(_12400_),
    .B1(_12399_));
 sg13g2_nand2_1 _19379_ (.Y(_12401_),
    .A(net964),
    .B(_12315_));
 sg13g2_o21ai_1 _19380_ (.B1(_12401_),
    .Y(_00475_),
    .A1(_12316_),
    .A2(_12400_));
 sg13g2_nor2_1 _19381_ (.A(_09947_),
    .B(_11907_),
    .Y(_12402_));
 sg13g2_buf_2 _19382_ (.A(_12402_),
    .X(_12403_));
 sg13g2_nor2b_1 _19383_ (.A(_12403_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_12404_));
 sg13g2_a21oi_1 _19384_ (.A1(net966),
    .A2(_12403_),
    .Y(_12405_),
    .B1(_12404_));
 sg13g2_nand2_1 _19385_ (.Y(_12406_),
    .A(net971),
    .B(_12315_));
 sg13g2_o21ai_1 _19386_ (.B1(_12406_),
    .Y(_00476_),
    .A1(net48),
    .A2(_12405_));
 sg13g2_nor2b_1 _19387_ (.A(_12403_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_12407_));
 sg13g2_a21oi_1 _19388_ (.A1(net965),
    .A2(_12403_),
    .Y(_12408_),
    .B1(_12407_));
 sg13g2_nand2_1 _19389_ (.Y(_12409_),
    .A(net970),
    .B(_12315_));
 sg13g2_o21ai_1 _19390_ (.B1(_12409_),
    .Y(_00477_),
    .A1(net48),
    .A2(_12408_));
 sg13g2_nor2b_1 _19391_ (.A(_12403_),
    .B_N(\cpu.dcache.r_data[4][6] ),
    .Y(_12410_));
 sg13g2_a21oi_1 _19392_ (.A1(net968),
    .A2(_12403_),
    .Y(_12411_),
    .B1(_12410_));
 sg13g2_nand2_1 _19393_ (.Y(_12412_),
    .A(net969),
    .B(_12315_));
 sg13g2_o21ai_1 _19394_ (.B1(_12412_),
    .Y(_00478_),
    .A1(net48),
    .A2(_12411_));
 sg13g2_nor2b_1 _19395_ (.A(_12403_),
    .B_N(\cpu.dcache.r_data[4][7] ),
    .Y(_12413_));
 sg13g2_a21oi_1 _19396_ (.A1(net967),
    .A2(_12403_),
    .Y(_12414_),
    .B1(_12413_));
 sg13g2_nand2_1 _19397_ (.Y(_12415_),
    .A(net976),
    .B(_12315_));
 sg13g2_o21ai_1 _19398_ (.B1(_12415_),
    .Y(_00479_),
    .A1(net48),
    .A2(_12414_));
 sg13g2_nor2b_1 _19399_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_12416_));
 sg13g2_a21oi_1 _19400_ (.A1(net966),
    .A2(_12326_),
    .Y(_12417_),
    .B1(_12416_));
 sg13g2_nand2_1 _19401_ (.Y(_12418_),
    .A(net485),
    .B(_12323_));
 sg13g2_o21ai_1 _19402_ (.B1(_12418_),
    .Y(_00480_),
    .A1(net47),
    .A2(_12417_));
 sg13g2_nor2b_1 _19403_ (.A(_12326_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_12419_));
 sg13g2_a21oi_1 _19404_ (.A1(_12297_),
    .A2(_12326_),
    .Y(_12420_),
    .B1(_12419_));
 sg13g2_nand2_1 _19405_ (.Y(_12421_),
    .A(net484),
    .B(_12323_));
 sg13g2_o21ai_1 _19406_ (.B1(_12421_),
    .Y(_00481_),
    .A1(net47),
    .A2(_12420_));
 sg13g2_nand2_1 _19407_ (.Y(_12422_),
    .A(net772),
    .B(net773));
 sg13g2_buf_1 _19408_ (.A(_12422_),
    .X(_12423_));
 sg13g2_buf_1 _19409_ (.A(_12423_),
    .X(_12424_));
 sg13g2_nor2_1 _19410_ (.A(net534),
    .B(_11920_),
    .Y(_12425_));
 sg13g2_buf_2 _19411_ (.A(_12425_),
    .X(_12426_));
 sg13g2_buf_1 _19412_ (.A(_12426_),
    .X(_12427_));
 sg13g2_nor2_1 _19413_ (.A(net534),
    .B(_11774_),
    .Y(_12428_));
 sg13g2_buf_2 _19414_ (.A(_12428_),
    .X(_12429_));
 sg13g2_nor2b_1 _19415_ (.A(_12429_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_12430_));
 sg13g2_a21oi_1 _19416_ (.A1(net966),
    .A2(_12429_),
    .Y(_12431_),
    .B1(_12430_));
 sg13g2_nand2_1 _19417_ (.Y(_12432_),
    .A(net860),
    .B(net45));
 sg13g2_o21ai_1 _19418_ (.B1(_12432_),
    .Y(_00482_),
    .A1(net45),
    .A2(_12431_));
 sg13g2_nor2_1 _19419_ (.A(net534),
    .B(_11933_),
    .Y(_12433_));
 sg13g2_buf_1 _19420_ (.A(_12433_),
    .X(_12434_));
 sg13g2_buf_1 _19421_ (.A(_12434_),
    .X(_12435_));
 sg13g2_nor2_1 _19422_ (.A(_12424_),
    .B(_11797_),
    .Y(_12436_));
 sg13g2_buf_2 _19423_ (.A(_12436_),
    .X(_12437_));
 sg13g2_nor2b_1 _19424_ (.A(_12437_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_12438_));
 sg13g2_a21oi_1 _19425_ (.A1(net968),
    .A2(_12437_),
    .Y(_12439_),
    .B1(_12438_));
 sg13g2_nand2_1 _19426_ (.Y(_12440_),
    .A(_11805_),
    .B(net44));
 sg13g2_o21ai_1 _19427_ (.B1(_12440_),
    .Y(_00483_),
    .A1(net44),
    .A2(_12439_));
 sg13g2_nor2b_1 _19428_ (.A(_12437_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_12441_));
 sg13g2_a21oi_1 _19429_ (.A1(net967),
    .A2(_12437_),
    .Y(_12442_),
    .B1(_12441_));
 sg13g2_nand2_1 _19430_ (.Y(_12443_),
    .A(_11815_),
    .B(net44));
 sg13g2_o21ai_1 _19431_ (.B1(_12443_),
    .Y(_00484_),
    .A1(net44),
    .A2(_12442_));
 sg13g2_nor2_2 _19432_ (.A(net534),
    .B(_11823_),
    .Y(_12444_));
 sg13g2_mux2_1 _19433_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(net1073),
    .S(_12444_),
    .X(_12445_));
 sg13g2_nor2_1 _19434_ (.A(_12434_),
    .B(_12445_),
    .Y(_12446_));
 sg13g2_a21oi_1 _19435_ (.A1(net423),
    .A2(net44),
    .Y(_00485_),
    .B1(_12446_));
 sg13g2_mux2_1 _19436_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(net1072),
    .S(_12444_),
    .X(_12447_));
 sg13g2_nor2_1 _19437_ (.A(_12434_),
    .B(_12447_),
    .Y(_12448_));
 sg13g2_a21oi_1 _19438_ (.A1(net422),
    .A2(net44),
    .Y(_00486_),
    .B1(_12448_));
 sg13g2_mux2_1 _19439_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(net1071),
    .S(_12444_),
    .X(_12449_));
 sg13g2_nor2_1 _19440_ (.A(_12434_),
    .B(_12449_),
    .Y(_12450_));
 sg13g2_a21oi_1 _19441_ (.A1(_11899_),
    .A2(_12435_),
    .Y(_00487_),
    .B1(_12450_));
 sg13g2_mux2_1 _19442_ (.A0(\cpu.dcache.r_data[5][15] ),
    .A1(net1070),
    .S(_12444_),
    .X(_12451_));
 sg13g2_nor2_1 _19443_ (.A(_12434_),
    .B(_12451_),
    .Y(_12452_));
 sg13g2_a21oi_1 _19444_ (.A1(net420),
    .A2(_12435_),
    .Y(_00488_),
    .B1(_12452_));
 sg13g2_nor2_1 _19445_ (.A(net534),
    .B(_11963_),
    .Y(_12453_));
 sg13g2_buf_2 _19446_ (.A(_12453_),
    .X(_12454_));
 sg13g2_buf_1 _19447_ (.A(_12454_),
    .X(_12455_));
 sg13g2_nor2_1 _19448_ (.A(net534),
    .B(_11846_),
    .Y(_12456_));
 sg13g2_buf_2 _19449_ (.A(_12456_),
    .X(_12457_));
 sg13g2_nor2b_1 _19450_ (.A(_12457_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_12458_));
 sg13g2_a21oi_1 _19451_ (.A1(_12291_),
    .A2(_12457_),
    .Y(_12459_),
    .B1(_12458_));
 sg13g2_nand2_1 _19452_ (.Y(_12460_),
    .A(net860),
    .B(net43));
 sg13g2_o21ai_1 _19453_ (.B1(_12460_),
    .Y(_00489_),
    .A1(net43),
    .A2(_12459_));
 sg13g2_nor2b_1 _19454_ (.A(_12457_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_12461_));
 sg13g2_a21oi_1 _19455_ (.A1(net965),
    .A2(_12457_),
    .Y(_12462_),
    .B1(_12461_));
 sg13g2_nand2_1 _19456_ (.Y(_12463_),
    .A(net857),
    .B(net43));
 sg13g2_o21ai_1 _19457_ (.B1(_12463_),
    .Y(_00490_),
    .A1(net43),
    .A2(_12462_));
 sg13g2_nor2b_1 _19458_ (.A(_12457_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12464_));
 sg13g2_a21oi_1 _19459_ (.A1(net968),
    .A2(_12457_),
    .Y(_12465_),
    .B1(_12464_));
 sg13g2_nand2_1 _19460_ (.Y(_12466_),
    .A(net856),
    .B(_12454_));
 sg13g2_o21ai_1 _19461_ (.B1(_12466_),
    .Y(_00491_),
    .A1(net43),
    .A2(_12465_));
 sg13g2_nor2b_1 _19462_ (.A(_12457_),
    .B_N(\cpu.dcache.r_data[5][19] ),
    .Y(_12467_));
 sg13g2_a21oi_1 _19463_ (.A1(net967),
    .A2(_12457_),
    .Y(_12468_),
    .B1(_12467_));
 sg13g2_nand2_1 _19464_ (.Y(_12469_),
    .A(_12358_),
    .B(_12454_));
 sg13g2_o21ai_1 _19465_ (.B1(_12469_),
    .Y(_00492_),
    .A1(net43),
    .A2(_12468_));
 sg13g2_nor2b_1 _19466_ (.A(_12429_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_12470_));
 sg13g2_a21oi_1 _19467_ (.A1(net965),
    .A2(_12429_),
    .Y(_12471_),
    .B1(_12470_));
 sg13g2_nand2_1 _19468_ (.Y(_12472_),
    .A(_12120_),
    .B(_12427_));
 sg13g2_o21ai_1 _19469_ (.B1(_12472_),
    .Y(_00493_),
    .A1(_12427_),
    .A2(_12471_));
 sg13g2_nor2_1 _19470_ (.A(_12423_),
    .B(_11862_),
    .Y(_12473_));
 sg13g2_buf_2 _19471_ (.A(_12473_),
    .X(_12474_));
 sg13g2_nor2b_1 _19472_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_12475_));
 sg13g2_a21oi_1 _19473_ (.A1(_12291_),
    .A2(_12474_),
    .Y(_12476_),
    .B1(_12475_));
 sg13g2_nand2_1 _19474_ (.Y(_12477_),
    .A(net971),
    .B(_12454_));
 sg13g2_o21ai_1 _19475_ (.B1(_12477_),
    .Y(_00494_),
    .A1(net43),
    .A2(_12476_));
 sg13g2_nor2b_1 _19476_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_12478_));
 sg13g2_a21oi_1 _19477_ (.A1(net965),
    .A2(_12474_),
    .Y(_12479_),
    .B1(_12478_));
 sg13g2_nand2_1 _19478_ (.Y(_12480_),
    .A(net970),
    .B(_12454_));
 sg13g2_o21ai_1 _19479_ (.B1(_12480_),
    .Y(_00495_),
    .A1(_12455_),
    .A2(_12479_));
 sg13g2_nor2b_1 _19480_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[5][22] ),
    .Y(_12481_));
 sg13g2_a21oi_1 _19481_ (.A1(net968),
    .A2(_12474_),
    .Y(_12482_),
    .B1(_12481_));
 sg13g2_nand2_1 _19482_ (.Y(_12483_),
    .A(net969),
    .B(_12454_));
 sg13g2_o21ai_1 _19483_ (.B1(_12483_),
    .Y(_00496_),
    .A1(net43),
    .A2(_12482_));
 sg13g2_nor2b_1 _19484_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[5][23] ),
    .Y(_12484_));
 sg13g2_a21oi_1 _19485_ (.A1(net967),
    .A2(_12474_),
    .Y(_12485_),
    .B1(_12484_));
 sg13g2_nand2_1 _19486_ (.Y(_12486_),
    .A(_12058_),
    .B(_12454_));
 sg13g2_o21ai_1 _19487_ (.B1(_12486_),
    .Y(_00497_),
    .A1(_12455_),
    .A2(_12485_));
 sg13g2_nor2_1 _19488_ (.A(net534),
    .B(_12009_),
    .Y(_12487_));
 sg13g2_buf_1 _19489_ (.A(_12487_),
    .X(_12488_));
 sg13g2_buf_1 _19490_ (.A(_12488_),
    .X(_12489_));
 sg13g2_buf_1 _19491_ (.A(net1076),
    .X(_12490_));
 sg13g2_nor2_1 _19492_ (.A(net597),
    .B(_12015_),
    .Y(_12491_));
 sg13g2_buf_1 _19493_ (.A(_12491_),
    .X(_12492_));
 sg13g2_nor2b_1 _19494_ (.A(net481),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_12493_));
 sg13g2_a21oi_1 _19495_ (.A1(_12490_),
    .A2(_12492_),
    .Y(_12494_),
    .B1(_12493_));
 sg13g2_nand2_1 _19496_ (.Y(_12495_),
    .A(_11876_),
    .B(net42));
 sg13g2_o21ai_1 _19497_ (.B1(_12495_),
    .Y(_00498_),
    .A1(net42),
    .A2(_12494_));
 sg13g2_buf_1 _19498_ (.A(net1069),
    .X(_12496_));
 sg13g2_nor2b_1 _19499_ (.A(net481),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_12497_));
 sg13g2_a21oi_1 _19500_ (.A1(net962),
    .A2(net481),
    .Y(_12498_),
    .B1(_12497_));
 sg13g2_nand2_1 _19501_ (.Y(_12499_),
    .A(_11884_),
    .B(net42));
 sg13g2_o21ai_1 _19502_ (.B1(_12499_),
    .Y(_00499_),
    .A1(_12489_),
    .A2(_12498_));
 sg13g2_buf_1 _19503_ (.A(net1075),
    .X(_12500_));
 sg13g2_nor2b_1 _19504_ (.A(net481),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_12501_));
 sg13g2_a21oi_1 _19505_ (.A1(_12500_),
    .A2(net481),
    .Y(_12502_),
    .B1(_12501_));
 sg13g2_nand2_1 _19506_ (.Y(_12503_),
    .A(_11805_),
    .B(_12488_));
 sg13g2_o21ai_1 _19507_ (.B1(_12503_),
    .Y(_00500_),
    .A1(net42),
    .A2(_12502_));
 sg13g2_buf_1 _19508_ (.A(net1074),
    .X(_12504_));
 sg13g2_nor2b_1 _19509_ (.A(net481),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_12505_));
 sg13g2_a21oi_1 _19510_ (.A1(net960),
    .A2(net481),
    .Y(_12506_),
    .B1(_12505_));
 sg13g2_nand2_1 _19511_ (.Y(_12507_),
    .A(_11815_),
    .B(_12488_));
 sg13g2_o21ai_1 _19512_ (.B1(_12507_),
    .Y(_00501_),
    .A1(net42),
    .A2(_12506_));
 sg13g2_nor2_2 _19513_ (.A(_12424_),
    .B(_11890_),
    .Y(_12508_));
 sg13g2_mux2_1 _19514_ (.A0(\cpu.dcache.r_data[5][28] ),
    .A1(_11949_),
    .S(_12508_),
    .X(_12509_));
 sg13g2_nor2_1 _19515_ (.A(_12488_),
    .B(_12509_),
    .Y(_12510_));
 sg13g2_a21oi_1 _19516_ (.A1(_11820_),
    .A2(net42),
    .Y(_00502_),
    .B1(_12510_));
 sg13g2_mux2_1 _19517_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(net1072),
    .S(_12508_),
    .X(_12511_));
 sg13g2_nor2_1 _19518_ (.A(_12488_),
    .B(_12511_),
    .Y(_12512_));
 sg13g2_a21oi_1 _19519_ (.A1(_11830_),
    .A2(net42),
    .Y(_00503_),
    .B1(_12512_));
 sg13g2_nor2b_1 _19520_ (.A(_12429_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_12513_));
 sg13g2_a21oi_1 _19521_ (.A1(net961),
    .A2(_12429_),
    .Y(_12514_),
    .B1(_12513_));
 sg13g2_nand2_1 _19522_ (.Y(_12515_),
    .A(_12160_),
    .B(_12426_));
 sg13g2_o21ai_1 _19523_ (.B1(_12515_),
    .Y(_00504_),
    .A1(net45),
    .A2(_12514_));
 sg13g2_mux2_1 _19524_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(_11956_),
    .S(_12508_),
    .X(_12516_));
 sg13g2_nor2_1 _19525_ (.A(_12488_),
    .B(_12516_),
    .Y(_12517_));
 sg13g2_a21oi_1 _19526_ (.A1(_11837_),
    .A2(net42),
    .Y(_00505_),
    .B1(_12517_));
 sg13g2_mux2_1 _19527_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(_11959_),
    .S(_12508_),
    .X(_12518_));
 sg13g2_nor2_1 _19528_ (.A(_12488_),
    .B(_12518_),
    .Y(_12519_));
 sg13g2_a21oi_1 _19529_ (.A1(_11842_),
    .A2(_12489_),
    .Y(_00506_),
    .B1(_12519_));
 sg13g2_nor2b_1 _19530_ (.A(_12429_),
    .B_N(\cpu.dcache.r_data[5][3] ),
    .Y(_12520_));
 sg13g2_a21oi_1 _19531_ (.A1(net960),
    .A2(_12429_),
    .Y(_12521_),
    .B1(_12520_));
 sg13g2_nand2_1 _19532_ (.Y(_12522_),
    .A(net964),
    .B(_12426_));
 sg13g2_o21ai_1 _19533_ (.B1(_12522_),
    .Y(_00507_),
    .A1(net45),
    .A2(_12521_));
 sg13g2_nor2_1 _19534_ (.A(net597),
    .B(_11907_),
    .Y(_12523_));
 sg13g2_buf_2 _19535_ (.A(_12523_),
    .X(_12524_));
 sg13g2_nor2b_1 _19536_ (.A(_12524_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_12525_));
 sg13g2_a21oi_1 _19537_ (.A1(net963),
    .A2(_12524_),
    .Y(_12526_),
    .B1(_12525_));
 sg13g2_nand2_1 _19538_ (.Y(_12527_),
    .A(net971),
    .B(_12426_));
 sg13g2_o21ai_1 _19539_ (.B1(_12527_),
    .Y(_00508_),
    .A1(net45),
    .A2(_12526_));
 sg13g2_nor2b_1 _19540_ (.A(_12524_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_12528_));
 sg13g2_a21oi_1 _19541_ (.A1(net962),
    .A2(_12524_),
    .Y(_12529_),
    .B1(_12528_));
 sg13g2_nand2_1 _19542_ (.Y(_12530_),
    .A(_12177_),
    .B(_12426_));
 sg13g2_o21ai_1 _19543_ (.B1(_12530_),
    .Y(_00509_),
    .A1(net45),
    .A2(_12529_));
 sg13g2_nor2b_1 _19544_ (.A(_12524_),
    .B_N(\cpu.dcache.r_data[5][6] ),
    .Y(_12531_));
 sg13g2_a21oi_1 _19545_ (.A1(net961),
    .A2(_12524_),
    .Y(_12532_),
    .B1(_12531_));
 sg13g2_nand2_1 _19546_ (.Y(_12533_),
    .A(_12181_),
    .B(_12426_));
 sg13g2_o21ai_1 _19547_ (.B1(_12533_),
    .Y(_00510_),
    .A1(net45),
    .A2(_12532_));
 sg13g2_nor2b_1 _19548_ (.A(_12524_),
    .B_N(\cpu.dcache.r_data[5][7] ),
    .Y(_12534_));
 sg13g2_a21oi_1 _19549_ (.A1(net960),
    .A2(_12524_),
    .Y(_12535_),
    .B1(_12534_));
 sg13g2_nand2_1 _19550_ (.Y(_12536_),
    .A(net976),
    .B(_12426_));
 sg13g2_o21ai_1 _19551_ (.B1(_12536_),
    .Y(_00511_),
    .A1(net45),
    .A2(_12535_));
 sg13g2_nor2b_1 _19552_ (.A(_12437_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_12537_));
 sg13g2_a21oi_1 _19553_ (.A1(net963),
    .A2(_12437_),
    .Y(_12538_),
    .B1(_12537_));
 sg13g2_nand2_1 _19554_ (.Y(_12539_),
    .A(_11876_),
    .B(_12434_));
 sg13g2_o21ai_1 _19555_ (.B1(_12539_),
    .Y(_00512_),
    .A1(net44),
    .A2(_12538_));
 sg13g2_nor2b_1 _19556_ (.A(_12437_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_12540_));
 sg13g2_a21oi_1 _19557_ (.A1(net962),
    .A2(_12437_),
    .Y(_12541_),
    .B1(_12540_));
 sg13g2_nand2_1 _19558_ (.Y(_12542_),
    .A(_11884_),
    .B(_12434_));
 sg13g2_o21ai_1 _19559_ (.B1(_12542_),
    .Y(_00513_),
    .A1(net44),
    .A2(_12541_));
 sg13g2_nand2_1 _19560_ (.Y(_12543_),
    .A(_09091_),
    .B(_09283_));
 sg13g2_buf_1 _19561_ (.A(_12543_),
    .X(_12544_));
 sg13g2_buf_1 _19562_ (.A(net533),
    .X(_12545_));
 sg13g2_nor2_1 _19563_ (.A(net480),
    .B(_11920_),
    .Y(_12546_));
 sg13g2_buf_1 _19564_ (.A(_12546_),
    .X(_12547_));
 sg13g2_buf_1 _19565_ (.A(_12547_),
    .X(_12548_));
 sg13g2_nor2_1 _19566_ (.A(net480),
    .B(_11774_),
    .Y(_12549_));
 sg13g2_buf_2 _19567_ (.A(_12549_),
    .X(_12550_));
 sg13g2_nor2b_1 _19568_ (.A(_12550_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_12551_));
 sg13g2_a21oi_1 _19569_ (.A1(net963),
    .A2(_12550_),
    .Y(_12552_),
    .B1(_12551_));
 sg13g2_nand2_1 _19570_ (.Y(_12553_),
    .A(_11971_),
    .B(net41));
 sg13g2_o21ai_1 _19571_ (.B1(_12553_),
    .Y(_00514_),
    .A1(net41),
    .A2(_12552_));
 sg13g2_nor2_1 _19572_ (.A(net480),
    .B(_11933_),
    .Y(_12554_));
 sg13g2_buf_2 _19573_ (.A(_12554_),
    .X(_12555_));
 sg13g2_buf_1 _19574_ (.A(_12555_),
    .X(_12556_));
 sg13g2_nor2_1 _19575_ (.A(net533),
    .B(_11797_),
    .Y(_12557_));
 sg13g2_buf_2 _19576_ (.A(_12557_),
    .X(_12558_));
 sg13g2_nor2b_1 _19577_ (.A(_12558_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_12559_));
 sg13g2_a21oi_1 _19578_ (.A1(net961),
    .A2(_12558_),
    .Y(_12560_),
    .B1(_12559_));
 sg13g2_nand2_1 _19579_ (.Y(_12561_),
    .A(_11805_),
    .B(net40));
 sg13g2_o21ai_1 _19580_ (.B1(_12561_),
    .Y(_00515_),
    .A1(net40),
    .A2(_12560_));
 sg13g2_nor2b_1 _19581_ (.A(_12558_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_12562_));
 sg13g2_a21oi_1 _19582_ (.A1(net960),
    .A2(_12558_),
    .Y(_12563_),
    .B1(_12562_));
 sg13g2_nand2_1 _19583_ (.Y(_12564_),
    .A(_11815_),
    .B(net40));
 sg13g2_o21ai_1 _19584_ (.B1(_12564_),
    .Y(_00516_),
    .A1(net40),
    .A2(_12563_));
 sg13g2_nor2_2 _19585_ (.A(net480),
    .B(_11823_),
    .Y(_12565_));
 sg13g2_mux2_1 _19586_ (.A0(\cpu.dcache.r_data[6][12] ),
    .A1(net1076),
    .S(_12565_),
    .X(_12566_));
 sg13g2_nor2_1 _19587_ (.A(_12555_),
    .B(_12566_),
    .Y(_12567_));
 sg13g2_a21oi_1 _19588_ (.A1(_11820_),
    .A2(net40),
    .Y(_00517_),
    .B1(_12567_));
 sg13g2_mux2_1 _19589_ (.A0(\cpu.dcache.r_data[6][13] ),
    .A1(_11973_),
    .S(_12565_),
    .X(_12568_));
 sg13g2_nor2_1 _19590_ (.A(_12555_),
    .B(_12568_),
    .Y(_12569_));
 sg13g2_a21oi_1 _19591_ (.A1(_11830_),
    .A2(_12556_),
    .Y(_00518_),
    .B1(_12569_));
 sg13g2_mux2_1 _19592_ (.A0(\cpu.dcache.r_data[6][14] ),
    .A1(net1075),
    .S(_12565_),
    .X(_12570_));
 sg13g2_nor2_1 _19593_ (.A(_12555_),
    .B(_12570_),
    .Y(_12571_));
 sg13g2_a21oi_1 _19594_ (.A1(_11837_),
    .A2(net40),
    .Y(_00519_),
    .B1(_12571_));
 sg13g2_mux2_1 _19595_ (.A0(\cpu.dcache.r_data[6][15] ),
    .A1(net1074),
    .S(_12565_),
    .X(_12572_));
 sg13g2_nor2_1 _19596_ (.A(_12555_),
    .B(_12572_),
    .Y(_12573_));
 sg13g2_a21oi_1 _19597_ (.A1(_11842_),
    .A2(_12556_),
    .Y(_00520_),
    .B1(_12573_));
 sg13g2_nor2_1 _19598_ (.A(net480),
    .B(_11963_),
    .Y(_12574_));
 sg13g2_buf_2 _19599_ (.A(_12574_),
    .X(_12575_));
 sg13g2_buf_1 _19600_ (.A(_12575_),
    .X(_12576_));
 sg13g2_nor2_1 _19601_ (.A(net533),
    .B(_11846_),
    .Y(_12577_));
 sg13g2_buf_2 _19602_ (.A(_12577_),
    .X(_12578_));
 sg13g2_nor2b_1 _19603_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_12579_));
 sg13g2_a21oi_1 _19604_ (.A1(net963),
    .A2(_12578_),
    .Y(_12580_),
    .B1(_12579_));
 sg13g2_buf_1 _19605_ (.A(_09895_),
    .X(_12581_));
 sg13g2_nand2_1 _19606_ (.Y(_12582_),
    .A(_12581_),
    .B(net39));
 sg13g2_o21ai_1 _19607_ (.B1(_12582_),
    .Y(_00521_),
    .A1(net39),
    .A2(_12580_));
 sg13g2_nor2b_1 _19608_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_12583_));
 sg13g2_a21oi_1 _19609_ (.A1(net962),
    .A2(_12578_),
    .Y(_12584_),
    .B1(_12583_));
 sg13g2_nand2_1 _19610_ (.Y(_12585_),
    .A(net857),
    .B(net39));
 sg13g2_o21ai_1 _19611_ (.B1(_12585_),
    .Y(_00522_),
    .A1(net39),
    .A2(_12584_));
 sg13g2_nor2b_1 _19612_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_12586_));
 sg13g2_a21oi_1 _19613_ (.A1(net961),
    .A2(_12578_),
    .Y(_12587_),
    .B1(_12586_));
 sg13g2_nand2_1 _19614_ (.Y(_12588_),
    .A(net856),
    .B(_12575_));
 sg13g2_o21ai_1 _19615_ (.B1(_12588_),
    .Y(_00523_),
    .A1(net39),
    .A2(_12587_));
 sg13g2_nor2b_1 _19616_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[6][19] ),
    .Y(_02684_));
 sg13g2_a21oi_1 _19617_ (.A1(net960),
    .A2(_12578_),
    .Y(_02685_),
    .B1(_02684_));
 sg13g2_nand2_1 _19618_ (.Y(_02686_),
    .A(net964),
    .B(_12575_));
 sg13g2_o21ai_1 _19619_ (.B1(_02686_),
    .Y(_00524_),
    .A1(net39),
    .A2(_02685_));
 sg13g2_nor2b_1 _19620_ (.A(_12550_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_02687_));
 sg13g2_a21oi_1 _19621_ (.A1(net962),
    .A2(_12550_),
    .Y(_02688_),
    .B1(_02687_));
 sg13g2_nand2_1 _19622_ (.Y(_02689_),
    .A(net857),
    .B(_12548_));
 sg13g2_o21ai_1 _19623_ (.B1(_02689_),
    .Y(_00525_),
    .A1(_12548_),
    .A2(_02688_));
 sg13g2_nor2_1 _19624_ (.A(_12544_),
    .B(_11862_),
    .Y(_02690_));
 sg13g2_buf_2 _19625_ (.A(_02690_),
    .X(_02691_));
 sg13g2_nor2b_1 _19626_ (.A(_02691_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_02692_));
 sg13g2_a21oi_1 _19627_ (.A1(net963),
    .A2(_02691_),
    .Y(_02693_),
    .B1(_02692_));
 sg13g2_nand2_1 _19628_ (.Y(_02694_),
    .A(_12173_),
    .B(_12575_));
 sg13g2_o21ai_1 _19629_ (.B1(_02694_),
    .Y(_00526_),
    .A1(net39),
    .A2(_02693_));
 sg13g2_nor2b_1 _19630_ (.A(_02691_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_02695_));
 sg13g2_a21oi_1 _19631_ (.A1(net962),
    .A2(_02691_),
    .Y(_02696_),
    .B1(_02695_));
 sg13g2_nand2_1 _19632_ (.Y(_02697_),
    .A(_12177_),
    .B(_12575_));
 sg13g2_o21ai_1 _19633_ (.B1(_02697_),
    .Y(_00527_),
    .A1(_12576_),
    .A2(_02696_));
 sg13g2_nor2b_1 _19634_ (.A(_02691_),
    .B_N(\cpu.dcache.r_data[6][22] ),
    .Y(_02698_));
 sg13g2_a21oi_1 _19635_ (.A1(net961),
    .A2(_02691_),
    .Y(_02699_),
    .B1(_02698_));
 sg13g2_nand2_1 _19636_ (.Y(_02700_),
    .A(_12181_),
    .B(_12575_));
 sg13g2_o21ai_1 _19637_ (.B1(_02700_),
    .Y(_00528_),
    .A1(net39),
    .A2(_02699_));
 sg13g2_nor2b_1 _19638_ (.A(_02691_),
    .B_N(\cpu.dcache.r_data[6][23] ),
    .Y(_02701_));
 sg13g2_a21oi_1 _19639_ (.A1(net960),
    .A2(_02691_),
    .Y(_02702_),
    .B1(_02701_));
 sg13g2_nand2_1 _19640_ (.Y(_02703_),
    .A(_12058_),
    .B(_12575_));
 sg13g2_o21ai_1 _19641_ (.B1(_02703_),
    .Y(_00529_),
    .A1(_12576_),
    .A2(_02702_));
 sg13g2_nor2_1 _19642_ (.A(net480),
    .B(_12009_),
    .Y(_02704_));
 sg13g2_buf_1 _19643_ (.A(_02704_),
    .X(_02705_));
 sg13g2_buf_1 _19644_ (.A(_02705_),
    .X(_02706_));
 sg13g2_nor2_1 _19645_ (.A(net533),
    .B(_12015_),
    .Y(_02707_));
 sg13g2_buf_1 _19646_ (.A(_02707_),
    .X(_02708_));
 sg13g2_nor2b_1 _19647_ (.A(net418),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02709_));
 sg13g2_a21oi_1 _19648_ (.A1(_12490_),
    .A2(net418),
    .Y(_02710_),
    .B1(_02709_));
 sg13g2_nand2_1 _19649_ (.Y(_02711_),
    .A(_11876_),
    .B(_02706_));
 sg13g2_o21ai_1 _19650_ (.B1(_02711_),
    .Y(_00530_),
    .A1(_02706_),
    .A2(_02710_));
 sg13g2_nor2b_1 _19651_ (.A(net418),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02712_));
 sg13g2_a21oi_1 _19652_ (.A1(_12496_),
    .A2(net418),
    .Y(_02713_),
    .B1(_02712_));
 sg13g2_nand2_1 _19653_ (.Y(_02714_),
    .A(_11884_),
    .B(net38));
 sg13g2_o21ai_1 _19654_ (.B1(_02714_),
    .Y(_00531_),
    .A1(net38),
    .A2(_02713_));
 sg13g2_nor2b_1 _19655_ (.A(net418),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02715_));
 sg13g2_a21oi_1 _19656_ (.A1(_12500_),
    .A2(net418),
    .Y(_02716_),
    .B1(_02715_));
 sg13g2_nand2_1 _19657_ (.Y(_02717_),
    .A(_11805_),
    .B(_02705_));
 sg13g2_o21ai_1 _19658_ (.B1(_02717_),
    .Y(_00532_),
    .A1(net38),
    .A2(_02716_));
 sg13g2_nor2b_1 _19659_ (.A(_02708_),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02718_));
 sg13g2_a21oi_1 _19660_ (.A1(_12504_),
    .A2(_02708_),
    .Y(_02719_),
    .B1(_02718_));
 sg13g2_nand2_1 _19661_ (.Y(_02720_),
    .A(_11815_),
    .B(_02705_));
 sg13g2_o21ai_1 _19662_ (.B1(_02720_),
    .Y(_00533_),
    .A1(net38),
    .A2(_02719_));
 sg13g2_nor2_2 _19663_ (.A(_12545_),
    .B(_11890_),
    .Y(_02721_));
 sg13g2_mux2_1 _19664_ (.A0(\cpu.dcache.r_data[6][28] ),
    .A1(net1076),
    .S(_02721_),
    .X(_02722_));
 sg13g2_nor2_1 _19665_ (.A(_02705_),
    .B(_02722_),
    .Y(_02723_));
 sg13g2_a21oi_1 _19666_ (.A1(_11820_),
    .A2(net38),
    .Y(_00534_),
    .B1(_02723_));
 sg13g2_mux2_1 _19667_ (.A0(\cpu.dcache.r_data[6][29] ),
    .A1(net1069),
    .S(_02721_),
    .X(_02724_));
 sg13g2_nor2_1 _19668_ (.A(_02705_),
    .B(_02724_),
    .Y(_02725_));
 sg13g2_a21oi_1 _19669_ (.A1(_11830_),
    .A2(net38),
    .Y(_00535_),
    .B1(_02725_));
 sg13g2_nor2b_1 _19670_ (.A(_12550_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02726_));
 sg13g2_a21oi_1 _19671_ (.A1(net961),
    .A2(_12550_),
    .Y(_02727_),
    .B1(_02726_));
 sg13g2_nand2_1 _19672_ (.Y(_02728_),
    .A(net856),
    .B(_12547_));
 sg13g2_o21ai_1 _19673_ (.B1(_02728_),
    .Y(_00536_),
    .A1(net41),
    .A2(_02727_));
 sg13g2_mux2_1 _19674_ (.A0(\cpu.dcache.r_data[6][30] ),
    .A1(net1075),
    .S(_02721_),
    .X(_02729_));
 sg13g2_nor2_1 _19675_ (.A(_02705_),
    .B(_02729_),
    .Y(_02730_));
 sg13g2_a21oi_1 _19676_ (.A1(_11837_),
    .A2(net38),
    .Y(_00537_),
    .B1(_02730_));
 sg13g2_mux2_1 _19677_ (.A0(\cpu.dcache.r_data[6][31] ),
    .A1(net1074),
    .S(_02721_),
    .X(_02731_));
 sg13g2_nor2_1 _19678_ (.A(_02705_),
    .B(_02731_),
    .Y(_02732_));
 sg13g2_a21oi_1 _19679_ (.A1(_11842_),
    .A2(net38),
    .Y(_00538_),
    .B1(_02732_));
 sg13g2_nor2b_1 _19680_ (.A(_12550_),
    .B_N(\cpu.dcache.r_data[6][3] ),
    .Y(_02733_));
 sg13g2_a21oi_1 _19681_ (.A1(net960),
    .A2(_12550_),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nand2_1 _19682_ (.Y(_02735_),
    .A(_12358_),
    .B(_12547_));
 sg13g2_o21ai_1 _19683_ (.B1(_02735_),
    .Y(_00539_),
    .A1(net41),
    .A2(_02734_));
 sg13g2_nor2_1 _19684_ (.A(net533),
    .B(_11907_),
    .Y(_02736_));
 sg13g2_buf_2 _19685_ (.A(_02736_),
    .X(_02737_));
 sg13g2_nor2b_1 _19686_ (.A(_02737_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02738_));
 sg13g2_a21oi_1 _19687_ (.A1(net963),
    .A2(_02737_),
    .Y(_02739_),
    .B1(_02738_));
 sg13g2_nand2_1 _19688_ (.Y(_02740_),
    .A(net971),
    .B(_12547_));
 sg13g2_o21ai_1 _19689_ (.B1(_02740_),
    .Y(_00540_),
    .A1(net41),
    .A2(_02739_));
 sg13g2_nor2b_1 _19690_ (.A(_02737_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02741_));
 sg13g2_a21oi_1 _19691_ (.A1(net962),
    .A2(_02737_),
    .Y(_02742_),
    .B1(_02741_));
 sg13g2_nand2_1 _19692_ (.Y(_02743_),
    .A(net970),
    .B(_12547_));
 sg13g2_o21ai_1 _19693_ (.B1(_02743_),
    .Y(_00541_),
    .A1(net41),
    .A2(_02742_));
 sg13g2_nor2b_1 _19694_ (.A(_02737_),
    .B_N(\cpu.dcache.r_data[6][6] ),
    .Y(_02744_));
 sg13g2_a21oi_1 _19695_ (.A1(net961),
    .A2(_02737_),
    .Y(_02745_),
    .B1(_02744_));
 sg13g2_nand2_1 _19696_ (.Y(_02746_),
    .A(net969),
    .B(_12547_));
 sg13g2_o21ai_1 _19697_ (.B1(_02746_),
    .Y(_00542_),
    .A1(net41),
    .A2(_02745_));
 sg13g2_nor2b_1 _19698_ (.A(_02737_),
    .B_N(\cpu.dcache.r_data[6][7] ),
    .Y(_02747_));
 sg13g2_a21oi_1 _19699_ (.A1(net960),
    .A2(_02737_),
    .Y(_02748_),
    .B1(_02747_));
 sg13g2_nand2_1 _19700_ (.Y(_02749_),
    .A(_10000_),
    .B(_12547_));
 sg13g2_o21ai_1 _19701_ (.B1(_02749_),
    .Y(_00543_),
    .A1(net41),
    .A2(_02748_));
 sg13g2_nor2b_1 _19702_ (.A(_12558_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02750_));
 sg13g2_a21oi_1 _19703_ (.A1(net963),
    .A2(_12558_),
    .Y(_02751_),
    .B1(_02750_));
 sg13g2_nand2_1 _19704_ (.Y(_02752_),
    .A(_11876_),
    .B(_12555_));
 sg13g2_o21ai_1 _19705_ (.B1(_02752_),
    .Y(_00544_),
    .A1(net40),
    .A2(_02751_));
 sg13g2_nor2b_1 _19706_ (.A(_12558_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02753_));
 sg13g2_a21oi_1 _19707_ (.A1(_12496_),
    .A2(_12558_),
    .Y(_02754_),
    .B1(_02753_));
 sg13g2_nand2_1 _19708_ (.Y(_02755_),
    .A(_11884_),
    .B(_12555_));
 sg13g2_o21ai_1 _19709_ (.B1(_02755_),
    .Y(_00545_),
    .A1(net40),
    .A2(_02754_));
 sg13g2_buf_1 _19710_ (.A(_09817_),
    .X(_02756_));
 sg13g2_nor2_1 _19711_ (.A(net479),
    .B(_11920_),
    .Y(_02757_));
 sg13g2_buf_2 _19712_ (.A(_02757_),
    .X(_02758_));
 sg13g2_buf_1 _19713_ (.A(_02758_),
    .X(_02759_));
 sg13g2_nor2_1 _19714_ (.A(net479),
    .B(_11774_),
    .Y(_02760_));
 sg13g2_buf_2 _19715_ (.A(_02760_),
    .X(_02761_));
 sg13g2_nor2b_1 _19716_ (.A(_02761_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02762_));
 sg13g2_a21oi_1 _19717_ (.A1(net963),
    .A2(_02761_),
    .Y(_02763_),
    .B1(_02762_));
 sg13g2_nand2_1 _19718_ (.Y(_02764_),
    .A(_12581_),
    .B(net37));
 sg13g2_o21ai_1 _19719_ (.B1(_02764_),
    .Y(_00546_),
    .A1(_02759_),
    .A2(_02763_));
 sg13g2_nor2_1 _19720_ (.A(net479),
    .B(_11933_),
    .Y(_02765_));
 sg13g2_buf_1 _19721_ (.A(_02765_),
    .X(_02766_));
 sg13g2_buf_1 _19722_ (.A(_02766_),
    .X(_02767_));
 sg13g2_nor2_1 _19723_ (.A(net479),
    .B(_11797_),
    .Y(_02768_));
 sg13g2_buf_2 _19724_ (.A(_02768_),
    .X(_02769_));
 sg13g2_nor2b_1 _19725_ (.A(_02769_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02770_));
 sg13g2_a21oi_1 _19726_ (.A1(net961),
    .A2(_02769_),
    .Y(_02771_),
    .B1(_02770_));
 sg13g2_nand2_1 _19727_ (.Y(_02772_),
    .A(_11805_),
    .B(net36));
 sg13g2_o21ai_1 _19728_ (.B1(_02772_),
    .Y(_00547_),
    .A1(net36),
    .A2(_02771_));
 sg13g2_nor2b_1 _19729_ (.A(_02769_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02773_));
 sg13g2_a21oi_1 _19730_ (.A1(_12504_),
    .A2(_02769_),
    .Y(_02774_),
    .B1(_02773_));
 sg13g2_nand2_1 _19731_ (.Y(_02775_),
    .A(_11815_),
    .B(net36));
 sg13g2_o21ai_1 _19732_ (.B1(_02775_),
    .Y(_00548_),
    .A1(net36),
    .A2(_02774_));
 sg13g2_nor2_2 _19733_ (.A(net479),
    .B(_11823_),
    .Y(_02776_));
 sg13g2_mux2_1 _19734_ (.A0(\cpu.dcache.r_data[7][12] ),
    .A1(_11924_),
    .S(_02776_),
    .X(_02777_));
 sg13g2_nor2_1 _19735_ (.A(_02766_),
    .B(_02777_),
    .Y(_02778_));
 sg13g2_a21oi_1 _19736_ (.A1(_11820_),
    .A2(net36),
    .Y(_00549_),
    .B1(_02778_));
 sg13g2_mux2_1 _19737_ (.A0(\cpu.dcache.r_data[7][13] ),
    .A1(net1069),
    .S(_02776_),
    .X(_02779_));
 sg13g2_nor2_1 _19738_ (.A(_02766_),
    .B(_02779_),
    .Y(_02780_));
 sg13g2_a21oi_1 _19739_ (.A1(_11830_),
    .A2(_02767_),
    .Y(_00550_),
    .B1(_02780_));
 sg13g2_mux2_1 _19740_ (.A0(\cpu.dcache.r_data[7][14] ),
    .A1(_11937_),
    .S(_02776_),
    .X(_02781_));
 sg13g2_nor2_1 _19741_ (.A(_02766_),
    .B(_02781_),
    .Y(_02782_));
 sg13g2_a21oi_1 _19742_ (.A1(_11837_),
    .A2(_02767_),
    .Y(_00551_),
    .B1(_02782_));
 sg13g2_mux2_1 _19743_ (.A0(\cpu.dcache.r_data[7][15] ),
    .A1(net1074),
    .S(_02776_),
    .X(_02783_));
 sg13g2_nor2_1 _19744_ (.A(_02766_),
    .B(_02783_),
    .Y(_02784_));
 sg13g2_a21oi_1 _19745_ (.A1(_11842_),
    .A2(net36),
    .Y(_00552_),
    .B1(_02784_));
 sg13g2_nor2_1 _19746_ (.A(net479),
    .B(_11963_),
    .Y(_02785_));
 sg13g2_buf_2 _19747_ (.A(_02785_),
    .X(_02786_));
 sg13g2_buf_1 _19748_ (.A(_02786_),
    .X(_02787_));
 sg13g2_buf_2 _19749_ (.A(net1076),
    .X(_02788_));
 sg13g2_nor2_1 _19750_ (.A(net479),
    .B(_11846_),
    .Y(_02789_));
 sg13g2_buf_2 _19751_ (.A(_02789_),
    .X(_02790_));
 sg13g2_nor2b_1 _19752_ (.A(_02790_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02791_));
 sg13g2_a21oi_1 _19753_ (.A1(net958),
    .A2(_02790_),
    .Y(_02792_),
    .B1(_02791_));
 sg13g2_nand2_1 _19754_ (.Y(_02793_),
    .A(net959),
    .B(net35));
 sg13g2_o21ai_1 _19755_ (.B1(_02793_),
    .Y(_00553_),
    .A1(net35),
    .A2(_02792_));
 sg13g2_nor2b_1 _19756_ (.A(_02790_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02794_));
 sg13g2_a21oi_1 _19757_ (.A1(net962),
    .A2(_02790_),
    .Y(_02795_),
    .B1(_02794_));
 sg13g2_nand2_1 _19758_ (.Y(_02796_),
    .A(net857),
    .B(net35));
 sg13g2_o21ai_1 _19759_ (.B1(_02796_),
    .Y(_00554_),
    .A1(_02787_),
    .A2(_02795_));
 sg13g2_buf_2 _19760_ (.A(net1075),
    .X(_02797_));
 sg13g2_nor2b_1 _19761_ (.A(_02790_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02798_));
 sg13g2_a21oi_1 _19762_ (.A1(net957),
    .A2(_02790_),
    .Y(_02799_),
    .B1(_02798_));
 sg13g2_nand2_1 _19763_ (.Y(_02800_),
    .A(net856),
    .B(_02786_));
 sg13g2_o21ai_1 _19764_ (.B1(_02800_),
    .Y(_00555_),
    .A1(net35),
    .A2(_02799_));
 sg13g2_buf_2 _19765_ (.A(net1074),
    .X(_02801_));
 sg13g2_nor2b_1 _19766_ (.A(_02790_),
    .B_N(\cpu.dcache.r_data[7][19] ),
    .Y(_02802_));
 sg13g2_a21oi_1 _19767_ (.A1(net956),
    .A2(_02790_),
    .Y(_02803_),
    .B1(_02802_));
 sg13g2_nand2_1 _19768_ (.Y(_02804_),
    .A(net964),
    .B(_02786_));
 sg13g2_o21ai_1 _19769_ (.B1(_02804_),
    .Y(_00556_),
    .A1(net35),
    .A2(_02803_));
 sg13g2_buf_2 _19770_ (.A(net1069),
    .X(_02805_));
 sg13g2_nor2b_1 _19771_ (.A(_02761_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02806_));
 sg13g2_a21oi_1 _19772_ (.A1(net955),
    .A2(_02761_),
    .Y(_02807_),
    .B1(_02806_));
 sg13g2_buf_1 _19773_ (.A(_09904_),
    .X(_02808_));
 sg13g2_nand2_1 _19774_ (.Y(_02809_),
    .A(net954),
    .B(net37));
 sg13g2_o21ai_1 _19775_ (.B1(_02809_),
    .Y(_00557_),
    .A1(net37),
    .A2(_02807_));
 sg13g2_nor2_1 _19776_ (.A(_09817_),
    .B(_11862_),
    .Y(_02810_));
 sg13g2_buf_2 _19777_ (.A(_02810_),
    .X(_02811_));
 sg13g2_nor2b_1 _19778_ (.A(_02811_),
    .B_N(\cpu.dcache.r_data[7][20] ),
    .Y(_02812_));
 sg13g2_a21oi_1 _19779_ (.A1(net958),
    .A2(_02811_),
    .Y(_02813_),
    .B1(_02812_));
 sg13g2_nand2_1 _19780_ (.Y(_02814_),
    .A(net971),
    .B(_02786_));
 sg13g2_o21ai_1 _19781_ (.B1(_02814_),
    .Y(_00558_),
    .A1(_02787_),
    .A2(_02813_));
 sg13g2_nor2b_1 _19782_ (.A(_02811_),
    .B_N(\cpu.dcache.r_data[7][21] ),
    .Y(_02815_));
 sg13g2_a21oi_1 _19783_ (.A1(net955),
    .A2(_02811_),
    .Y(_02816_),
    .B1(_02815_));
 sg13g2_nand2_1 _19784_ (.Y(_02817_),
    .A(net970),
    .B(_02786_));
 sg13g2_o21ai_1 _19785_ (.B1(_02817_),
    .Y(_00559_),
    .A1(net35),
    .A2(_02816_));
 sg13g2_nor2b_1 _19786_ (.A(_02811_),
    .B_N(\cpu.dcache.r_data[7][22] ),
    .Y(_02818_));
 sg13g2_a21oi_1 _19787_ (.A1(net957),
    .A2(_02811_),
    .Y(_02819_),
    .B1(_02818_));
 sg13g2_nand2_1 _19788_ (.Y(_02820_),
    .A(net969),
    .B(_02786_));
 sg13g2_o21ai_1 _19789_ (.B1(_02820_),
    .Y(_00560_),
    .A1(net35),
    .A2(_02819_));
 sg13g2_nor2b_1 _19790_ (.A(_02811_),
    .B_N(\cpu.dcache.r_data[7][23] ),
    .Y(_02821_));
 sg13g2_a21oi_1 _19791_ (.A1(net956),
    .A2(_02811_),
    .Y(_02822_),
    .B1(_02821_));
 sg13g2_nand2_1 _19792_ (.Y(_02823_),
    .A(net1012),
    .B(_02786_));
 sg13g2_o21ai_1 _19793_ (.B1(_02823_),
    .Y(_00561_),
    .A1(net35),
    .A2(_02822_));
 sg13g2_nor2_1 _19794_ (.A(_02756_),
    .B(_12009_),
    .Y(_02824_));
 sg13g2_buf_1 _19795_ (.A(_02824_),
    .X(_02825_));
 sg13g2_buf_1 _19796_ (.A(_02825_),
    .X(_02826_));
 sg13g2_nor2_1 _19797_ (.A(_09817_),
    .B(_12015_),
    .Y(_02827_));
 sg13g2_buf_1 _19798_ (.A(_02827_),
    .X(_02828_));
 sg13g2_nor2b_1 _19799_ (.A(net417),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02829_));
 sg13g2_a21oi_1 _19800_ (.A1(net958),
    .A2(net417),
    .Y(_02830_),
    .B1(_02829_));
 sg13g2_nand2_1 _19801_ (.Y(_02831_),
    .A(_11876_),
    .B(net34));
 sg13g2_o21ai_1 _19802_ (.B1(_02831_),
    .Y(_00562_),
    .A1(net34),
    .A2(_02830_));
 sg13g2_nor2b_1 _19803_ (.A(net417),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02832_));
 sg13g2_a21oi_1 _19804_ (.A1(net955),
    .A2(net417),
    .Y(_02833_),
    .B1(_02832_));
 sg13g2_nand2_1 _19805_ (.Y(_02834_),
    .A(_11884_),
    .B(_02826_));
 sg13g2_o21ai_1 _19806_ (.B1(_02834_),
    .Y(_00563_),
    .A1(net34),
    .A2(_02833_));
 sg13g2_nor2b_1 _19807_ (.A(_02828_),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02835_));
 sg13g2_a21oi_1 _19808_ (.A1(net957),
    .A2(_02828_),
    .Y(_02836_),
    .B1(_02835_));
 sg13g2_nand2_1 _19809_ (.Y(_02837_),
    .A(_11805_),
    .B(_02825_));
 sg13g2_o21ai_1 _19810_ (.B1(_02837_),
    .Y(_00564_),
    .A1(net34),
    .A2(_02836_));
 sg13g2_nor2b_1 _19811_ (.A(net417),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02838_));
 sg13g2_a21oi_1 _19812_ (.A1(net956),
    .A2(net417),
    .Y(_02839_),
    .B1(_02838_));
 sg13g2_nand2_1 _19813_ (.Y(_02840_),
    .A(_11815_),
    .B(_02825_));
 sg13g2_o21ai_1 _19814_ (.B1(_02840_),
    .Y(_00565_),
    .A1(net34),
    .A2(_02839_));
 sg13g2_nor2_2 _19815_ (.A(_02756_),
    .B(_11890_),
    .Y(_02841_));
 sg13g2_mux2_1 _19816_ (.A0(\cpu.dcache.r_data[7][28] ),
    .A1(net1076),
    .S(_02841_),
    .X(_02842_));
 sg13g2_nor2_1 _19817_ (.A(_02825_),
    .B(_02842_),
    .Y(_02843_));
 sg13g2_a21oi_1 _19818_ (.A1(_11820_),
    .A2(net34),
    .Y(_00566_),
    .B1(_02843_));
 sg13g2_mux2_1 _19819_ (.A0(\cpu.dcache.r_data[7][29] ),
    .A1(net1069),
    .S(_02841_),
    .X(_02844_));
 sg13g2_nor2_1 _19820_ (.A(_02825_),
    .B(_02844_),
    .Y(_02845_));
 sg13g2_a21oi_1 _19821_ (.A1(_11830_),
    .A2(net34),
    .Y(_00567_),
    .B1(_02845_));
 sg13g2_nor2b_1 _19822_ (.A(_02761_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02846_));
 sg13g2_a21oi_1 _19823_ (.A1(net957),
    .A2(_02761_),
    .Y(_02847_),
    .B1(_02846_));
 sg13g2_buf_1 _19824_ (.A(net1018),
    .X(_02848_));
 sg13g2_nand2_1 _19825_ (.Y(_02849_),
    .A(net855),
    .B(_02758_));
 sg13g2_o21ai_1 _19826_ (.B1(_02849_),
    .Y(_00568_),
    .A1(net37),
    .A2(_02847_));
 sg13g2_mux2_1 _19827_ (.A0(\cpu.dcache.r_data[7][30] ),
    .A1(net1075),
    .S(_02841_),
    .X(_02850_));
 sg13g2_nor2_1 _19828_ (.A(_02825_),
    .B(_02850_),
    .Y(_02851_));
 sg13g2_a21oi_1 _19829_ (.A1(_11837_),
    .A2(net34),
    .Y(_00569_),
    .B1(_02851_));
 sg13g2_mux2_1 _19830_ (.A0(\cpu.dcache.r_data[7][31] ),
    .A1(_11944_),
    .S(_02841_),
    .X(_02852_));
 sg13g2_nor2_1 _19831_ (.A(_02825_),
    .B(_02852_),
    .Y(_02853_));
 sg13g2_a21oi_1 _19832_ (.A1(_11842_),
    .A2(_02826_),
    .Y(_00570_),
    .B1(_02853_));
 sg13g2_nor2b_1 _19833_ (.A(_02761_),
    .B_N(\cpu.dcache.r_data[7][3] ),
    .Y(_02854_));
 sg13g2_a21oi_1 _19834_ (.A1(net956),
    .A2(_02761_),
    .Y(_02855_),
    .B1(_02854_));
 sg13g2_nand2_1 _19835_ (.Y(_02856_),
    .A(net964),
    .B(_02758_));
 sg13g2_o21ai_1 _19836_ (.B1(_02856_),
    .Y(_00571_),
    .A1(net37),
    .A2(_02855_));
 sg13g2_nor2_1 _19837_ (.A(_09817_),
    .B(_11907_),
    .Y(_02857_));
 sg13g2_buf_2 _19838_ (.A(_02857_),
    .X(_02858_));
 sg13g2_nor2b_1 _19839_ (.A(_02858_),
    .B_N(\cpu.dcache.r_data[7][4] ),
    .Y(_02859_));
 sg13g2_a21oi_1 _19840_ (.A1(net958),
    .A2(_02858_),
    .Y(_02860_),
    .B1(_02859_));
 sg13g2_nand2_1 _19841_ (.Y(_02861_),
    .A(net1016),
    .B(_02758_));
 sg13g2_o21ai_1 _19842_ (.B1(_02861_),
    .Y(_00572_),
    .A1(net37),
    .A2(_02860_));
 sg13g2_nor2b_1 _19843_ (.A(_02858_),
    .B_N(\cpu.dcache.r_data[7][5] ),
    .Y(_02862_));
 sg13g2_a21oi_1 _19844_ (.A1(net955),
    .A2(_02858_),
    .Y(_02863_),
    .B1(_02862_));
 sg13g2_nand2_1 _19845_ (.Y(_02864_),
    .A(_09928_),
    .B(_02758_));
 sg13g2_o21ai_1 _19846_ (.B1(_02864_),
    .Y(_00573_),
    .A1(net37),
    .A2(_02863_));
 sg13g2_nor2b_1 _19847_ (.A(_02858_),
    .B_N(\cpu.dcache.r_data[7][6] ),
    .Y(_02865_));
 sg13g2_a21oi_1 _19848_ (.A1(net957),
    .A2(_02858_),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_nand2_1 _19849_ (.Y(_02867_),
    .A(_09934_),
    .B(_02758_));
 sg13g2_o21ai_1 _19850_ (.B1(_02867_),
    .Y(_00574_),
    .A1(net37),
    .A2(_02866_));
 sg13g2_nor2b_1 _19851_ (.A(_02858_),
    .B_N(\cpu.dcache.r_data[7][7] ),
    .Y(_02868_));
 sg13g2_a21oi_1 _19852_ (.A1(net956),
    .A2(_02858_),
    .Y(_02869_),
    .B1(_02868_));
 sg13g2_nand2_1 _19853_ (.Y(_02870_),
    .A(_10000_),
    .B(_02758_));
 sg13g2_o21ai_1 _19854_ (.B1(_02870_),
    .Y(_00575_),
    .A1(_02759_),
    .A2(_02869_));
 sg13g2_nor2b_1 _19855_ (.A(_02769_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_02871_));
 sg13g2_a21oi_1 _19856_ (.A1(net958),
    .A2(_02769_),
    .Y(_02872_),
    .B1(_02871_));
 sg13g2_nand2_1 _19857_ (.Y(_02873_),
    .A(_11876_),
    .B(_02766_));
 sg13g2_o21ai_1 _19858_ (.B1(_02873_),
    .Y(_00576_),
    .A1(net36),
    .A2(_02872_));
 sg13g2_nor2b_1 _19859_ (.A(_02769_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_02874_));
 sg13g2_a21oi_1 _19860_ (.A1(net955),
    .A2(_02769_),
    .Y(_02875_),
    .B1(_02874_));
 sg13g2_nand2_1 _19861_ (.Y(_02876_),
    .A(_11884_),
    .B(_02766_));
 sg13g2_o21ai_1 _19862_ (.B1(_02876_),
    .Y(_00577_),
    .A1(net36),
    .A2(_02875_));
 sg13g2_nand2_1 _19863_ (.Y(_02877_),
    .A(_09653_),
    .B(_11783_));
 sg13g2_buf_1 _19864_ (.A(_09107_),
    .X(_02878_));
 sg13g2_buf_1 _19865_ (.A(\cpu.d_rstrobe_d ),
    .X(_02879_));
 sg13g2_nand2b_1 _19866_ (.Y(_02880_),
    .B(net994),
    .A_N(_02879_));
 sg13g2_or4_1 _19867_ (.A(net854),
    .B(_09223_),
    .C(_08764_),
    .D(_02880_),
    .X(_02881_));
 sg13g2_nand2_1 _19868_ (.Y(_02882_),
    .A(_02877_),
    .B(_02881_));
 sg13g2_buf_2 _19869_ (.A(_02882_),
    .X(_02883_));
 sg13g2_xor2_1 _19870_ (.B(_11766_),
    .A(_02879_),
    .X(_02884_));
 sg13g2_nand3_1 _19871_ (.B(net863),
    .C(_02884_),
    .A(_12013_),
    .Y(_02885_));
 sg13g2_a21oi_1 _19872_ (.A1(_02885_),
    .A2(_02877_),
    .Y(_02886_),
    .B1(_11764_));
 sg13g2_mux2_1 _19873_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_02883_),
    .S(_02886_),
    .X(_00578_));
 sg13g2_buf_1 _19874_ (.A(net493),
    .X(_02887_));
 sg13g2_buf_1 _19875_ (.A(net416),
    .X(_02888_));
 sg13g2_nand2_1 _19876_ (.Y(_02889_),
    .A(_02885_),
    .B(_02877_));
 sg13g2_buf_2 _19877_ (.A(_02889_),
    .X(_02890_));
 sg13g2_nand2_1 _19878_ (.Y(_02891_),
    .A(net372),
    .B(_02890_));
 sg13g2_mux2_1 _19879_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[1] ),
    .S(_02891_),
    .X(_00579_));
 sg13g2_buf_1 _19880_ (.A(net548),
    .X(_02892_));
 sg13g2_buf_1 _19881_ (.A(_02892_),
    .X(_02893_));
 sg13g2_nand2_1 _19882_ (.Y(_02894_),
    .A(net415),
    .B(_02890_));
 sg13g2_mux2_1 _19883_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[2] ),
    .S(_02894_),
    .X(_00580_));
 sg13g2_buf_1 _19884_ (.A(net546),
    .X(_02895_));
 sg13g2_buf_1 _19885_ (.A(net477),
    .X(_02896_));
 sg13g2_nand2_1 _19886_ (.Y(_02897_),
    .A(net414),
    .B(_02890_));
 sg13g2_mux2_1 _19887_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[3] ),
    .S(_02897_),
    .X(_00581_));
 sg13g2_nand2_1 _19888_ (.Y(_02898_),
    .A(net598),
    .B(_02890_));
 sg13g2_mux2_1 _19889_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[4] ),
    .S(_02898_),
    .X(_00582_));
 sg13g2_buf_1 _19890_ (.A(net545),
    .X(_02899_));
 sg13g2_buf_1 _19891_ (.A(net476),
    .X(_02900_));
 sg13g2_nand2_1 _19892_ (.Y(_02901_),
    .A(_02900_),
    .B(_02890_));
 sg13g2_mux2_1 _19893_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[5] ),
    .S(_02901_),
    .X(_00583_));
 sg13g2_buf_1 _19894_ (.A(net612),
    .X(_02902_));
 sg13g2_buf_1 _19895_ (.A(net532),
    .X(_02903_));
 sg13g2_nand2_1 _19896_ (.Y(_02904_),
    .A(net475),
    .B(_02890_));
 sg13g2_mux2_1 _19897_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[6] ),
    .S(_02904_),
    .X(_00584_));
 sg13g2_buf_1 _19898_ (.A(_09391_),
    .X(_02905_));
 sg13g2_buf_1 _19899_ (.A(net531),
    .X(_02906_));
 sg13g2_nand2_1 _19900_ (.Y(_02907_),
    .A(_02906_),
    .B(_02890_));
 sg13g2_mux2_1 _19901_ (.A0(_02883_),
    .A1(\cpu.dcache.r_dirty[7] ),
    .S(_02907_),
    .X(_00585_));
 sg13g2_buf_1 _19902_ (.A(net865),
    .X(_02908_));
 sg13g2_buf_1 _19903_ (.A(_11873_),
    .X(_02909_));
 sg13g2_buf_1 _19904_ (.A(_11873_),
    .X(_02910_));
 sg13g2_nand2_1 _19905_ (.Y(_02911_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(_02910_));
 sg13g2_o21ai_1 _19906_ (.B1(_02911_),
    .Y(_00589_),
    .A1(net729),
    .A2(net337));
 sg13g2_mux2_1 _19907_ (.A0(net438),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(net337),
    .X(_00590_));
 sg13g2_mux2_1 _19908_ (.A0(net435),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net337),
    .X(_00591_));
 sg13g2_mux2_1 _19909_ (.A0(net432),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(_02909_),
    .X(_00592_));
 sg13g2_mux2_1 _19910_ (.A0(net439),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net337),
    .X(_00593_));
 sg13g2_mux2_1 _19911_ (.A0(net433),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net337),
    .X(_00594_));
 sg13g2_mux2_1 _19912_ (.A0(net430),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(net337),
    .X(_00595_));
 sg13g2_mux2_1 _19913_ (.A0(net434),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net337),
    .X(_00596_));
 sg13g2_mux2_1 _19914_ (.A0(net431),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(_02909_),
    .X(_00597_));
 sg13g2_inv_1 _19915_ (.Y(_02912_),
    .A(net437));
 sg13g2_nand2_1 _19916_ (.Y(_02913_),
    .A(\cpu.dcache.r_tag[0][23] ),
    .B(_11873_));
 sg13g2_o21ai_1 _19917_ (.B1(_02913_),
    .Y(_00598_),
    .A1(_02912_),
    .A2(net337));
 sg13g2_buf_2 _19918_ (.A(_09010_),
    .X(_02914_));
 sg13g2_buf_1 _19919_ (.A(net953),
    .X(_02915_));
 sg13g2_buf_2 _19920_ (.A(net853),
    .X(_02916_));
 sg13g2_mux2_1 _19921_ (.A0(net728),
    .A1(\cpu.dcache.r_tag[0][6] ),
    .S(net336),
    .X(_00599_));
 sg13g2_buf_1 _19922_ (.A(net1037),
    .X(_02917_));
 sg13g2_buf_2 _19923_ (.A(net852),
    .X(_02918_));
 sg13g2_mux2_1 _19924_ (.A0(net727),
    .A1(\cpu.dcache.r_tag[0][7] ),
    .S(net336),
    .X(_00600_));
 sg13g2_buf_1 _19925_ (.A(net1038),
    .X(_02919_));
 sg13g2_buf_2 _19926_ (.A(net851),
    .X(_02920_));
 sg13g2_mux2_1 _19927_ (.A0(net726),
    .A1(\cpu.dcache.r_tag[0][8] ),
    .S(net336),
    .X(_00601_));
 sg13g2_buf_1 _19928_ (.A(_10627_),
    .X(_02921_));
 sg13g2_buf_2 _19929_ (.A(net952),
    .X(_02922_));
 sg13g2_mux2_1 _19930_ (.A0(net850),
    .A1(\cpu.dcache.r_tag[0][9] ),
    .S(_02910_),
    .X(_00602_));
 sg13g2_buf_1 _19931_ (.A(_10652_),
    .X(_02923_));
 sg13g2_buf_2 _19932_ (.A(net951),
    .X(_02924_));
 sg13g2_mux2_1 _19933_ (.A0(net849),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(net336),
    .X(_00603_));
 sg13g2_buf_1 _19934_ (.A(_10078_),
    .X(_02925_));
 sg13g2_buf_1 _19935_ (.A(net950),
    .X(_02926_));
 sg13g2_mux2_1 _19936_ (.A0(net848),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(net336),
    .X(_00604_));
 sg13g2_mux2_1 _19937_ (.A0(net344),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net336),
    .X(_00605_));
 sg13g2_mux2_1 _19938_ (.A0(net376),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(net336),
    .X(_00606_));
 sg13g2_mux2_1 _19939_ (.A0(net436),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net336),
    .X(_00607_));
 sg13g2_buf_2 _19940_ (.A(_11726_),
    .X(_02927_));
 sg13g2_buf_1 _19941_ (.A(net643),
    .X(_02928_));
 sg13g2_buf_1 _19942_ (.A(_12017_),
    .X(_02929_));
 sg13g2_mux2_1 _19943_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net596),
    .S(net412),
    .X(_00608_));
 sg13g2_mux2_1 _19944_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net438),
    .S(net412),
    .X(_00609_));
 sg13g2_mux2_1 _19945_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net435),
    .S(net412),
    .X(_00610_));
 sg13g2_mux2_1 _19946_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net432),
    .S(net412),
    .X(_00611_));
 sg13g2_mux2_1 _19947_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net439),
    .S(net412),
    .X(_00612_));
 sg13g2_mux2_1 _19948_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net433),
    .S(net412),
    .X(_00613_));
 sg13g2_mux2_1 _19949_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net430),
    .S(_02929_),
    .X(_00614_));
 sg13g2_mux2_1 _19950_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net434),
    .S(net412),
    .X(_00615_));
 sg13g2_mux2_1 _19951_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net431),
    .S(net412),
    .X(_00616_));
 sg13g2_mux2_1 _19952_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(net437),
    .S(_02929_),
    .X(_00617_));
 sg13g2_buf_1 _19953_ (.A(net853),
    .X(_02930_));
 sg13g2_buf_1 _19954_ (.A(net483),
    .X(_02931_));
 sg13g2_mux2_1 _19955_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net725),
    .S(net411),
    .X(_00618_));
 sg13g2_buf_1 _19956_ (.A(net852),
    .X(_02932_));
 sg13g2_mux2_1 _19957_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(_02932_),
    .S(net411),
    .X(_00619_));
 sg13g2_buf_1 _19958_ (.A(net851),
    .X(_02933_));
 sg13g2_mux2_1 _19959_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net723),
    .S(_02931_),
    .X(_00620_));
 sg13g2_buf_1 _19960_ (.A(net952),
    .X(_02934_));
 sg13g2_mux2_1 _19961_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net847),
    .S(net411),
    .X(_00621_));
 sg13g2_buf_1 _19962_ (.A(net951),
    .X(_02935_));
 sg13g2_mux2_1 _19963_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net846),
    .S(net411),
    .X(_00622_));
 sg13g2_buf_1 _19964_ (.A(net950),
    .X(_02936_));
 sg13g2_mux2_1 _19965_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(_02936_),
    .S(_02931_),
    .X(_00623_));
 sg13g2_mux2_1 _19966_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net344),
    .S(net411),
    .X(_00624_));
 sg13g2_mux2_1 _19967_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net376),
    .S(net411),
    .X(_00625_));
 sg13g2_mux2_1 _19968_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net436),
    .S(net411),
    .X(_00626_));
 sg13g2_buf_1 _19969_ (.A(net535),
    .X(_02937_));
 sg13g2_mux2_1 _19970_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net596),
    .S(net473),
    .X(_00627_));
 sg13g2_mux2_1 _19971_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net438),
    .S(net473),
    .X(_00628_));
 sg13g2_mux2_1 _19972_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net435),
    .S(net473),
    .X(_00629_));
 sg13g2_mux2_1 _19973_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net432),
    .S(_02937_),
    .X(_00630_));
 sg13g2_mux2_1 _19974_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net439),
    .S(net473),
    .X(_00631_));
 sg13g2_mux2_1 _19975_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net433),
    .S(net473),
    .X(_00632_));
 sg13g2_mux2_1 _19976_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net430),
    .S(net473),
    .X(_00633_));
 sg13g2_mux2_1 _19977_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net434),
    .S(net473),
    .X(_00634_));
 sg13g2_mux2_1 _19978_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net431),
    .S(net473),
    .X(_00635_));
 sg13g2_mux2_1 _19979_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(net437),
    .S(_02937_),
    .X(_00636_));
 sg13g2_buf_1 _19980_ (.A(net853),
    .X(_02938_));
 sg13g2_buf_1 _19981_ (.A(net535),
    .X(_02939_));
 sg13g2_mux2_1 _19982_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net722),
    .S(net472),
    .X(_00637_));
 sg13g2_buf_1 _19983_ (.A(net852),
    .X(_02940_));
 sg13g2_mux2_1 _19984_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net721),
    .S(net472),
    .X(_00638_));
 sg13g2_buf_1 _19985_ (.A(net851),
    .X(_02941_));
 sg13g2_mux2_1 _19986_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net720),
    .S(net472),
    .X(_00639_));
 sg13g2_buf_1 _19987_ (.A(net952),
    .X(_02942_));
 sg13g2_mux2_1 _19988_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net844),
    .S(net472),
    .X(_00640_));
 sg13g2_buf_1 _19989_ (.A(net951),
    .X(_02943_));
 sg13g2_mux2_1 _19990_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net843),
    .S(_02939_),
    .X(_00641_));
 sg13g2_buf_1 _19991_ (.A(net950),
    .X(_02944_));
 sg13g2_mux2_1 _19992_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net842),
    .S(_02939_),
    .X(_00642_));
 sg13g2_mux2_1 _19993_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net344),
    .S(net472),
    .X(_00643_));
 sg13g2_mux2_1 _19994_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net376),
    .S(net472),
    .X(_00644_));
 sg13g2_mux2_1 _19995_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(_09493_),
    .S(net472),
    .X(_00645_));
 sg13g2_buf_1 _19996_ (.A(_12261_),
    .X(_02945_));
 sg13g2_mux2_1 _19997_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net596),
    .S(_02945_),
    .X(_00646_));
 sg13g2_mux2_1 _19998_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net438),
    .S(net371),
    .X(_00647_));
 sg13g2_mux2_1 _19999_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net435),
    .S(net371),
    .X(_00648_));
 sg13g2_mux2_1 _20000_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net432),
    .S(_02945_),
    .X(_00649_));
 sg13g2_mux2_1 _20001_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net439),
    .S(net371),
    .X(_00650_));
 sg13g2_mux2_1 _20002_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(net433),
    .S(net371),
    .X(_00651_));
 sg13g2_mux2_1 _20003_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(_09631_),
    .S(net371),
    .X(_00652_));
 sg13g2_mux2_1 _20004_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net434),
    .S(net371),
    .X(_00653_));
 sg13g2_mux2_1 _20005_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net431),
    .S(net371),
    .X(_00654_));
 sg13g2_mux2_1 _20006_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(net437),
    .S(net371),
    .X(_00655_));
 sg13g2_buf_1 _20007_ (.A(_12261_),
    .X(_02946_));
 sg13g2_mux2_1 _20008_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net722),
    .S(net370),
    .X(_00656_));
 sg13g2_mux2_1 _20009_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net721),
    .S(net370),
    .X(_00657_));
 sg13g2_mux2_1 _20010_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net720),
    .S(net370),
    .X(_00658_));
 sg13g2_mux2_1 _20011_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net844),
    .S(net370),
    .X(_00659_));
 sg13g2_mux2_1 _20012_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net843),
    .S(_02946_),
    .X(_00660_));
 sg13g2_mux2_1 _20013_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net842),
    .S(_02946_),
    .X(_00661_));
 sg13g2_mux2_1 _20014_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net344),
    .S(net370),
    .X(_00662_));
 sg13g2_mux2_1 _20015_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(_09316_),
    .S(net370),
    .X(_00663_));
 sg13g2_mux2_1 _20016_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(_09493_),
    .S(net370),
    .X(_00664_));
 sg13g2_buf_1 _20017_ (.A(_12380_),
    .X(_02947_));
 sg13g2_buf_1 _20018_ (.A(_12380_),
    .X(_02948_));
 sg13g2_nand2_1 _20019_ (.Y(_02949_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net409));
 sg13g2_o21ai_1 _20020_ (.B1(_02949_),
    .Y(_00665_),
    .A1(net729),
    .A2(net410));
 sg13g2_mux2_1 _20021_ (.A0(net438),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net410),
    .X(_00666_));
 sg13g2_mux2_1 _20022_ (.A0(net435),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net410),
    .X(_00667_));
 sg13g2_mux2_1 _20023_ (.A0(net432),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(_02947_),
    .X(_00668_));
 sg13g2_mux2_1 _20024_ (.A0(net439),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net410),
    .X(_00669_));
 sg13g2_mux2_1 _20025_ (.A0(net433),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net410),
    .X(_00670_));
 sg13g2_mux2_1 _20026_ (.A0(net430),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(_02947_),
    .X(_00671_));
 sg13g2_mux2_1 _20027_ (.A0(net434),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net410),
    .X(_00672_));
 sg13g2_mux2_1 _20028_ (.A0(net431),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(net410),
    .X(_00673_));
 sg13g2_nand2_1 _20029_ (.Y(_02950_),
    .A(\cpu.dcache.r_tag[4][23] ),
    .B(_12380_));
 sg13g2_o21ai_1 _20030_ (.B1(_02950_),
    .Y(_00674_),
    .A1(_02912_),
    .A2(net410));
 sg13g2_mux2_1 _20031_ (.A0(net728),
    .A1(\cpu.dcache.r_tag[4][6] ),
    .S(net409),
    .X(_00675_));
 sg13g2_mux2_1 _20032_ (.A0(net727),
    .A1(\cpu.dcache.r_tag[4][7] ),
    .S(net409),
    .X(_00676_));
 sg13g2_mux2_1 _20033_ (.A0(net726),
    .A1(\cpu.dcache.r_tag[4][8] ),
    .S(net409),
    .X(_00677_));
 sg13g2_mux2_1 _20034_ (.A0(net850),
    .A1(\cpu.dcache.r_tag[4][9] ),
    .S(_02948_),
    .X(_00678_));
 sg13g2_mux2_1 _20035_ (.A0(net849),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(_02948_),
    .X(_00679_));
 sg13g2_mux2_1 _20036_ (.A0(net848),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(net409),
    .X(_00680_));
 sg13g2_mux2_1 _20037_ (.A0(net344),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net409),
    .X(_00681_));
 sg13g2_mux2_1 _20038_ (.A0(net376),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net409),
    .X(_00682_));
 sg13g2_mux2_1 _20039_ (.A0(net436),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(net409),
    .X(_00683_));
 sg13g2_inv_1 _20040_ (.Y(_02951_),
    .A(\cpu.dcache.r_tag[5][5] ));
 sg13g2_buf_1 _20041_ (.A(net481),
    .X(_02952_));
 sg13g2_buf_1 _20042_ (.A(_12491_),
    .X(_02953_));
 sg13g2_nand2_1 _20043_ (.Y(_02954_),
    .A(net643),
    .B(net471));
 sg13g2_o21ai_1 _20044_ (.B1(_02954_),
    .Y(_00684_),
    .A1(_02951_),
    .A2(net408));
 sg13g2_mux2_1 _20045_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net438),
    .S(net408),
    .X(_00685_));
 sg13g2_mux2_1 _20046_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(net435),
    .S(net408),
    .X(_00686_));
 sg13g2_mux2_1 _20047_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(net432),
    .S(net408),
    .X(_00687_));
 sg13g2_mux2_1 _20048_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net439),
    .S(net408),
    .X(_00688_));
 sg13g2_mux2_1 _20049_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net433),
    .S(net408),
    .X(_00689_));
 sg13g2_mux2_1 _20050_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net430),
    .S(_02952_),
    .X(_00690_));
 sg13g2_mux2_1 _20051_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(net434),
    .S(net408),
    .X(_00691_));
 sg13g2_mux2_1 _20052_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net431),
    .S(net408),
    .X(_00692_));
 sg13g2_mux2_1 _20053_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(net437),
    .S(_02952_),
    .X(_00693_));
 sg13g2_mux2_1 _20054_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(net722),
    .S(net471),
    .X(_00694_));
 sg13g2_mux2_1 _20055_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(net721),
    .S(net471),
    .X(_00695_));
 sg13g2_mux2_1 _20056_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(net720),
    .S(_02953_),
    .X(_00696_));
 sg13g2_mux2_1 _20057_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(net844),
    .S(net471),
    .X(_00697_));
 sg13g2_mux2_1 _20058_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(net843),
    .S(net471),
    .X(_00698_));
 sg13g2_mux2_1 _20059_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(net842),
    .S(_02953_),
    .X(_00699_));
 sg13g2_mux2_1 _20060_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net344),
    .S(net471),
    .X(_00700_));
 sg13g2_mux2_1 _20061_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net376),
    .S(net471),
    .X(_00701_));
 sg13g2_mux2_1 _20062_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net436),
    .S(net471),
    .X(_00702_));
 sg13g2_buf_1 _20063_ (.A(net418),
    .X(_02955_));
 sg13g2_mux2_1 _20064_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net596),
    .S(_02955_),
    .X(_00703_));
 sg13g2_mux2_1 _20065_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(_09444_),
    .S(net369),
    .X(_00704_));
 sg13g2_mux2_1 _20066_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(_09515_),
    .S(net369),
    .X(_00705_));
 sg13g2_mux2_1 _20067_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(net432),
    .S(net369),
    .X(_00706_));
 sg13g2_mux2_1 _20068_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(_09342_),
    .S(_02955_),
    .X(_00707_));
 sg13g2_mux2_1 _20069_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(_09562_),
    .S(net369),
    .X(_00708_));
 sg13g2_mux2_1 _20070_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(net430),
    .S(net369),
    .X(_00709_));
 sg13g2_mux2_1 _20071_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net434),
    .S(net369),
    .X(_00710_));
 sg13g2_mux2_1 _20072_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(net431),
    .S(net369),
    .X(_00711_));
 sg13g2_buf_1 _20073_ (.A(_02707_),
    .X(_02956_));
 sg13g2_mux2_1 _20074_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(net437),
    .S(net407),
    .X(_00712_));
 sg13g2_mux2_1 _20075_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(net722),
    .S(net407),
    .X(_00713_));
 sg13g2_mux2_1 _20076_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net721),
    .S(net407),
    .X(_00714_));
 sg13g2_mux2_1 _20077_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net720),
    .S(net407),
    .X(_00715_));
 sg13g2_mux2_1 _20078_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(net844),
    .S(_02956_),
    .X(_00716_));
 sg13g2_inv_1 _20079_ (.Y(_02957_),
    .A(\cpu.dcache.r_tag[6][10] ));
 sg13g2_nand2_1 _20080_ (.Y(_02958_),
    .A(net951),
    .B(_02956_));
 sg13g2_o21ai_1 _20081_ (.B1(_02958_),
    .Y(_00717_),
    .A1(_02957_),
    .A2(net369));
 sg13g2_mux2_1 _20082_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(net842),
    .S(net407),
    .X(_00718_));
 sg13g2_mux2_1 _20083_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(_09249_),
    .S(net407),
    .X(_00719_));
 sg13g2_mux2_1 _20084_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(_09316_),
    .S(net407),
    .X(_00720_));
 sg13g2_mux2_1 _20085_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net436),
    .S(net407),
    .X(_00721_));
 sg13g2_buf_1 _20086_ (.A(net417),
    .X(_02959_));
 sg13g2_mux2_1 _20087_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net596),
    .S(net368),
    .X(_00722_));
 sg13g2_mux2_1 _20088_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(_09444_),
    .S(net368),
    .X(_00723_));
 sg13g2_mux2_1 _20089_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(_09515_),
    .S(net368),
    .X(_00724_));
 sg13g2_mux2_1 _20090_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(_09586_),
    .S(_02959_),
    .X(_00725_));
 sg13g2_mux2_1 _20091_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(_09342_),
    .S(net368),
    .X(_00726_));
 sg13g2_mux2_1 _20092_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net433),
    .S(net368),
    .X(_00727_));
 sg13g2_mux2_1 _20093_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net430),
    .S(net368),
    .X(_00728_));
 sg13g2_mux2_1 _20094_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(net434),
    .S(net368),
    .X(_00729_));
 sg13g2_mux2_1 _20095_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(_09609_),
    .S(net368),
    .X(_00730_));
 sg13g2_mux2_1 _20096_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09467_),
    .S(_02959_),
    .X(_00731_));
 sg13g2_buf_1 _20097_ (.A(net417),
    .X(_02960_));
 sg13g2_mux2_1 _20098_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net722),
    .S(net367),
    .X(_00732_));
 sg13g2_mux2_1 _20099_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net721),
    .S(net367),
    .X(_00733_));
 sg13g2_mux2_1 _20100_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net720),
    .S(_02960_),
    .X(_00734_));
 sg13g2_mux2_1 _20101_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net844),
    .S(net367),
    .X(_00735_));
 sg13g2_mux2_1 _20102_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net843),
    .S(_02960_),
    .X(_00736_));
 sg13g2_mux2_1 _20103_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(net842),
    .S(net367),
    .X(_00737_));
 sg13g2_mux2_1 _20104_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(_09249_),
    .S(net367),
    .X(_00738_));
 sg13g2_mux2_1 _20105_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net376),
    .S(net367),
    .X(_00739_));
 sg13g2_mux2_1 _20106_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(net436),
    .S(net367),
    .X(_00740_));
 sg13g2_nor2_1 _20107_ (.A(_08223_),
    .B(_08922_),
    .Y(_02961_));
 sg13g2_buf_1 _20108_ (.A(_02961_),
    .X(_02962_));
 sg13g2_buf_1 _20109_ (.A(_09718_),
    .X(_02963_));
 sg13g2_buf_1 _20110_ (.A(_08307_),
    .X(_02964_));
 sg13g2_nor2_1 _20111_ (.A(_08292_),
    .B(net241),
    .Y(_02965_));
 sg13g2_buf_2 _20112_ (.A(_02965_),
    .X(_02966_));
 sg13g2_buf_1 _20113_ (.A(_08293_),
    .X(_02967_));
 sg13g2_nor2_1 _20114_ (.A(_08882_),
    .B(net240),
    .Y(_02968_));
 sg13g2_buf_1 _20115_ (.A(_02968_),
    .X(_02969_));
 sg13g2_a21oi_1 _20116_ (.A1(_08248_),
    .A2(_02966_),
    .Y(_02970_),
    .B1(_02969_));
 sg13g2_nor2_1 _20117_ (.A(net161),
    .B(_02970_),
    .Y(_02971_));
 sg13g2_a21oi_1 _20118_ (.A1(net147),
    .A2(net146),
    .Y(_02972_),
    .B1(_02971_));
 sg13g2_nand2_1 _20119_ (.Y(_02973_),
    .A(_10176_),
    .B(net91));
 sg13g2_o21ai_1 _20120_ (.B1(_02973_),
    .Y(_00749_),
    .A1(_09762_),
    .A2(_02972_));
 sg13g2_buf_1 _20121_ (.A(net241),
    .X(_02974_));
 sg13g2_buf_1 _20122_ (.A(net161),
    .X(_02975_));
 sg13g2_buf_1 _20123_ (.A(_08922_),
    .X(_02976_));
 sg13g2_nand2_1 _20124_ (.Y(_02977_),
    .A(net160),
    .B(net240));
 sg13g2_a21oi_1 _20125_ (.A1(net145),
    .A2(_02977_),
    .Y(_02978_),
    .B1(_02969_));
 sg13g2_buf_1 _20126_ (.A(_08292_),
    .X(_02979_));
 sg13g2_nor2_1 _20127_ (.A(_08223_),
    .B(net315),
    .Y(_02980_));
 sg13g2_buf_1 _20128_ (.A(_08882_),
    .X(_02981_));
 sg13g2_nand2_1 _20129_ (.Y(_02982_),
    .A(net164),
    .B(net206));
 sg13g2_nand2_1 _20130_ (.Y(_02983_),
    .A(_08884_),
    .B(_02982_));
 sg13g2_a22oi_1 _20131_ (.Y(_02984_),
    .B1(_02983_),
    .B2(net166),
    .A2(_02980_),
    .A1(net165));
 sg13g2_o21ai_1 _20132_ (.B1(_02984_),
    .Y(_02985_),
    .A1(net207),
    .A2(_02978_));
 sg13g2_nor2_1 _20133_ (.A(_09762_),
    .B(_02985_),
    .Y(_02986_));
 sg13g2_a21oi_1 _20134_ (.A1(net1033),
    .A2(net91),
    .Y(_00750_),
    .B1(_02986_));
 sg13g2_buf_1 _20135_ (.A(_08924_),
    .X(_02987_));
 sg13g2_buf_1 _20136_ (.A(_08271_),
    .X(_02988_));
 sg13g2_nand2_1 _20137_ (.Y(_02989_),
    .A(net239),
    .B(net315));
 sg13g2_nor3_1 _20138_ (.A(net109),
    .B(net121),
    .C(_02989_),
    .Y(_02990_));
 sg13g2_a21o_1 _20139_ (.A2(net111),
    .A1(\cpu.cond[1] ),
    .B1(_02990_),
    .X(_00751_));
 sg13g2_buf_1 _20140_ (.A(net315),
    .X(_02991_));
 sg13g2_buf_1 _20141_ (.A(_02976_),
    .X(_02992_));
 sg13g2_a21oi_1 _20142_ (.A1(_02991_),
    .A2(_02982_),
    .Y(_02993_),
    .B1(net144));
 sg13g2_mux2_1 _20143_ (.A0(_02993_),
    .A1(\cpu.cond[2] ),
    .S(net106),
    .X(_00752_));
 sg13g2_nand3_1 _20144_ (.B(_08925_),
    .C(_08992_),
    .A(_08919_),
    .Y(_02994_));
 sg13g2_nand2_1 _20145_ (.Y(_02995_),
    .A(_09202_),
    .B(_08997_));
 sg13g2_o21ai_1 _20146_ (.B1(_02995_),
    .Y(_00753_),
    .A1(_08928_),
    .A2(_02994_));
 sg13g2_nand2_1 _20147_ (.Y(_02996_),
    .A(net206),
    .B(_08309_));
 sg13g2_buf_2 _20148_ (.A(_02996_),
    .X(_02997_));
 sg13g2_nand2_1 _20149_ (.Y(_02998_),
    .A(\cpu.icache.r_data[7][8] ),
    .B(_08178_));
 sg13g2_a22oi_1 _20150_ (.Y(_02999_),
    .B1(net499),
    .B2(\cpu.icache.r_data[1][8] ),
    .A2(net447),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_a22oi_1 _20151_ (.Y(_03000_),
    .B1(_08201_),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(net622),
    .A1(\cpu.icache.r_data[4][8] ));
 sg13g2_a22oi_1 _20152_ (.Y(_03001_),
    .B1(net502),
    .B2(\cpu.icache.r_data[5][8] ),
    .A2(net621),
    .A1(\cpu.icache.r_data[6][8] ));
 sg13g2_nand4_1 _20153_ (.B(_02999_),
    .C(_03000_),
    .A(_02998_),
    .Y(_03002_),
    .D(_03001_));
 sg13g2_nand2_1 _20154_ (.Y(_03003_),
    .A(_00174_),
    .B(net452));
 sg13g2_o21ai_1 _20155_ (.B1(_03003_),
    .Y(_03004_),
    .A1(_08158_),
    .A2(_03002_));
 sg13g2_nor2_1 _20156_ (.A(_00175_),
    .B(net387),
    .Y(_03005_));
 sg13g2_mux2_1 _20157_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(net799),
    .X(_03006_));
 sg13g2_a22oi_1 _20158_ (.Y(_03007_),
    .B1(_03006_),
    .B2(_08320_),
    .A2(net689),
    .A1(\cpu.icache.r_data[5][24] ));
 sg13g2_nor2_1 _20159_ (.A(_08226_),
    .B(_03007_),
    .Y(_03008_));
 sg13g2_a22oi_1 _20160_ (.Y(_03009_),
    .B1(_08166_),
    .B2(\cpu.icache.r_data[1][24] ),
    .A2(_08173_),
    .A1(\cpu.icache.r_data[2][24] ));
 sg13g2_a22oi_1 _20161_ (.Y(_03010_),
    .B1(net503),
    .B2(\cpu.icache.r_data[7][24] ),
    .A2(net450),
    .A1(\cpu.icache.r_data[3][24] ));
 sg13g2_nand2_1 _20162_ (.Y(_03011_),
    .A(_03009_),
    .B(_03010_));
 sg13g2_nor4_1 _20163_ (.A(net913),
    .B(_03005_),
    .C(_03008_),
    .D(_03011_),
    .Y(_03012_));
 sg13g2_a21oi_1 _20164_ (.A1(net913),
    .A2(_03004_),
    .Y(_03013_),
    .B1(_03012_));
 sg13g2_buf_1 _20165_ (.A(_03013_),
    .X(_03014_));
 sg13g2_nand2_1 _20166_ (.Y(_03015_),
    .A(\cpu.icache.r_data[7][9] ),
    .B(_08177_));
 sg13g2_a22oi_1 _20167_ (.Y(_03016_),
    .B1(_08165_),
    .B2(\cpu.icache.r_data[1][9] ),
    .A2(_08172_),
    .A1(\cpu.icache.r_data[2][9] ));
 sg13g2_a22oi_1 _20168_ (.Y(_03017_),
    .B1(net501),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(net622),
    .A1(\cpu.icache.r_data[4][9] ));
 sg13g2_a22oi_1 _20169_ (.Y(_03018_),
    .B1(net502),
    .B2(\cpu.icache.r_data[5][9] ),
    .A2(net621),
    .A1(\cpu.icache.r_data[6][9] ));
 sg13g2_nand4_1 _20170_ (.B(_03016_),
    .C(_03017_),
    .A(_03015_),
    .Y(_03019_),
    .D(_03018_));
 sg13g2_nand2_1 _20171_ (.Y(_03020_),
    .A(_00176_),
    .B(net506));
 sg13g2_o21ai_1 _20172_ (.B1(_03020_),
    .Y(_03021_),
    .A1(net452),
    .A2(_03019_));
 sg13g2_nor2_1 _20173_ (.A(_00177_),
    .B(_08211_),
    .Y(_03022_));
 sg13g2_mux2_1 _20174_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(net799),
    .X(_03023_));
 sg13g2_a22oi_1 _20175_ (.Y(_03024_),
    .B1(_03023_),
    .B2(_08320_),
    .A2(_08196_),
    .A1(\cpu.icache.r_data[7][25] ));
 sg13g2_nor2_1 _20176_ (.A(net691),
    .B(_03024_),
    .Y(_03025_));
 sg13g2_a22oi_1 _20177_ (.Y(_03026_),
    .B1(net502),
    .B2(\cpu.icache.r_data[5][25] ),
    .A2(_08217_),
    .A1(\cpu.icache.r_data[1][25] ));
 sg13g2_a22oi_1 _20178_ (.Y(_03027_),
    .B1(_08200_),
    .B2(\cpu.icache.r_data[3][25] ),
    .A2(_08214_),
    .A1(\cpu.icache.r_data[2][25] ));
 sg13g2_nand2_1 _20179_ (.Y(_03028_),
    .A(_03026_),
    .B(_03027_));
 sg13g2_nor4_1 _20180_ (.A(_08312_),
    .B(_03022_),
    .C(_03025_),
    .D(_03028_),
    .Y(_03029_));
 sg13g2_a21oi_1 _20181_ (.A1(_08312_),
    .A2(_03021_),
    .Y(_03030_),
    .B1(_03029_));
 sg13g2_buf_1 _20182_ (.A(_03030_),
    .X(_03031_));
 sg13g2_nand2_1 _20183_ (.Y(_03032_),
    .A(\cpu.icache.r_data[4][7] ),
    .B(_08183_));
 sg13g2_a22oi_1 _20184_ (.Y(_03033_),
    .B1(_08177_),
    .B2(\cpu.icache.r_data[7][7] ),
    .A2(_08172_),
    .A1(\cpu.icache.r_data[2][7] ));
 sg13g2_a22oi_1 _20185_ (.Y(_03034_),
    .B1(_08264_),
    .B2(\cpu.icache.r_data[3][7] ),
    .A2(_08185_),
    .A1(\cpu.icache.r_data[5][7] ));
 sg13g2_nand2b_1 _20186_ (.Y(_03035_),
    .B(_08233_),
    .A_N(_03034_));
 sg13g2_a22oi_1 _20187_ (.Y(_03036_),
    .B1(net499),
    .B2(\cpu.icache.r_data[1][7] ),
    .A2(_08195_),
    .A1(\cpu.icache.r_data[6][7] ));
 sg13g2_nand4_1 _20188_ (.B(_03033_),
    .C(_03035_),
    .A(_03032_),
    .Y(_03037_),
    .D(_03036_));
 sg13g2_nand2_1 _20189_ (.Y(_03038_),
    .A(_00172_),
    .B(net452));
 sg13g2_o21ai_1 _20190_ (.B1(_03038_),
    .Y(_03039_),
    .A1(net452),
    .A2(_03037_));
 sg13g2_nand2_1 _20191_ (.Y(_03040_),
    .A(\cpu.icache.r_data[7][23] ),
    .B(_08178_));
 sg13g2_a22oi_1 _20192_ (.Y(_03041_),
    .B1(_08217_),
    .B2(\cpu.icache.r_data[1][23] ),
    .A2(_08195_),
    .A1(\cpu.icache.r_data[6][23] ));
 sg13g2_a22oi_1 _20193_ (.Y(_03042_),
    .B1(net447),
    .B2(\cpu.icache.r_data[2][23] ),
    .A2(_08183_),
    .A1(\cpu.icache.r_data[4][23] ));
 sg13g2_a22oi_1 _20194_ (.Y(_03043_),
    .B1(_08189_),
    .B2(\cpu.icache.r_data[5][23] ),
    .A2(_08200_),
    .A1(\cpu.icache.r_data[3][23] ));
 sg13g2_nand4_1 _20195_ (.B(_03041_),
    .C(_03042_),
    .A(_03040_),
    .Y(_03044_),
    .D(_03043_));
 sg13g2_nor2_1 _20196_ (.A(_00173_),
    .B(_08212_),
    .Y(_03045_));
 sg13g2_o21ai_1 _20197_ (.B1(_08142_),
    .Y(_03046_),
    .A1(_03044_),
    .A2(_03045_));
 sg13g2_o21ai_1 _20198_ (.B1(_03046_),
    .Y(_03047_),
    .A1(net1060),
    .A2(_03039_));
 sg13g2_buf_1 _20199_ (.A(_03047_),
    .X(_03048_));
 sg13g2_nor3_1 _20200_ (.A(net205),
    .B(net204),
    .C(_03048_),
    .Y(_03049_));
 sg13g2_nand2_1 _20201_ (.Y(_03050_),
    .A(_09712_),
    .B(_03049_));
 sg13g2_nor3_1 _20202_ (.A(_02987_),
    .B(_02997_),
    .C(_03050_),
    .Y(_03051_));
 sg13g2_nand3_1 _20203_ (.B(_08992_),
    .C(_03051_),
    .A(_08947_),
    .Y(_03052_));
 sg13g2_nand2_1 _20204_ (.Y(_03053_),
    .A(\cpu.dec.do_flush_all ),
    .B(net108));
 sg13g2_o21ai_1 _20205_ (.B1(_03053_),
    .Y(_00754_),
    .A1(net92),
    .A2(_03052_));
 sg13g2_nand2_1 _20206_ (.Y(_03054_),
    .A(net239),
    .B(_02966_));
 sg13g2_nor3_1 _20207_ (.A(_08893_),
    .B(net121),
    .C(_03054_),
    .Y(_03055_));
 sg13g2_a21o_1 _20208_ (.A2(net111),
    .A1(\cpu.dec.do_flush_write ),
    .B1(_03055_),
    .X(_00755_));
 sg13g2_nor2_1 _20209_ (.A(_08924_),
    .B(_02997_),
    .Y(_03056_));
 sg13g2_buf_1 _20210_ (.A(_08880_),
    .X(_03057_));
 sg13g2_nor2_1 _20211_ (.A(_09718_),
    .B(_08922_),
    .Y(_03058_));
 sg13g2_mux2_1 _20212_ (.A0(_03058_),
    .A1(net240),
    .S(net239),
    .X(_03059_));
 sg13g2_a21oi_1 _20213_ (.A1(_02974_),
    .A2(_03059_),
    .Y(_03060_),
    .B1(_02980_));
 sg13g2_nor2_1 _20214_ (.A(net237),
    .B(_03060_),
    .Y(_03061_));
 sg13g2_a21oi_1 _20215_ (.A1(net343),
    .A2(_03056_),
    .Y(_03062_),
    .B1(_03061_));
 sg13g2_buf_1 _20216_ (.A(_08946_),
    .X(_03063_));
 sg13g2_nand2_1 _20217_ (.Y(_03064_),
    .A(net160),
    .B(net203));
 sg13g2_o21ai_1 _20218_ (.B1(_03064_),
    .Y(_03065_),
    .A1(net160),
    .A2(_03057_));
 sg13g2_nor2_1 _20219_ (.A(_02967_),
    .B(_08307_),
    .Y(_03066_));
 sg13g2_nand3_1 _20220_ (.B(_03065_),
    .C(_03066_),
    .A(net145),
    .Y(_03067_));
 sg13g2_o21ai_1 _20221_ (.B1(_03067_),
    .Y(_03068_),
    .A1(_02962_),
    .A2(_03062_));
 sg13g2_mux2_1 _20222_ (.A0(_03068_),
    .A1(_10921_),
    .S(net106),
    .X(_00756_));
 sg13g2_inv_1 _20223_ (.Y(_03069_),
    .A(\cpu.dec.imm[10] ));
 sg13g2_buf_1 _20224_ (.A(net109),
    .X(_03070_));
 sg13g2_nand2_1 _20225_ (.Y(_03071_),
    .A(net206),
    .B(net241));
 sg13g2_buf_2 _20226_ (.A(_03071_),
    .X(_03072_));
 sg13g2_o21ai_1 _20227_ (.B1(_03058_),
    .Y(_03073_),
    .A1(net203),
    .A2(_03072_));
 sg13g2_buf_1 _20228_ (.A(_03073_),
    .X(_03074_));
 sg13g2_inv_1 _20229_ (.Y(_03075_),
    .A(_03074_));
 sg13g2_or2_1 _20230_ (.X(_03076_),
    .B(_08307_),
    .A(_08292_));
 sg13g2_buf_2 _20231_ (.A(_03076_),
    .X(_03077_));
 sg13g2_inv_1 _20232_ (.Y(_03078_),
    .A(net205));
 sg13g2_nand2b_1 _20233_ (.Y(_03079_),
    .B(_08292_),
    .A_N(_08307_));
 sg13g2_nor2_1 _20234_ (.A(net239),
    .B(_03079_),
    .Y(_03080_));
 sg13g2_buf_1 _20235_ (.A(_03080_),
    .X(_03081_));
 sg13g2_nand2_1 _20236_ (.Y(_03082_),
    .A(net190),
    .B(_02969_));
 sg13g2_buf_2 _20237_ (.A(_03082_),
    .X(_03083_));
 sg13g2_nand2_1 _20238_ (.Y(_03084_),
    .A(_03072_),
    .B(_03083_));
 sg13g2_a21oi_1 _20239_ (.A1(net203),
    .A2(_03081_),
    .Y(_03085_),
    .B1(_03084_));
 sg13g2_o21ai_1 _20240_ (.B1(_03085_),
    .Y(_03086_),
    .A1(_03077_),
    .A2(_03078_));
 sg13g2_nor2_1 _20241_ (.A(_08924_),
    .B(_09741_),
    .Y(_03087_));
 sg13g2_buf_2 _20242_ (.A(_03087_),
    .X(_03088_));
 sg13g2_inv_1 _20243_ (.Y(_03089_),
    .A(_08946_));
 sg13g2_nand2_1 _20244_ (.Y(_03090_),
    .A(net206),
    .B(_03066_));
 sg13g2_buf_2 _20245_ (.A(_03090_),
    .X(_03091_));
 sg13g2_o21ai_1 _20246_ (.B1(_03083_),
    .Y(_03092_),
    .A1(_03089_),
    .A2(_03091_));
 sg13g2_a22oi_1 _20247_ (.Y(_03093_),
    .B1(_03088_),
    .B2(_03092_),
    .A2(_03086_),
    .A1(_03075_));
 sg13g2_nor2_1 _20248_ (.A(_08271_),
    .B(_03077_),
    .Y(_03094_));
 sg13g2_buf_1 _20249_ (.A(_03094_),
    .X(_03095_));
 sg13g2_nand2_1 _20250_ (.Y(_03096_),
    .A(_08922_),
    .B(_03095_));
 sg13g2_o21ai_1 _20251_ (.B1(_03096_),
    .Y(_03097_),
    .A1(_08922_),
    .A2(_08311_));
 sg13g2_nand3_1 _20252_ (.B(_03063_),
    .C(_03097_),
    .A(net161),
    .Y(_03098_));
 sg13g2_nor2b_1 _20253_ (.A(_09761_),
    .B_N(_03098_),
    .Y(_03099_));
 sg13g2_buf_2 _20254_ (.A(_03099_),
    .X(_03100_));
 sg13g2_a22oi_1 _20255_ (.Y(_00757_),
    .B1(_03093_),
    .B2(_03100_),
    .A2(net86),
    .A1(_03069_));
 sg13g2_inv_1 _20256_ (.Y(_03101_),
    .A(\cpu.dec.imm[11] ));
 sg13g2_o21ai_1 _20257_ (.B1(_03083_),
    .Y(_03102_),
    .A1(net237),
    .A2(_03091_));
 sg13g2_nor2_1 _20258_ (.A(_08271_),
    .B(_02967_),
    .Y(_03103_));
 sg13g2_buf_2 _20259_ (.A(_03103_),
    .X(_03104_));
 sg13g2_nor2_1 _20260_ (.A(_08917_),
    .B(_03104_),
    .Y(_03105_));
 sg13g2_o21ai_1 _20261_ (.B1(net239),
    .Y(_03106_),
    .A1(_08309_),
    .A2(_08917_));
 sg13g2_o21ai_1 _20262_ (.B1(_03106_),
    .Y(_03107_),
    .A1(net241),
    .A2(_03105_));
 sg13g2_buf_1 _20263_ (.A(_03107_),
    .X(_03108_));
 sg13g2_or3_1 _20264_ (.A(_08334_),
    .B(_03031_),
    .C(_03048_),
    .X(_03109_));
 sg13g2_nor2_1 _20265_ (.A(_03078_),
    .B(_03109_),
    .Y(_03110_));
 sg13g2_buf_1 _20266_ (.A(_03110_),
    .X(_03111_));
 sg13g2_a21oi_1 _20267_ (.A1(_03089_),
    .A2(net143),
    .Y(_03112_),
    .B1(_03091_));
 sg13g2_buf_1 _20268_ (.A(_03112_),
    .X(_03113_));
 sg13g2_o21ai_1 _20269_ (.B1(_03113_),
    .Y(_03114_),
    .A1(_08919_),
    .A2(net143));
 sg13g2_nand2_1 _20270_ (.Y(_03115_),
    .A(_03108_),
    .B(_03114_));
 sg13g2_a22oi_1 _20271_ (.Y(_03116_),
    .B1(_03115_),
    .B2(_03075_),
    .A2(_03102_),
    .A1(_03088_));
 sg13g2_a22oi_1 _20272_ (.Y(_00758_),
    .B1(_03100_),
    .B2(_03116_),
    .A2(net86),
    .A1(_03101_));
 sg13g2_inv_1 _20273_ (.Y(_03117_),
    .A(\cpu.dec.imm[12] ));
 sg13g2_nand2_1 _20274_ (.Y(_03118_),
    .A(net249),
    .B(_03081_));
 sg13g2_nand2_1 _20275_ (.Y(_03119_),
    .A(_03083_),
    .B(_03118_));
 sg13g2_o21ai_1 _20276_ (.B1(_03113_),
    .Y(_03120_),
    .A1(net249),
    .A2(net143));
 sg13g2_nand2_1 _20277_ (.Y(_03121_),
    .A(_03108_),
    .B(_03120_));
 sg13g2_a22oi_1 _20278_ (.Y(_03122_),
    .B1(_03121_),
    .B2(_03075_),
    .A2(_03119_),
    .A1(_03088_));
 sg13g2_a22oi_1 _20279_ (.Y(_00759_),
    .B1(_03100_),
    .B2(_03122_),
    .A2(net86),
    .A1(_03117_));
 sg13g2_and3_1 _20280_ (.X(_03123_),
    .A(net238),
    .B(net165),
    .C(_03072_));
 sg13g2_o21ai_1 _20281_ (.B1(_03113_),
    .Y(_03124_),
    .A1(net165),
    .A2(net143));
 sg13g2_nand2_1 _20282_ (.Y(_03125_),
    .A(_03108_),
    .B(_03124_));
 sg13g2_a22oi_1 _20283_ (.Y(_03126_),
    .B1(_03125_),
    .B2(_03075_),
    .A2(_03123_),
    .A1(_09720_));
 sg13g2_a22oi_1 _20284_ (.Y(_00760_),
    .B1(_03100_),
    .B2(_03126_),
    .A2(net86),
    .A1(_11240_));
 sg13g2_inv_1 _20285_ (.Y(_03127_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_o21ai_1 _20286_ (.B1(_03083_),
    .Y(_03128_),
    .A1(_08887_),
    .A2(_03091_));
 sg13g2_nand2_1 _20287_ (.Y(_03129_),
    .A(_03088_),
    .B(_03128_));
 sg13g2_o21ai_1 _20288_ (.B1(_03113_),
    .Y(_03130_),
    .A1(net191),
    .A2(net143));
 sg13g2_a21oi_1 _20289_ (.A1(_03108_),
    .A2(_03130_),
    .Y(_03131_),
    .B1(_03074_));
 sg13g2_nor2b_1 _20290_ (.A(_03131_),
    .B_N(_03100_),
    .Y(_03132_));
 sg13g2_a22oi_1 _20291_ (.Y(_00761_),
    .B1(_03129_),
    .B2(_03132_),
    .A2(net86),
    .A1(_03127_));
 sg13g2_inv_1 _20292_ (.Y(_03133_),
    .A(\cpu.dec.imm[15] ));
 sg13g2_o21ai_1 _20293_ (.B1(_03083_),
    .Y(_03134_),
    .A1(net191),
    .A2(_03091_));
 sg13g2_nand2_1 _20294_ (.Y(_03135_),
    .A(_03088_),
    .B(_03134_));
 sg13g2_a22oi_1 _20295_ (.Y(_00762_),
    .B1(_03132_),
    .B2(_03135_),
    .A2(net86),
    .A1(_03133_));
 sg13g2_or2_1 _20296_ (.X(_03136_),
    .B(_03056_),
    .A(_02971_));
 sg13g2_buf_1 _20297_ (.A(_02988_),
    .X(_03137_));
 sg13g2_nand2_1 _20298_ (.Y(_03138_),
    .A(_02979_),
    .B(_02964_));
 sg13g2_o21ai_1 _20299_ (.B1(_03138_),
    .Y(_03139_),
    .A1(net166),
    .A2(_03077_));
 sg13g2_a21oi_1 _20300_ (.A1(_02979_),
    .A2(_03111_),
    .Y(_03140_),
    .B1(_02964_));
 sg13g2_or2_1 _20301_ (.X(_03141_),
    .B(_03140_),
    .A(net160));
 sg13g2_nor2b_1 _20302_ (.A(_03139_),
    .B_N(_03141_),
    .Y(_03142_));
 sg13g2_nor2_1 _20303_ (.A(_02963_),
    .B(net147),
    .Y(_03143_));
 sg13g2_o21ai_1 _20304_ (.B1(_03143_),
    .Y(_03144_),
    .A1(net202),
    .A2(_03142_));
 sg13g2_a22oi_1 _20305_ (.Y(_03145_),
    .B1(_03144_),
    .B2(net249),
    .A2(_03136_),
    .A1(net346));
 sg13g2_nand2_1 _20306_ (.Y(_03146_),
    .A(_10888_),
    .B(net108));
 sg13g2_o21ai_1 _20307_ (.B1(_03146_),
    .Y(_00763_),
    .A1(net92),
    .A2(_03145_));
 sg13g2_nand2_1 _20308_ (.Y(_03147_),
    .A(_08223_),
    .B(_03072_));
 sg13g2_nand2_1 _20309_ (.Y(_03148_),
    .A(_03081_),
    .B(net143));
 sg13g2_nand2_1 _20310_ (.Y(_03149_),
    .A(net147),
    .B(net346));
 sg13g2_o21ai_1 _20311_ (.B1(_03149_),
    .Y(_03150_),
    .A1(net237),
    .A2(_03148_));
 sg13g2_a21oi_1 _20312_ (.A1(_08335_),
    .A2(_03147_),
    .Y(_03151_),
    .B1(_02992_));
 sg13g2_o21ai_1 _20313_ (.B1(_03151_),
    .Y(_03152_),
    .A1(_03147_),
    .A2(_03150_));
 sg13g2_nand2_1 _20314_ (.Y(_03153_),
    .A(_09718_),
    .B(_08922_));
 sg13g2_buf_2 _20315_ (.A(_03153_),
    .X(_03154_));
 sg13g2_a221oi_1 _20316_ (.B2(_08335_),
    .C1(_03154_),
    .B1(_03095_),
    .A1(net238),
    .Y(_03155_),
    .A2(net237));
 sg13g2_nor2_1 _20317_ (.A(net238),
    .B(_03095_),
    .Y(_03156_));
 sg13g2_nand2_1 _20318_ (.Y(_03157_),
    .A(_09723_),
    .B(_03156_));
 sg13g2_a21oi_1 _20319_ (.A1(_03077_),
    .A2(_03138_),
    .Y(_03158_),
    .B1(_02988_));
 sg13g2_nand2_1 _20320_ (.Y(_03159_),
    .A(net189),
    .B(_03158_));
 sg13g2_a21oi_1 _20321_ (.A1(_03149_),
    .A2(_03159_),
    .Y(_03160_),
    .B1(net121));
 sg13g2_a221oi_1 _20322_ (.B2(_03157_),
    .C1(_03160_),
    .B1(_03155_),
    .A1(net203),
    .Y(_03161_),
    .A2(_03136_));
 sg13g2_nand2_1 _20323_ (.Y(_03162_),
    .A(_03152_),
    .B(_03161_));
 sg13g2_mux2_1 _20324_ (.A0(_03162_),
    .A1(_10811_),
    .S(net106),
    .X(_00764_));
 sg13g2_inv_1 _20325_ (.Y(_03163_),
    .A(_03148_));
 sg13g2_a22oi_1 _20326_ (.Y(_03164_),
    .B1(_02969_),
    .B2(net189),
    .A2(_03063_),
    .A1(_08886_));
 sg13g2_o21ai_1 _20327_ (.B1(_03164_),
    .Y(_03165_),
    .A1(_03057_),
    .A2(_03077_));
 sg13g2_a21oi_1 _20328_ (.A1(net191),
    .A2(_03163_),
    .Y(_03166_),
    .B1(_03165_));
 sg13g2_nand2_1 _20329_ (.Y(_03167_),
    .A(_03058_),
    .B(_03072_));
 sg13g2_o21ai_1 _20330_ (.B1(_03164_),
    .Y(_03168_),
    .A1(net237),
    .A2(_02997_));
 sg13g2_nor2_1 _20331_ (.A(_03089_),
    .B(_03154_),
    .Y(_03169_));
 sg13g2_a22oi_1 _20332_ (.Y(_03170_),
    .B1(_03147_),
    .B2(_02977_),
    .A2(_03095_),
    .A1(net160));
 sg13g2_nor2_1 _20333_ (.A(_08887_),
    .B(_03170_),
    .Y(_03171_));
 sg13g2_a221oi_1 _20334_ (.B2(_03156_),
    .C1(_03171_),
    .B1(_03169_),
    .A1(_09720_),
    .Y(_03172_),
    .A2(_03168_));
 sg13g2_o21ai_1 _20335_ (.B1(_03172_),
    .Y(_03173_),
    .A1(_03166_),
    .A2(_03167_));
 sg13g2_mux2_1 _20336_ (.A0(_03173_),
    .A1(_10852_),
    .S(_09768_),
    .X(_00765_));
 sg13g2_o21ai_1 _20337_ (.B1(_03143_),
    .Y(_03174_),
    .A1(_03137_),
    .A2(_03141_));
 sg13g2_a22oi_1 _20338_ (.Y(_03175_),
    .B1(_03174_),
    .B2(net165),
    .A2(_02971_),
    .A1(net191));
 sg13g2_nand2_1 _20339_ (.Y(_03176_),
    .A(\cpu.dec.imm[4] ),
    .B(net108));
 sg13g2_o21ai_1 _20340_ (.B1(_03176_),
    .Y(_00766_),
    .A1(net92),
    .A2(_03175_));
 sg13g2_nor2_1 _20341_ (.A(net161),
    .B(net240),
    .Y(_03177_));
 sg13g2_o21ai_1 _20342_ (.B1(net202),
    .Y(_03178_),
    .A1(_08309_),
    .A2(_03177_));
 sg13g2_o21ai_1 _20343_ (.B1(_03058_),
    .Y(_03179_),
    .A1(_03079_),
    .A2(_03111_));
 sg13g2_nand3_1 _20344_ (.B(_03178_),
    .C(_03179_),
    .A(_03154_),
    .Y(_03180_));
 sg13g2_nor2_1 _20345_ (.A(net237),
    .B(_03066_),
    .Y(_03181_));
 sg13g2_and2_1 _20346_ (.A(_08311_),
    .B(net146),
    .X(_03182_));
 sg13g2_buf_1 _20347_ (.A(_03182_),
    .X(_03183_));
 sg13g2_a22oi_1 _20348_ (.Y(_03184_),
    .B1(_03181_),
    .B2(_03183_),
    .A2(_03180_),
    .A1(net343));
 sg13g2_nand2_1 _20349_ (.Y(_03185_),
    .A(\cpu.dec.imm[5] ),
    .B(net108));
 sg13g2_o21ai_1 _20350_ (.B1(_03185_),
    .Y(_00767_),
    .A1(net92),
    .A2(_03184_));
 sg13g2_buf_1 _20351_ (.A(_03048_),
    .X(_03186_));
 sg13g2_a21o_1 _20352_ (.A2(_03186_),
    .A1(_02966_),
    .B1(_02963_),
    .X(_03187_));
 sg13g2_nor2_1 _20353_ (.A(_02975_),
    .B(net237),
    .Y(_03188_));
 sg13g2_a22oi_1 _20354_ (.Y(_03189_),
    .B1(_03188_),
    .B2(_02969_),
    .A2(_03187_),
    .A1(_08249_));
 sg13g2_a21oi_1 _20355_ (.A1(_03072_),
    .A2(_03148_),
    .Y(_03190_),
    .B1(net125));
 sg13g2_nor2_1 _20356_ (.A(_03154_),
    .B(_03156_),
    .Y(_03191_));
 sg13g2_o21ai_1 _20357_ (.B1(net346),
    .Y(_03192_),
    .A1(_03190_),
    .A2(_03191_));
 sg13g2_nor2_1 _20358_ (.A(net315),
    .B(_08886_),
    .Y(_03193_));
 sg13g2_nand2_1 _20359_ (.Y(_03194_),
    .A(net146),
    .B(_03149_));
 sg13g2_a21oi_1 _20360_ (.A1(net181),
    .A2(_03193_),
    .Y(_03195_),
    .B1(_03194_));
 sg13g2_a21oi_1 _20361_ (.A1(_03189_),
    .A2(_03192_),
    .Y(_03196_),
    .B1(_03195_));
 sg13g2_mux2_1 _20362_ (.A0(_03196_),
    .A1(\cpu.dec.imm[6] ),
    .S(net106),
    .X(_00768_));
 sg13g2_inv_1 _20363_ (.Y(_03197_),
    .A(\cpu.dec.imm[7] ));
 sg13g2_nand2_1 _20364_ (.Y(_03198_),
    .A(net240),
    .B(net146));
 sg13g2_a21o_1 _20365_ (.A2(net207),
    .A1(net202),
    .B1(_03078_),
    .X(_03199_));
 sg13g2_nand2b_1 _20366_ (.Y(_03200_),
    .B(_03169_),
    .A_N(_03138_));
 sg13g2_o21ai_1 _20367_ (.B1(_03200_),
    .Y(_03201_),
    .A1(_03198_),
    .A2(_03199_));
 sg13g2_a221oi_1 _20368_ (.B2(net203),
    .C1(_03201_),
    .B1(_03190_),
    .A1(net249),
    .Y(_03202_),
    .A2(_02971_));
 sg13g2_a22oi_1 _20369_ (.Y(_00769_),
    .B1(_03100_),
    .B2(_03202_),
    .A2(_03070_),
    .A1(_03197_));
 sg13g2_inv_1 _20370_ (.Y(_03203_),
    .A(\cpu.dec.imm[8] ));
 sg13g2_nand2_1 _20371_ (.Y(_03204_),
    .A(net343),
    .B(_03081_));
 sg13g2_nand2_1 _20372_ (.Y(_03205_),
    .A(_03083_),
    .B(_03204_));
 sg13g2_inv_1 _20373_ (.Y(_03206_),
    .A(net204));
 sg13g2_nor2_1 _20374_ (.A(_02991_),
    .B(_03206_),
    .Y(_03207_));
 sg13g2_o21ai_1 _20375_ (.B1(_03113_),
    .Y(_03208_),
    .A1(net343),
    .A2(net143));
 sg13g2_a21oi_1 _20376_ (.A1(_02966_),
    .A2(net204),
    .Y(_03209_),
    .B1(_03084_));
 sg13g2_a21oi_1 _20377_ (.A1(_03208_),
    .A2(_03209_),
    .Y(_03210_),
    .B1(_03074_));
 sg13g2_a221oi_1 _20378_ (.B2(_03183_),
    .C1(_03210_),
    .B1(_03207_),
    .A1(_03088_),
    .Y(_03211_),
    .A2(_03205_));
 sg13g2_a22oi_1 _20379_ (.Y(_00770_),
    .B1(_03100_),
    .B2(_03211_),
    .A2(_03070_),
    .A1(_03203_));
 sg13g2_o21ai_1 _20380_ (.B1(_03113_),
    .Y(_03212_),
    .A1(net346),
    .A2(net143));
 sg13g2_a21oi_1 _20381_ (.A1(net189),
    .A2(_02966_),
    .Y(_03213_),
    .B1(_03084_));
 sg13g2_nand2_1 _20382_ (.Y(_03214_),
    .A(_03212_),
    .B(_03213_));
 sg13g2_o21ai_1 _20383_ (.B1(_03083_),
    .Y(_03215_),
    .A1(_09723_),
    .A2(_03091_));
 sg13g2_a22oi_1 _20384_ (.Y(_03216_),
    .B1(_03215_),
    .B2(_03088_),
    .A2(_03214_),
    .A1(_03075_));
 sg13g2_a22oi_1 _20385_ (.Y(_00771_),
    .B1(_03100_),
    .B2(_03216_),
    .A2(net92),
    .A1(_11048_));
 sg13g2_buf_1 _20386_ (.A(net911),
    .X(_03217_));
 sg13g2_nand3_1 _20387_ (.B(_09721_),
    .C(_03051_),
    .A(net719),
    .Y(_03218_));
 sg13g2_buf_2 _20388_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03219_));
 sg13g2_buf_1 _20389_ (.A(_08840_),
    .X(_03220_));
 sg13g2_nand2_1 _20390_ (.Y(_03221_),
    .A(_03219_),
    .B(net98));
 sg13g2_o21ai_1 _20391_ (.B1(_03221_),
    .Y(_00772_),
    .A1(net110),
    .A2(_03218_));
 sg13g2_nand2_1 _20392_ (.Y(_03222_),
    .A(_09720_),
    .B(_03158_));
 sg13g2_nand2_1 _20393_ (.Y(_03223_),
    .A(\cpu.dec.io ),
    .B(_03220_));
 sg13g2_o21ai_1 _20394_ (.B1(_03223_),
    .Y(_00773_),
    .A1(_08845_),
    .A2(_03222_));
 sg13g2_or2_1 _20395_ (.X(_03224_),
    .B(_08986_),
    .A(net346));
 sg13g2_buf_1 _20396_ (.A(_03224_),
    .X(_03225_));
 sg13g2_nor3_1 _20397_ (.A(_08881_),
    .B(_08946_),
    .C(_03225_),
    .Y(_03226_));
 sg13g2_buf_2 _20398_ (.A(_03226_),
    .X(_03227_));
 sg13g2_nand3_1 _20399_ (.B(_09742_),
    .C(_03227_),
    .A(_09730_),
    .Y(_03228_));
 sg13g2_nand2_1 _20400_ (.Y(_03229_),
    .A(\cpu.dec.jmp ),
    .B(net98));
 sg13g2_o21ai_1 _20401_ (.B1(_03229_),
    .Y(_00774_),
    .A1(net110),
    .A2(_03228_));
 sg13g2_nand2_1 _20402_ (.Y(_03230_),
    .A(_02981_),
    .B(net315));
 sg13g2_a21oi_1 _20403_ (.A1(net160),
    .A2(net207),
    .Y(_03231_),
    .B1(net145));
 sg13g2_nor3_1 _20404_ (.A(net109),
    .B(_03230_),
    .C(_03231_),
    .Y(_03232_));
 sg13g2_a21o_1 _20405_ (.A2(net111),
    .A1(_11337_),
    .B1(_03232_),
    .X(_00775_));
 sg13g2_nor3_1 _20406_ (.A(net109),
    .B(_08991_),
    .C(_08926_),
    .Y(_03233_));
 sg13g2_a21o_1 _20407_ (.A2(_08841_),
    .A1(_09197_),
    .B1(_03233_),
    .X(_00776_));
 sg13g2_nor3_1 _20408_ (.A(net161),
    .B(net206),
    .C(_08888_),
    .Y(_03234_));
 sg13g2_nor3_1 _20409_ (.A(net164),
    .B(net202),
    .C(net165),
    .Y(_03235_));
 sg13g2_nor3_1 _20410_ (.A(_08884_),
    .B(_03234_),
    .C(_03235_),
    .Y(_03236_));
 sg13g2_a21oi_1 _20411_ (.A1(_08887_),
    .A2(net165),
    .Y(_03237_),
    .B1(_08888_));
 sg13g2_nor3_1 _20412_ (.A(net160),
    .B(_08311_),
    .C(_03237_),
    .Y(_03238_));
 sg13g2_a21oi_1 _20413_ (.A1(net144),
    .A2(_03236_),
    .Y(_03239_),
    .B1(_03238_));
 sg13g2_nor3_1 _20414_ (.A(net109),
    .B(net146),
    .C(_03239_),
    .Y(_03240_));
 sg13g2_a21o_1 _20415_ (.A2(net111),
    .A1(_10950_),
    .B1(_03240_),
    .X(_00777_));
 sg13g2_nor2_1 _20416_ (.A(net181),
    .B(_03227_),
    .Y(_03241_));
 sg13g2_a21oi_1 _20417_ (.A1(_08917_),
    .A2(_03227_),
    .Y(_03242_),
    .B1(_03241_));
 sg13g2_a22oi_1 _20418_ (.Y(_03243_),
    .B1(_03242_),
    .B2(net147),
    .A2(net181),
    .A1(net206));
 sg13g2_a21oi_1 _20419_ (.A1(_03077_),
    .A2(net181),
    .Y(_03244_),
    .B1(_03095_));
 sg13g2_nand2_1 _20420_ (.Y(_03245_),
    .A(_03077_),
    .B(net146));
 sg13g2_inv_1 _20421_ (.Y(_03246_),
    .A(_03245_));
 sg13g2_o21ai_1 _20422_ (.B1(_03246_),
    .Y(_03247_),
    .A1(net202),
    .A2(net343));
 sg13g2_o21ai_1 _20423_ (.B1(_03247_),
    .Y(_03248_),
    .A1(net125),
    .A2(_03244_));
 sg13g2_mux2_1 _20424_ (.A0(net181),
    .A1(net343),
    .S(net241),
    .X(_03249_));
 sg13g2_a22oi_1 _20425_ (.Y(_03250_),
    .B1(_03104_),
    .B2(_03249_),
    .A2(net181),
    .A1(net147));
 sg13g2_nor2_1 _20426_ (.A(net121),
    .B(_03250_),
    .Y(_03251_));
 sg13g2_a21oi_1 _20427_ (.A1(_02989_),
    .A2(_03248_),
    .Y(_03252_),
    .B1(_03251_));
 sg13g2_o21ai_1 _20428_ (.B1(_03252_),
    .Y(_03253_),
    .A1(_03154_),
    .A2(_03243_));
 sg13g2_mux2_1 _20429_ (.A0(_03253_),
    .A1(\cpu.dec.r_rd[0] ),
    .S(_09768_),
    .X(_00778_));
 sg13g2_nor2_1 _20430_ (.A(net202),
    .B(_03245_),
    .Y(_03254_));
 sg13g2_o21ai_1 _20431_ (.B1(net202),
    .Y(_03255_),
    .A1(_08884_),
    .A2(_03227_));
 sg13g2_a21oi_1 _20432_ (.A1(_08884_),
    .A2(_03230_),
    .Y(_03256_),
    .B1(net125));
 sg13g2_a21o_1 _20433_ (.A2(_03255_),
    .A1(_09742_),
    .B1(_03256_),
    .X(_03257_));
 sg13g2_a21oi_1 _20434_ (.A1(net315),
    .A2(_09723_),
    .Y(_03258_),
    .B1(net239));
 sg13g2_nor2_1 _20435_ (.A(net238),
    .B(_03078_),
    .Y(_03259_));
 sg13g2_o21ai_1 _20436_ (.B1(net207),
    .Y(_03260_),
    .A1(_03258_),
    .A2(_03259_));
 sg13g2_nand3b_1 _20437_ (.B(net205),
    .C(_03104_),
    .Y(_03261_),
    .A_N(net207));
 sg13g2_nand2_1 _20438_ (.Y(_03262_),
    .A(_08880_),
    .B(_08946_));
 sg13g2_or4_1 _20439_ (.A(_08990_),
    .B(net190),
    .C(_03050_),
    .D(_03262_),
    .X(_03263_));
 sg13g2_or2_1 _20440_ (.X(_03264_),
    .B(_03263_),
    .A(_09763_));
 sg13g2_a221oi_1 _20441_ (.B2(_09741_),
    .C1(net121),
    .B1(_03264_),
    .A1(_03260_),
    .Y(_03265_),
    .A2(_03261_));
 sg13g2_a221oi_1 _20442_ (.B2(net205),
    .C1(_03265_),
    .B1(_03257_),
    .A1(net346),
    .Y(_03266_),
    .A2(_03254_));
 sg13g2_nand2_1 _20443_ (.Y(_03267_),
    .A(\cpu.dec.r_rd[1] ),
    .B(net98));
 sg13g2_o21ai_1 _20444_ (.B1(_03267_),
    .Y(_00779_),
    .A1(_08845_),
    .A2(_03266_));
 sg13g2_nor2_1 _20445_ (.A(net241),
    .B(net204),
    .Y(_03268_));
 sg13g2_a21oi_1 _20446_ (.A1(net207),
    .A2(_03089_),
    .Y(_03269_),
    .B1(_03268_));
 sg13g2_a22oi_1 _20447_ (.Y(_03270_),
    .B1(_03104_),
    .B2(_03269_),
    .A2(net204),
    .A1(net147));
 sg13g2_nor2_1 _20448_ (.A(net121),
    .B(_03270_),
    .Y(_03271_));
 sg13g2_a221oi_1 _20449_ (.B2(net204),
    .C1(_03271_),
    .B1(_03257_),
    .A1(net203),
    .Y(_03272_),
    .A2(_03254_));
 sg13g2_nand2_1 _20450_ (.Y(_03273_),
    .A(\cpu.dec.r_rd[2] ),
    .B(net98));
 sg13g2_o21ai_1 _20451_ (.B1(_03273_),
    .Y(_00780_),
    .A1(net110),
    .A2(_03272_));
 sg13g2_inv_1 _20452_ (.Y(_03274_),
    .A(\cpu.dec.r_rd[3] ));
 sg13g2_a21oi_1 _20453_ (.A1(net315),
    .A2(net189),
    .Y(_03275_),
    .B1(net241));
 sg13g2_o21ai_1 _20454_ (.B1(_03230_),
    .Y(_03276_),
    .A1(_08311_),
    .A2(_03227_));
 sg13g2_a21oi_1 _20455_ (.A1(net189),
    .A2(_03276_),
    .Y(_03277_),
    .B1(_08223_));
 sg13g2_nor3_1 _20456_ (.A(net161),
    .B(net166),
    .C(_03104_),
    .Y(_03278_));
 sg13g2_nor4_1 _20457_ (.A(_02969_),
    .B(_03275_),
    .C(_03277_),
    .D(_03278_),
    .Y(_03279_));
 sg13g2_o21ai_1 _20458_ (.B1(net144),
    .Y(_03280_),
    .A1(_09741_),
    .A2(_03279_));
 sg13g2_inv_1 _20459_ (.Y(_03281_),
    .A(_03143_));
 sg13g2_a21oi_1 _20460_ (.A1(net144),
    .A2(_03281_),
    .Y(_03282_),
    .B1(_03279_));
 sg13g2_a21oi_1 _20461_ (.A1(_02975_),
    .A2(_03280_),
    .Y(_03283_),
    .B1(_03282_));
 sg13g2_nor3_1 _20462_ (.A(_09761_),
    .B(_03254_),
    .C(_03283_),
    .Y(_03284_));
 sg13g2_a21oi_1 _20463_ (.A1(_03274_),
    .A2(net86),
    .Y(_00781_),
    .B1(_03284_));
 sg13g2_o21ai_1 _20464_ (.B1(_08886_),
    .Y(_03285_),
    .A1(_08915_),
    .A2(_03227_));
 sg13g2_inv_1 _20465_ (.Y(_03286_),
    .A(_03285_));
 sg13g2_o21ai_1 _20466_ (.B1(_09742_),
    .Y(_03287_),
    .A1(_03193_),
    .A2(_03286_));
 sg13g2_a21oi_1 _20467_ (.A1(_03077_),
    .A2(_03230_),
    .Y(_03288_),
    .B1(net160));
 sg13g2_o21ai_1 _20468_ (.B1(net164),
    .Y(_03289_),
    .A1(_03081_),
    .A2(_03288_));
 sg13g2_o21ai_1 _20469_ (.B1(_02992_),
    .Y(_03290_),
    .A1(net145),
    .A2(_09741_));
 sg13g2_nand2_1 _20470_ (.Y(_03291_),
    .A(_03289_),
    .B(_03290_));
 sg13g2_a22oi_1 _20471_ (.Y(_03292_),
    .B1(_03186_),
    .B2(_03198_),
    .A2(net146),
    .A1(net147));
 sg13g2_a21oi_1 _20472_ (.A1(_03287_),
    .A2(_03291_),
    .Y(_03293_),
    .B1(_03292_));
 sg13g2_mux2_1 _20473_ (.A0(_03293_),
    .A1(_10245_),
    .S(net91),
    .X(_00782_));
 sg13g2_o21ai_1 _20474_ (.B1(_03287_),
    .Y(_03294_),
    .A1(_08924_),
    .A2(_03081_));
 sg13g2_o21ai_1 _20475_ (.B1(_02981_),
    .Y(_03295_),
    .A1(net241),
    .A2(_03109_));
 sg13g2_a21oi_1 _20476_ (.A1(net315),
    .A2(_03295_),
    .Y(_03296_),
    .B1(_08309_));
 sg13g2_nor2_1 _20477_ (.A(_02976_),
    .B(_03296_),
    .Y(_03297_));
 sg13g2_o21ai_1 _20478_ (.B1(_03014_),
    .Y(_03298_),
    .A1(_03294_),
    .A2(_03297_));
 sg13g2_o21ai_1 _20479_ (.B1(_03298_),
    .Y(_03299_),
    .A1(net166),
    .A2(_02997_));
 sg13g2_a21oi_1 _20480_ (.A1(net205),
    .A2(_03294_),
    .Y(_03300_),
    .B1(net238));
 sg13g2_o21ai_1 _20481_ (.B1(_03183_),
    .Y(_03301_),
    .A1(net240),
    .A2(net205));
 sg13g2_o21ai_1 _20482_ (.B1(_03301_),
    .Y(_03302_),
    .A1(_03154_),
    .A2(_03300_));
 sg13g2_a21oi_1 _20483_ (.A1(net164),
    .A2(_03299_),
    .Y(_03303_),
    .B1(_03302_));
 sg13g2_nand2_1 _20484_ (.Y(_03304_),
    .A(_10277_),
    .B(net98));
 sg13g2_o21ai_1 _20485_ (.B1(_03304_),
    .Y(_00783_),
    .A1(net110),
    .A2(_03303_));
 sg13g2_nor3_1 _20486_ (.A(net125),
    .B(_02966_),
    .C(_03104_),
    .Y(_03305_));
 sg13g2_o21ai_1 _20487_ (.B1(_03206_),
    .Y(_03306_),
    .A1(net121),
    .A2(_02997_));
 sg13g2_o21ai_1 _20488_ (.B1(_03306_),
    .Y(_03307_),
    .A1(_03294_),
    .A2(_03305_));
 sg13g2_nand3_1 _20489_ (.B(net146),
    .C(net204),
    .A(net238),
    .Y(_03308_));
 sg13g2_a21oi_1 _20490_ (.A1(_03307_),
    .A2(_03308_),
    .Y(_03309_),
    .B1(net98));
 sg13g2_a21o_1 _20491_ (.A2(_08841_),
    .A1(_10275_),
    .B1(_03309_),
    .X(_00784_));
 sg13g2_nor2_1 _20492_ (.A(net164),
    .B(_02974_),
    .Y(_03310_));
 sg13g2_a21oi_1 _20493_ (.A1(net164),
    .A2(_08309_),
    .Y(_03311_),
    .B1(_03310_));
 sg13g2_nor2_1 _20494_ (.A(_09729_),
    .B(_03193_),
    .Y(_03312_));
 sg13g2_o21ai_1 _20495_ (.B1(_03312_),
    .Y(_03313_),
    .A1(_08335_),
    .A2(_03285_));
 sg13g2_o21ai_1 _20496_ (.B1(_03313_),
    .Y(_03314_),
    .A1(_03137_),
    .A2(_03311_));
 sg13g2_and2_1 _20497_ (.A(net164),
    .B(net207),
    .X(_03315_));
 sg13g2_nor3_1 _20498_ (.A(net144),
    .B(net238),
    .C(_03315_),
    .Y(_03316_));
 sg13g2_a221oi_1 _20499_ (.B2(net144),
    .C1(_03316_),
    .B1(_03314_),
    .A1(_03104_),
    .Y(_03317_),
    .A2(_03231_));
 sg13g2_mux2_1 _20500_ (.A0(_03317_),
    .A1(_10235_),
    .S(net106),
    .X(_00785_));
 sg13g2_nor2_1 _20501_ (.A(_03154_),
    .B(_02989_),
    .Y(_03318_));
 sg13g2_nand3_1 _20502_ (.B(_08950_),
    .C(_03225_),
    .A(_08888_),
    .Y(_03319_));
 sg13g2_a221oi_1 _20503_ (.B2(_08886_),
    .C1(net161),
    .B1(_03319_),
    .A1(net206),
    .Y(_03320_),
    .A2(_02966_));
 sg13g2_nor2_1 _20504_ (.A(net164),
    .B(_02989_),
    .Y(_03321_));
 sg13g2_o21ai_1 _20505_ (.B1(net144),
    .Y(_03322_),
    .A1(_03320_),
    .A2(_03321_));
 sg13g2_a221oi_1 _20506_ (.B2(net343),
    .C1(_09761_),
    .B1(_03322_),
    .A1(net181),
    .Y(_03323_),
    .A2(_03318_));
 sg13g2_a21oi_1 _20507_ (.A1(net662),
    .A2(net91),
    .Y(_00786_),
    .B1(_03323_));
 sg13g2_a221oi_1 _20508_ (.B2(net346),
    .C1(_09761_),
    .B1(_03322_),
    .A1(net205),
    .Y(_03324_),
    .A2(_03318_));
 sg13g2_a21oi_1 _20509_ (.A1(net661),
    .A2(net91),
    .Y(_00787_),
    .B1(_03324_));
 sg13g2_nand2b_1 _20510_ (.Y(_03325_),
    .B(net239),
    .A_N(net207));
 sg13g2_a21oi_1 _20511_ (.A1(_03072_),
    .A2(_03325_),
    .Y(_03326_),
    .B1(net145));
 sg13g2_a21oi_1 _20512_ (.A1(net145),
    .A2(net206),
    .Y(_03327_),
    .B1(net240));
 sg13g2_o21ai_1 _20513_ (.B1(net144),
    .Y(_03328_),
    .A1(_03326_),
    .A2(_03327_));
 sg13g2_a221oi_1 _20514_ (.B2(net203),
    .C1(_09761_),
    .B1(_03328_),
    .A1(net204),
    .Y(_03329_),
    .A2(_03318_));
 sg13g2_a21oi_1 _20515_ (.A1(net650),
    .A2(net91),
    .Y(_00788_),
    .B1(_03329_));
 sg13g2_a22oi_1 _20516_ (.Y(_03330_),
    .B1(_08880_),
    .B2(_08309_),
    .A2(_08335_),
    .A1(net238));
 sg13g2_nand3b_1 _20517_ (.B(net202),
    .C(net145),
    .Y(_03331_),
    .A_N(_03330_));
 sg13g2_nor2b_1 _20518_ (.A(_03320_),
    .B_N(_03331_),
    .Y(_03332_));
 sg13g2_nor3_1 _20519_ (.A(_03220_),
    .B(net166),
    .C(_03332_),
    .Y(_03333_));
 sg13g2_a21oi_1 _20520_ (.A1(_10859_),
    .A2(net86),
    .Y(_00789_),
    .B1(_03333_));
 sg13g2_mux2_1 _20521_ (.A0(_08988_),
    .A1(_10163_),
    .S(net106),
    .X(_00790_));
 sg13g2_nor3_1 _20522_ (.A(net109),
    .B(_08951_),
    .C(_03225_),
    .Y(_03334_));
 sg13g2_a21o_1 _20523_ (.A2(net111),
    .A1(_10076_),
    .B1(_03334_),
    .X(_00791_));
 sg13g2_nor4_1 _20524_ (.A(net125),
    .B(net249),
    .C(_08889_),
    .D(_08917_),
    .Y(_03335_));
 sg13g2_mux2_1 _20525_ (.A0(_03335_),
    .A1(\cpu.dec.r_set_cc ),
    .S(net106),
    .X(_00792_));
 sg13g2_a21oi_1 _20526_ (.A1(_09720_),
    .A2(_02966_),
    .Y(_03336_),
    .B1(_03321_));
 sg13g2_buf_1 _20527_ (.A(\cpu.dec.r_store ),
    .X(_03337_));
 sg13g2_nand2_1 _20528_ (.Y(_03338_),
    .A(_03337_),
    .B(net98));
 sg13g2_o21ai_1 _20529_ (.B1(_03338_),
    .Y(_00793_),
    .A1(net110),
    .A2(_03336_));
 sg13g2_nor3_1 _20530_ (.A(net121),
    .B(_02997_),
    .C(_03264_),
    .Y(_03339_));
 sg13g2_mux2_1 _20531_ (.A0(_03339_),
    .A1(\cpu.dec.r_swapsp ),
    .S(net108),
    .X(_00794_));
 sg13g2_nor4_1 _20532_ (.A(_08840_),
    .B(_09725_),
    .C(_02997_),
    .D(_03263_),
    .Y(_03340_));
 sg13g2_a21o_1 _20533_ (.A2(net111),
    .A1(\cpu.dec.r_sys_call ),
    .B1(_03340_),
    .X(_00795_));
 sg13g2_a21oi_1 _20534_ (.A1(net240),
    .A2(_03285_),
    .Y(_03341_),
    .B1(_09731_));
 sg13g2_nand2_1 _20535_ (.Y(_03342_),
    .A(net205),
    .B(net181));
 sg13g2_xnor2_1 _20536_ (.Y(_03343_),
    .A(_03206_),
    .B(_03342_));
 sg13g2_nor2_1 _20537_ (.A(net719),
    .B(_03343_),
    .Y(_03344_));
 sg13g2_o21ai_1 _20538_ (.B1(_03344_),
    .Y(_03345_),
    .A1(_03095_),
    .A2(_03341_));
 sg13g2_o21ai_1 _20539_ (.B1(_09741_),
    .Y(_03346_),
    .A1(net190),
    .A2(_09724_));
 sg13g2_a21o_1 _20540_ (.A2(_08991_),
    .A1(_08920_),
    .B1(_03346_),
    .X(_03347_));
 sg13g2_xnor2_1 _20541_ (.Y(_03348_),
    .A(net203),
    .B(_08987_));
 sg13g2_nor2_1 _20542_ (.A(_08737_),
    .B(net190),
    .Y(_03349_));
 sg13g2_a21oi_1 _20543_ (.A1(net911),
    .A2(net190),
    .Y(_03350_),
    .B1(_03349_));
 sg13g2_nand4_1 _20544_ (.B(_08880_),
    .C(_03348_),
    .A(_08886_),
    .Y(_03351_),
    .D(_03350_));
 sg13g2_nand4_1 _20545_ (.B(_03345_),
    .C(_03347_),
    .A(_03054_),
    .Y(_03352_),
    .D(_03351_));
 sg13g2_nor2_1 _20546_ (.A(net191),
    .B(_08916_),
    .Y(_03353_));
 sg13g2_nand2_1 _20547_ (.Y(_03354_),
    .A(_09731_),
    .B(net249));
 sg13g2_o21ai_1 _20548_ (.B1(_03354_),
    .Y(_03355_),
    .A1(_08355_),
    .A2(_08920_));
 sg13g2_a22oi_1 _20549_ (.Y(_03356_),
    .B1(_03355_),
    .B2(net165),
    .A2(_03353_),
    .A1(_09724_));
 sg13g2_nor4_1 _20550_ (.A(_08368_),
    .B(net189),
    .C(_03091_),
    .D(_03343_),
    .Y(_03357_));
 sg13g2_nor2_1 _20551_ (.A(net161),
    .B(_03357_),
    .Y(_03358_));
 sg13g2_o21ai_1 _20552_ (.B1(_03358_),
    .Y(_03359_),
    .A1(_08311_),
    .A2(_03356_));
 sg13g2_nand4_1 _20553_ (.B(_08881_),
    .C(_08916_),
    .A(_08334_),
    .Y(_03360_),
    .D(_08949_));
 sg13g2_a21oi_1 _20554_ (.A1(_08355_),
    .A2(_03360_),
    .Y(_03361_),
    .B1(_08884_));
 sg13g2_nand4_1 _20555_ (.B(_08917_),
    .C(_09712_),
    .A(net911),
    .Y(_03362_),
    .D(_03227_));
 sg13g2_nor2b_1 _20556_ (.A(_03054_),
    .B_N(_03362_),
    .Y(_03363_));
 sg13g2_nor2_1 _20557_ (.A(_08368_),
    .B(_10416_),
    .Y(_03364_));
 sg13g2_a21oi_1 _20558_ (.A1(_03079_),
    .A2(_03364_),
    .Y(_03365_),
    .B1(_08309_));
 sg13g2_nor2_1 _20559_ (.A(net239),
    .B(_03365_),
    .Y(_03366_));
 sg13g2_nor4_1 _20560_ (.A(_03357_),
    .B(_03361_),
    .C(_03363_),
    .D(_03366_),
    .Y(_03367_));
 sg13g2_nor2_1 _20561_ (.A(_02997_),
    .B(_03050_),
    .Y(_03368_));
 sg13g2_nor2_1 _20562_ (.A(net249),
    .B(_08947_),
    .Y(_03369_));
 sg13g2_o21ai_1 _20563_ (.B1(_03369_),
    .Y(_03370_),
    .A1(_09763_),
    .A2(_03262_));
 sg13g2_and4_1 _20564_ (.A(net719),
    .B(_08917_),
    .C(_03368_),
    .D(_03370_),
    .X(_03371_));
 sg13g2_nor3_1 _20565_ (.A(_02987_),
    .B(_03367_),
    .C(_03371_),
    .Y(_03372_));
 sg13g2_a221oi_1 _20566_ (.B2(net166),
    .C1(_03372_),
    .B1(_03359_),
    .A1(net145),
    .Y(_03373_),
    .A2(_03352_));
 sg13g2_nand2_1 _20567_ (.Y(_03374_),
    .A(net237),
    .B(_03049_));
 sg13g2_a221oi_1 _20568_ (.B2(_09730_),
    .C1(_03245_),
    .B1(_03374_),
    .A1(_03227_),
    .Y(_03375_),
    .A2(_03368_));
 sg13g2_nor3_1 _20569_ (.A(_09761_),
    .B(_03373_),
    .C(_03375_),
    .Y(_03376_));
 sg13g2_a21o_1 _20570_ (.A2(net111),
    .A1(_09018_),
    .B1(_03376_),
    .X(_00796_));
 sg13g2_buf_1 _20571_ (.A(net1032),
    .X(_03377_));
 sg13g2_buf_1 _20572_ (.A(_03377_),
    .X(_03378_));
 sg13g2_nand2b_1 _20573_ (.Y(_03379_),
    .B(net1011),
    .A_N(net1010));
 sg13g2_buf_1 _20574_ (.A(_03379_),
    .X(_03380_));
 sg13g2_nand3_1 _20575_ (.B(_10058_),
    .C(net1097),
    .A(net1096),
    .Y(_03381_));
 sg13g2_buf_1 _20576_ (.A(_03381_),
    .X(_03382_));
 sg13g2_nor2_1 _20577_ (.A(_03380_),
    .B(_03382_),
    .Y(_03383_));
 sg13g2_buf_2 _20578_ (.A(_03383_),
    .X(_03384_));
 sg13g2_buf_1 _20579_ (.A(_03384_),
    .X(_03385_));
 sg13g2_mux2_1 _20580_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net718),
    .S(net530),
    .X(_00801_));
 sg13g2_mux2_1 _20581_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net843),
    .S(_03385_),
    .X(_00802_));
 sg13g2_mux2_1 _20582_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net842),
    .S(_03385_),
    .X(_00803_));
 sg13g2_buf_1 _20583_ (.A(net675),
    .X(_03386_));
 sg13g2_buf_1 _20584_ (.A(net595),
    .X(_03387_));
 sg13g2_mux2_1 _20585_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net529),
    .S(net530),
    .X(_00804_));
 sg13g2_buf_1 _20586_ (.A(net611),
    .X(_03388_));
 sg13g2_buf_1 _20587_ (.A(net528),
    .X(_03389_));
 sg13g2_mux2_1 _20588_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net470),
    .S(net530),
    .X(_00805_));
 sg13g2_buf_1 _20589_ (.A(net672),
    .X(_03390_));
 sg13g2_buf_1 _20590_ (.A(net594),
    .X(_03391_));
 sg13g2_mux2_1 _20591_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net527),
    .S(net530),
    .X(_00806_));
 sg13g2_buf_1 _20592_ (.A(net890),
    .X(_03392_));
 sg13g2_buf_1 _20593_ (.A(net717),
    .X(_03393_));
 sg13g2_mux2_1 _20594_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net642),
    .S(net530),
    .X(_00807_));
 sg13g2_mux2_1 _20595_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net544),
    .S(net530),
    .X(_00808_));
 sg13g2_buf_1 _20596_ (.A(net551),
    .X(_03394_));
 sg13g2_buf_1 _20597_ (.A(net469),
    .X(_03395_));
 sg13g2_mux2_1 _20598_ (.A0(\cpu.ex.r_10[2] ),
    .A1(net406),
    .S(net530),
    .X(_00809_));
 sg13g2_buf_1 _20599_ (.A(net496),
    .X(_03396_));
 sg13g2_mux2_1 _20600_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net405),
    .S(net530),
    .X(_00810_));
 sg13g2_buf_2 _20601_ (.A(net424),
    .X(_03397_));
 sg13g2_buf_1 _20602_ (.A(net366),
    .X(_03398_));
 sg13g2_buf_1 _20603_ (.A(net335),
    .X(_03399_));
 sg13g2_mux2_1 _20604_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net314),
    .S(_03384_),
    .X(_00811_));
 sg13g2_mux2_1 _20605_ (.A0(\cpu.ex.r_10[5] ),
    .A1(net596),
    .S(_03384_),
    .X(_00812_));
 sg13g2_mux2_1 _20606_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net722),
    .S(_03384_),
    .X(_00813_));
 sg13g2_mux2_1 _20607_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net721),
    .S(_03384_),
    .X(_00814_));
 sg13g2_mux2_1 _20608_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net720),
    .S(_03384_),
    .X(_00815_));
 sg13g2_mux2_1 _20609_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net844),
    .S(_03384_),
    .X(_00816_));
 sg13g2_nand2_1 _20610_ (.Y(_03400_),
    .A(net1011),
    .B(net1010));
 sg13g2_nor2_1 _20611_ (.A(_03400_),
    .B(_03382_),
    .Y(_03401_));
 sg13g2_buf_2 _20612_ (.A(_03401_),
    .X(_03402_));
 sg13g2_buf_1 _20613_ (.A(_03402_),
    .X(_03403_));
 sg13g2_mux2_1 _20614_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net718),
    .S(net526),
    .X(_00817_));
 sg13g2_mux2_1 _20615_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net843),
    .S(net526),
    .X(_00818_));
 sg13g2_mux2_1 _20616_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net842),
    .S(_03403_),
    .X(_00819_));
 sg13g2_mux2_1 _20617_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net529),
    .S(net526),
    .X(_00820_));
 sg13g2_mux2_1 _20618_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net470),
    .S(net526),
    .X(_00821_));
 sg13g2_mux2_1 _20619_ (.A0(\cpu.ex.r_11[14] ),
    .A1(net527),
    .S(net526),
    .X(_00822_));
 sg13g2_mux2_1 _20620_ (.A0(\cpu.ex.r_11[15] ),
    .A1(_03393_),
    .S(net526),
    .X(_00823_));
 sg13g2_mux2_1 _20621_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net544),
    .S(_03403_),
    .X(_00824_));
 sg13g2_mux2_1 _20622_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net406),
    .S(net526),
    .X(_00825_));
 sg13g2_mux2_1 _20623_ (.A0(\cpu.ex.r_11[3] ),
    .A1(net405),
    .S(net526),
    .X(_00826_));
 sg13g2_mux2_1 _20624_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net314),
    .S(_03402_),
    .X(_00827_));
 sg13g2_mux2_1 _20625_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net596),
    .S(_03402_),
    .X(_00828_));
 sg13g2_mux2_1 _20626_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net722),
    .S(_03402_),
    .X(_00829_));
 sg13g2_mux2_1 _20627_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net721),
    .S(_03402_),
    .X(_00830_));
 sg13g2_mux2_1 _20628_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net720),
    .S(_03402_),
    .X(_00831_));
 sg13g2_mux2_1 _20629_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net844),
    .S(_03402_),
    .X(_00832_));
 sg13g2_nand3_1 _20630_ (.B(_10057_),
    .C(net1097),
    .A(net1096),
    .Y(_03404_));
 sg13g2_buf_1 _20631_ (.A(_03404_),
    .X(_03405_));
 sg13g2_nor3_1 _20632_ (.A(_10052_),
    .B(net1010),
    .C(_03405_),
    .Y(_03406_));
 sg13g2_buf_4 _20633_ (.X(_03407_),
    .A(_03406_));
 sg13g2_buf_1 _20634_ (.A(_03407_),
    .X(_03408_));
 sg13g2_mux2_1 _20635_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net718),
    .S(net593),
    .X(_00833_));
 sg13g2_mux2_1 _20636_ (.A0(\cpu.ex.r_12[10] ),
    .A1(net843),
    .S(net593),
    .X(_00834_));
 sg13g2_mux2_1 _20637_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net842),
    .S(net593),
    .X(_00835_));
 sg13g2_mux2_1 _20638_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net529),
    .S(net593),
    .X(_00836_));
 sg13g2_mux2_1 _20639_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net470),
    .S(_03408_),
    .X(_00837_));
 sg13g2_mux2_1 _20640_ (.A0(\cpu.ex.r_12[14] ),
    .A1(_03391_),
    .S(net593),
    .X(_00838_));
 sg13g2_mux2_1 _20641_ (.A0(\cpu.ex.r_12[15] ),
    .A1(_03393_),
    .S(net593),
    .X(_00839_));
 sg13g2_mux2_1 _20642_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net544),
    .S(net593),
    .X(_00840_));
 sg13g2_mux2_1 _20643_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net406),
    .S(net593),
    .X(_00841_));
 sg13g2_mux2_1 _20644_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net405),
    .S(_03407_),
    .X(_00842_));
 sg13g2_nand2_1 _20645_ (.Y(_03409_),
    .A(net335),
    .B(_03407_));
 sg13g2_o21ai_1 _20646_ (.B1(_03409_),
    .Y(_00843_),
    .A1(_10774_),
    .A2(_03408_));
 sg13g2_mux2_1 _20647_ (.A0(\cpu.ex.r_12[5] ),
    .A1(net596),
    .S(_03407_),
    .X(_00844_));
 sg13g2_mux2_1 _20648_ (.A0(\cpu.ex.r_12[6] ),
    .A1(net722),
    .S(_03407_),
    .X(_00845_));
 sg13g2_mux2_1 _20649_ (.A0(\cpu.ex.r_12[7] ),
    .A1(net721),
    .S(_03407_),
    .X(_00846_));
 sg13g2_mux2_1 _20650_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net720),
    .S(_03407_),
    .X(_00847_));
 sg13g2_mux2_1 _20651_ (.A0(\cpu.ex.r_12[9] ),
    .A1(net844),
    .S(_03407_),
    .X(_00848_));
 sg13g2_inv_1 _20652_ (.Y(_03410_),
    .A(net1011));
 sg13g2_nand2_1 _20653_ (.Y(_03411_),
    .A(_03410_),
    .B(_10054_));
 sg13g2_nor2_1 _20654_ (.A(_03405_),
    .B(_03411_),
    .Y(_03412_));
 sg13g2_buf_2 _20655_ (.A(_03412_),
    .X(_03413_));
 sg13g2_buf_1 _20656_ (.A(_03413_),
    .X(_03414_));
 sg13g2_mux2_1 _20657_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net718),
    .S(net525),
    .X(_00849_));
 sg13g2_mux2_1 _20658_ (.A0(\cpu.ex.r_13[10] ),
    .A1(net843),
    .S(net525),
    .X(_00850_));
 sg13g2_mux2_1 _20659_ (.A0(\cpu.ex.r_13[11] ),
    .A1(_02944_),
    .S(net525),
    .X(_00851_));
 sg13g2_mux2_1 _20660_ (.A0(\cpu.ex.r_13[12] ),
    .A1(_03387_),
    .S(net525),
    .X(_00852_));
 sg13g2_buf_1 _20661_ (.A(net528),
    .X(_03415_));
 sg13g2_mux2_1 _20662_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net468),
    .S(net525),
    .X(_00853_));
 sg13g2_buf_1 _20663_ (.A(_03390_),
    .X(_03416_));
 sg13g2_mux2_1 _20664_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net524),
    .S(net525),
    .X(_00854_));
 sg13g2_buf_1 _20665_ (.A(net717),
    .X(_03417_));
 sg13g2_mux2_1 _20666_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net641),
    .S(_03414_),
    .X(_00855_));
 sg13g2_mux2_1 _20667_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net544),
    .S(net525),
    .X(_00856_));
 sg13g2_mux2_1 _20668_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net406),
    .S(_03414_),
    .X(_00857_));
 sg13g2_mux2_1 _20669_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net405),
    .S(net525),
    .X(_00858_));
 sg13g2_mux2_1 _20670_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net314),
    .S(_03413_),
    .X(_00859_));
 sg13g2_mux2_1 _20671_ (.A0(\cpu.ex.r_13[5] ),
    .A1(_02928_),
    .S(_03413_),
    .X(_00860_));
 sg13g2_mux2_1 _20672_ (.A0(\cpu.ex.r_13[6] ),
    .A1(_02938_),
    .S(_03413_),
    .X(_00861_));
 sg13g2_mux2_1 _20673_ (.A0(\cpu.ex.r_13[7] ),
    .A1(_02940_),
    .S(_03413_),
    .X(_00862_));
 sg13g2_mux2_1 _20674_ (.A0(\cpu.ex.r_13[8] ),
    .A1(_02941_),
    .S(_03413_),
    .X(_00863_));
 sg13g2_mux2_1 _20675_ (.A0(\cpu.ex.r_13[9] ),
    .A1(_02942_),
    .S(_03413_),
    .X(_00864_));
 sg13g2_nor2_1 _20676_ (.A(_03380_),
    .B(_03405_),
    .Y(_03418_));
 sg13g2_buf_2 _20677_ (.A(_03418_),
    .X(_03419_));
 sg13g2_buf_1 _20678_ (.A(_03419_),
    .X(_03420_));
 sg13g2_mux2_1 _20679_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net718),
    .S(net523),
    .X(_00865_));
 sg13g2_mux2_1 _20680_ (.A0(\cpu.ex.r_14[10] ),
    .A1(_02943_),
    .S(net523),
    .X(_00866_));
 sg13g2_mux2_1 _20681_ (.A0(\cpu.ex.r_14[11] ),
    .A1(_02944_),
    .S(_03420_),
    .X(_00867_));
 sg13g2_mux2_1 _20682_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net529),
    .S(net523),
    .X(_00868_));
 sg13g2_mux2_1 _20683_ (.A0(\cpu.ex.r_14[13] ),
    .A1(net468),
    .S(net523),
    .X(_00869_));
 sg13g2_mux2_1 _20684_ (.A0(\cpu.ex.r_14[14] ),
    .A1(net524),
    .S(net523),
    .X(_00870_));
 sg13g2_mux2_1 _20685_ (.A0(\cpu.ex.r_14[15] ),
    .A1(net641),
    .S(net523),
    .X(_00871_));
 sg13g2_mux2_1 _20686_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net544),
    .S(_03420_),
    .X(_00872_));
 sg13g2_mux2_1 _20687_ (.A0(\cpu.ex.r_14[2] ),
    .A1(net406),
    .S(net523),
    .X(_00873_));
 sg13g2_mux2_1 _20688_ (.A0(\cpu.ex.r_14[3] ),
    .A1(net405),
    .S(net523),
    .X(_00874_));
 sg13g2_mux2_1 _20689_ (.A0(\cpu.ex.r_14[4] ),
    .A1(net314),
    .S(_03419_),
    .X(_00875_));
 sg13g2_mux2_1 _20690_ (.A0(\cpu.ex.r_14[5] ),
    .A1(_02928_),
    .S(_03419_),
    .X(_00876_));
 sg13g2_mux2_1 _20691_ (.A0(\cpu.ex.r_14[6] ),
    .A1(_02938_),
    .S(_03419_),
    .X(_00877_));
 sg13g2_mux2_1 _20692_ (.A0(\cpu.ex.r_14[7] ),
    .A1(_02940_),
    .S(_03419_),
    .X(_00878_));
 sg13g2_mux2_1 _20693_ (.A0(\cpu.ex.r_14[8] ),
    .A1(_02941_),
    .S(_03419_),
    .X(_00879_));
 sg13g2_mux2_1 _20694_ (.A0(\cpu.ex.r_14[9] ),
    .A1(_02942_),
    .S(_03419_),
    .X(_00880_));
 sg13g2_nor2_1 _20695_ (.A(_03400_),
    .B(_03405_),
    .Y(_03421_));
 sg13g2_buf_2 _20696_ (.A(_03421_),
    .X(_03422_));
 sg13g2_buf_1 _20697_ (.A(_03422_),
    .X(_03423_));
 sg13g2_mux2_1 _20698_ (.A0(\cpu.ex.r_15[0] ),
    .A1(_03378_),
    .S(net592),
    .X(_00881_));
 sg13g2_mux2_1 _20699_ (.A0(\cpu.ex.r_15[10] ),
    .A1(_02943_),
    .S(net592),
    .X(_00882_));
 sg13g2_buf_1 _20700_ (.A(net1094),
    .X(_03424_));
 sg13g2_mux2_1 _20701_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net949),
    .S(net592),
    .X(_00883_));
 sg13g2_mux2_1 _20702_ (.A0(\cpu.ex.r_15[12] ),
    .A1(net529),
    .S(net592),
    .X(_00884_));
 sg13g2_mux2_1 _20703_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net468),
    .S(_03423_),
    .X(_00885_));
 sg13g2_mux2_1 _20704_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net524),
    .S(_03423_),
    .X(_00886_));
 sg13g2_mux2_1 _20705_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net641),
    .S(net592),
    .X(_00887_));
 sg13g2_mux2_1 _20706_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net544),
    .S(net592),
    .X(_00888_));
 sg13g2_mux2_1 _20707_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net406),
    .S(net592),
    .X(_00889_));
 sg13g2_mux2_1 _20708_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net405),
    .S(net592),
    .X(_00890_));
 sg13g2_mux2_1 _20709_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net314),
    .S(_03422_),
    .X(_00891_));
 sg13g2_buf_1 _20710_ (.A(net643),
    .X(_03425_));
 sg13g2_mux2_1 _20711_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net591),
    .S(_03422_),
    .X(_00892_));
 sg13g2_buf_1 _20712_ (.A(net953),
    .X(_03426_));
 sg13g2_mux2_1 _20713_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net840),
    .S(_03422_),
    .X(_00893_));
 sg13g2_buf_1 _20714_ (.A(net852),
    .X(_03427_));
 sg13g2_mux2_1 _20715_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net716),
    .S(_03422_),
    .X(_00894_));
 sg13g2_buf_1 _20716_ (.A(net851),
    .X(_03428_));
 sg13g2_mux2_1 _20717_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net715),
    .S(_03422_),
    .X(_00895_));
 sg13g2_buf_1 _20718_ (.A(net952),
    .X(_03429_));
 sg13g2_mux2_1 _20719_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net839),
    .S(_03422_),
    .X(_00896_));
 sg13g2_nor3_1 _20720_ (.A(net1011),
    .B(_10054_),
    .C(_03382_),
    .Y(_03430_));
 sg13g2_buf_1 _20721_ (.A(_03430_),
    .X(_03431_));
 sg13g2_buf_1 _20722_ (.A(net590),
    .X(_03432_));
 sg13g2_mux2_1 _20723_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net718),
    .S(net522),
    .X(_00897_));
 sg13g2_buf_1 _20724_ (.A(net951),
    .X(_03433_));
 sg13g2_mux2_1 _20725_ (.A0(\cpu.ex.r_8[10] ),
    .A1(net838),
    .S(net522),
    .X(_00898_));
 sg13g2_mux2_1 _20726_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net949),
    .S(net522),
    .X(_00899_));
 sg13g2_mux2_1 _20727_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net529),
    .S(net522),
    .X(_00900_));
 sg13g2_mux2_1 _20728_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net468),
    .S(net522),
    .X(_00901_));
 sg13g2_nand2_1 _20729_ (.Y(_03434_),
    .A(net594),
    .B(net590));
 sg13g2_o21ai_1 _20730_ (.B1(_03434_),
    .Y(_00902_),
    .A1(_10560_),
    .A2(_03432_));
 sg13g2_mux2_1 _20731_ (.A0(\cpu.ex.r_8[15] ),
    .A1(net641),
    .S(_03432_),
    .X(_00903_));
 sg13g2_mux2_1 _20732_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net544),
    .S(net522),
    .X(_00904_));
 sg13g2_nand2_1 _20733_ (.Y(_03435_),
    .A(net469),
    .B(net590));
 sg13g2_o21ai_1 _20734_ (.B1(_03435_),
    .Y(_00905_),
    .A1(_10835_),
    .A2(net522));
 sg13g2_mux2_1 _20735_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net405),
    .S(net590),
    .X(_00906_));
 sg13g2_mux2_1 _20736_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net314),
    .S(net590),
    .X(_00907_));
 sg13g2_inv_1 _20737_ (.Y(_03436_),
    .A(\cpu.ex.r_8[5] ));
 sg13g2_nand2_1 _20738_ (.Y(_03437_),
    .A(net643),
    .B(net590));
 sg13g2_o21ai_1 _20739_ (.B1(_03437_),
    .Y(_00908_),
    .A1(_03436_),
    .A2(net522));
 sg13g2_mux2_1 _20740_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net840),
    .S(net590),
    .X(_00909_));
 sg13g2_mux2_1 _20741_ (.A0(\cpu.ex.r_8[7] ),
    .A1(net716),
    .S(net590),
    .X(_00910_));
 sg13g2_mux2_1 _20742_ (.A0(\cpu.ex.r_8[8] ),
    .A1(net715),
    .S(_03431_),
    .X(_00911_));
 sg13g2_mux2_1 _20743_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net839),
    .S(_03431_),
    .X(_00912_));
 sg13g2_nor2_1 _20744_ (.A(_03382_),
    .B(_03411_),
    .Y(_03438_));
 sg13g2_buf_1 _20745_ (.A(_03438_),
    .X(_03439_));
 sg13g2_buf_1 _20746_ (.A(net589),
    .X(_03440_));
 sg13g2_mux2_1 _20747_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net718),
    .S(_03440_),
    .X(_00913_));
 sg13g2_mux2_1 _20748_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net838),
    .S(net521),
    .X(_00914_));
 sg13g2_inv_1 _20749_ (.Y(_03441_),
    .A(\cpu.ex.r_9[11] ));
 sg13g2_nand2_1 _20750_ (.Y(_03442_),
    .A(net950),
    .B(net589));
 sg13g2_o21ai_1 _20751_ (.B1(_03442_),
    .Y(_00915_),
    .A1(_03441_),
    .A2(_03440_));
 sg13g2_mux2_1 _20752_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net529),
    .S(net521),
    .X(_00916_));
 sg13g2_mux2_1 _20753_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net468),
    .S(net521),
    .X(_00917_));
 sg13g2_mux2_1 _20754_ (.A0(\cpu.ex.r_9[14] ),
    .A1(net524),
    .S(net521),
    .X(_00918_));
 sg13g2_mux2_1 _20755_ (.A0(\cpu.ex.r_9[15] ),
    .A1(net641),
    .S(net521),
    .X(_00919_));
 sg13g2_mux2_1 _20756_ (.A0(\cpu.ex.r_9[1] ),
    .A1(_09944_),
    .S(net521),
    .X(_00920_));
 sg13g2_mux2_1 _20757_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net406),
    .S(net521),
    .X(_00921_));
 sg13g2_mux2_1 _20758_ (.A0(\cpu.ex.r_9[3] ),
    .A1(_03396_),
    .S(net589),
    .X(_00922_));
 sg13g2_mux2_1 _20759_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net314),
    .S(net589),
    .X(_00923_));
 sg13g2_mux2_1 _20760_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net591),
    .S(net589),
    .X(_00924_));
 sg13g2_mux2_1 _20761_ (.A0(\cpu.ex.r_9[6] ),
    .A1(net840),
    .S(net589),
    .X(_00925_));
 sg13g2_mux2_1 _20762_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net716),
    .S(_03439_),
    .X(_00926_));
 sg13g2_mux2_1 _20763_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net715),
    .S(net589),
    .X(_00927_));
 sg13g2_nand2_1 _20764_ (.Y(_03443_),
    .A(net952),
    .B(net589));
 sg13g2_o21ai_1 _20765_ (.B1(_03443_),
    .Y(_00928_),
    .A1(_10628_),
    .A2(net521));
 sg13g2_inv_1 _20766_ (.Y(_03444_),
    .A(_11363_));
 sg13g2_nor2_1 _20767_ (.A(_08766_),
    .B(_03444_),
    .Y(_03445_));
 sg13g2_buf_1 _20768_ (.A(_03445_),
    .X(_03446_));
 sg13g2_nor2_1 _20769_ (.A(_11357_),
    .B(_03446_),
    .Y(_03447_));
 sg13g2_buf_2 _20770_ (.A(_03447_),
    .X(_03448_));
 sg13g2_inv_1 _20771_ (.Y(_03449_),
    .A(_00194_));
 sg13g2_nor2b_1 _20772_ (.A(_10601_),
    .B_N(_10618_),
    .Y(_03450_));
 sg13g2_buf_1 _20773_ (.A(_10351_),
    .X(_03451_));
 sg13g2_buf_1 _20774_ (.A(net313),
    .X(_03452_));
 sg13g2_buf_1 _20775_ (.A(net236),
    .X(_03453_));
 sg13g2_mux2_1 _20776_ (.A0(_03449_),
    .A1(_03450_),
    .S(net201),
    .X(_03454_));
 sg13g2_buf_2 _20777_ (.A(_03454_),
    .X(_03455_));
 sg13g2_buf_1 _20778_ (.A(_03455_),
    .X(_03456_));
 sg13g2_buf_1 _20779_ (.A(_10205_),
    .X(_03457_));
 sg13g2_nand2b_1 _20780_ (.Y(_03458_),
    .B(net235),
    .A_N(_10621_));
 sg13g2_o21ai_1 _20781_ (.B1(_03458_),
    .Y(_03459_),
    .A1(net235),
    .A2(_10573_));
 sg13g2_buf_1 _20782_ (.A(_03459_),
    .X(_03460_));
 sg13g2_buf_1 _20783_ (.A(net159),
    .X(_03461_));
 sg13g2_nor2_1 _20784_ (.A(_00289_),
    .B(net236),
    .Y(_03462_));
 sg13g2_nand2_1 _20785_ (.Y(_03463_),
    .A(net236),
    .B(_10546_));
 sg13g2_nand2b_1 _20786_ (.Y(_03464_),
    .B(_03463_),
    .A_N(_03462_));
 sg13g2_buf_1 _20787_ (.A(_03464_),
    .X(_03465_));
 sg13g2_nand2_1 _20788_ (.Y(_03466_),
    .A(_03452_),
    .B(_10599_));
 sg13g2_o21ai_1 _20789_ (.B1(_03466_),
    .Y(_03467_),
    .A1(_00196_),
    .A2(_03452_));
 sg13g2_buf_2 _20790_ (.A(_03467_),
    .X(_03468_));
 sg13g2_a21oi_1 _20791_ (.A1(net182),
    .A2(_03465_),
    .Y(_03469_),
    .B1(_03468_));
 sg13g2_nand3_1 _20792_ (.B(_03468_),
    .C(_03465_),
    .A(net182),
    .Y(_03470_));
 sg13g2_o21ai_1 _20793_ (.B1(_03470_),
    .Y(_03471_),
    .A1(net187),
    .A2(_03469_));
 sg13g2_buf_1 _20794_ (.A(_03471_),
    .X(_03472_));
 sg13g2_xnor2_1 _20795_ (.Y(_03473_),
    .A(_11295_),
    .B(_03468_));
 sg13g2_buf_1 _20796_ (.A(_03473_),
    .X(_03474_));
 sg13g2_nor2b_1 _20797_ (.A(_03462_),
    .B_N(_03463_),
    .Y(_03475_));
 sg13g2_buf_1 _20798_ (.A(_03475_),
    .X(_03476_));
 sg13g2_xnor2_1 _20799_ (.Y(_03477_),
    .A(_11177_),
    .B(net158));
 sg13g2_nor2_1 _20800_ (.A(net120),
    .B(_03477_),
    .Y(_03478_));
 sg13g2_inv_1 _20801_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_nor2b_1 _20802_ (.A(_10677_),
    .B_N(_10692_),
    .Y(_03480_));
 sg13g2_nor2_1 _20803_ (.A(_10676_),
    .B(net236),
    .Y(_03481_));
 sg13g2_a21oi_1 _20804_ (.A1(net236),
    .A2(_03480_),
    .Y(_03482_),
    .B1(_03481_));
 sg13g2_buf_2 _20805_ (.A(_03482_),
    .X(_03483_));
 sg13g2_inv_1 _20806_ (.Y(_03484_),
    .A(_03483_));
 sg13g2_buf_1 _20807_ (.A(_03484_),
    .X(_03485_));
 sg13g2_nand2b_1 _20808_ (.Y(_03486_),
    .B(net235),
    .A_N(_10695_));
 sg13g2_o21ai_1 _20809_ (.B1(_03486_),
    .Y(_03487_),
    .A1(net235),
    .A2(_10715_));
 sg13g2_buf_1 _20810_ (.A(_03487_),
    .X(_03488_));
 sg13g2_or2_1 _20811_ (.X(_03489_),
    .B(_10285_),
    .A(_10222_));
 sg13g2_mux2_1 _20812_ (.A0(_00191_),
    .A1(_03489_),
    .S(net313),
    .X(_03490_));
 sg13g2_buf_1 _20813_ (.A(_03490_),
    .X(_03491_));
 sg13g2_o21ai_1 _20814_ (.B1(_10805_),
    .Y(_03492_),
    .A1(_10488_),
    .A2(_10490_));
 sg13g2_buf_1 _20815_ (.A(_03492_),
    .X(_03493_));
 sg13g2_nand3_1 _20816_ (.B(net200),
    .C(_03493_),
    .A(net341),
    .Y(_03494_));
 sg13g2_mux2_1 _20817_ (.A0(_10394_),
    .A1(_11669_),
    .S(_03451_),
    .X(_03495_));
 sg13g2_buf_1 _20818_ (.A(_03495_),
    .X(_03496_));
 sg13g2_nand4_1 _20819_ (.B(_03496_),
    .C(net200),
    .A(net317),
    .Y(_03497_),
    .D(_03493_));
 sg13g2_buf_1 _20820_ (.A(_03496_),
    .X(_03498_));
 sg13g2_nor2_1 _20821_ (.A(net340),
    .B(_10850_),
    .Y(_03499_));
 sg13g2_buf_2 _20822_ (.A(_03499_),
    .X(_03500_));
 sg13g2_nand3_1 _20823_ (.B(_03493_),
    .C(_03500_),
    .A(net180),
    .Y(_03501_));
 sg13g2_nand3_1 _20824_ (.B(_03497_),
    .C(_03501_),
    .A(_03494_),
    .Y(_03502_));
 sg13g2_or2_1 _20825_ (.X(_03503_),
    .B(_10490_),
    .A(_10488_));
 sg13g2_buf_1 _20826_ (.A(_03503_),
    .X(_03504_));
 sg13g2_buf_1 _20827_ (.A(_03504_),
    .X(_03505_));
 sg13g2_nand2_1 _20828_ (.Y(_03506_),
    .A(net317),
    .B(net200));
 sg13g2_nand2_1 _20829_ (.Y(_03507_),
    .A(net180),
    .B(net200));
 sg13g2_nand2_1 _20830_ (.Y(_03508_),
    .A(_08738_),
    .B(_10176_));
 sg13g2_a21o_1 _20831_ (.A2(_10181_),
    .A1(net379),
    .B1(_03508_),
    .X(_03509_));
 sg13g2_buf_2 _20832_ (.A(_03509_),
    .X(_03510_));
 sg13g2_nor2_1 _20833_ (.A(_10327_),
    .B(_10347_),
    .Y(_03511_));
 sg13g2_nand3_1 _20834_ (.B(_10188_),
    .C(_10200_),
    .A(_10187_),
    .Y(_03512_));
 sg13g2_nor4_1 _20835_ (.A(_08834_),
    .B(_03512_),
    .C(_10327_),
    .D(_10347_),
    .Y(_03513_));
 sg13g2_a22oi_1 _20836_ (.Y(_03514_),
    .B1(_03513_),
    .B2(_09026_),
    .A2(_03511_),
    .A1(_10203_));
 sg13g2_buf_1 _20837_ (.A(_03514_),
    .X(_03515_));
 sg13g2_and2_1 _20838_ (.A(_03510_),
    .B(_03515_),
    .X(_03516_));
 sg13g2_buf_2 _20839_ (.A(_03516_),
    .X(_03517_));
 sg13g2_nor2_1 _20840_ (.A(_10918_),
    .B(_10947_),
    .Y(_03518_));
 sg13g2_a21o_1 _20841_ (.A2(_10323_),
    .A1(_10298_),
    .B1(_10324_),
    .X(_03519_));
 sg13g2_buf_1 _20842_ (.A(_03519_),
    .X(_03520_));
 sg13g2_mux2_1 _20843_ (.A0(_10206_),
    .A1(_03520_),
    .S(net313),
    .X(_03521_));
 sg13g2_and3_1 _20844_ (.X(_03522_),
    .A(_03510_),
    .B(_11331_),
    .C(_03515_));
 sg13g2_a221oi_1 _20845_ (.B2(net426),
    .C1(_10325_),
    .B1(net427),
    .A1(net1056),
    .Y(_03523_),
    .A2(net1009));
 sg13g2_a221oi_1 _20846_ (.B2(net426),
    .C1(_10207_),
    .B1(net427),
    .A1(net1056),
    .Y(_03524_),
    .A2(net1009));
 sg13g2_mux2_1 _20847_ (.A0(_03523_),
    .A1(_03524_),
    .S(_10205_),
    .X(_03525_));
 sg13g2_a221oi_1 _20848_ (.B2(_03522_),
    .C1(_03525_),
    .B1(_03521_),
    .A1(_03517_),
    .Y(_03526_),
    .A2(_03518_));
 sg13g2_buf_2 _20849_ (.A(_03526_),
    .X(_03527_));
 sg13g2_a221oi_1 _20850_ (.B2(_03507_),
    .C1(_03527_),
    .B1(_03506_),
    .A1(net322),
    .Y(_03528_),
    .A2(net199));
 sg13g2_nand2_1 _20851_ (.Y(_03529_),
    .A(_03493_),
    .B(_03500_));
 sg13g2_nand3_1 _20852_ (.B(net180),
    .C(_03493_),
    .A(net341),
    .Y(_03530_));
 sg13g2_a21oi_1 _20853_ (.A1(_03529_),
    .A2(_03530_),
    .Y(_03531_),
    .B1(_03527_));
 sg13g2_or3_1 _20854_ (.A(_03502_),
    .B(_03528_),
    .C(_03531_),
    .X(_03532_));
 sg13g2_mux2_1 _20855_ (.A0(_10398_),
    .A1(_10430_),
    .S(net313),
    .X(_03533_));
 sg13g2_buf_1 _20856_ (.A(_03533_),
    .X(_03534_));
 sg13g2_nor2_1 _20857_ (.A(_03534_),
    .B(_11042_),
    .Y(_03535_));
 sg13g2_nand2b_1 _20858_ (.Y(_03536_),
    .B(net321),
    .A_N(net247));
 sg13g2_nor2_1 _20859_ (.A(_10203_),
    .B(_10399_),
    .Y(_03537_));
 sg13g2_nand2_1 _20860_ (.Y(_03538_),
    .A(net379),
    .B(_10202_));
 sg13g2_a221oi_1 _20861_ (.B2(_03538_),
    .C1(_10801_),
    .B1(_03537_),
    .A1(net236),
    .Y(_03539_),
    .A2(_10456_));
 sg13g2_a21o_1 _20862_ (.A2(_10999_),
    .A1(net247),
    .B1(_03539_),
    .X(_03540_));
 sg13g2_a22oi_1 _20863_ (.Y(_03541_),
    .B1(_03536_),
    .B2(_03540_),
    .A2(_11042_),
    .A1(_03534_));
 sg13g2_nand2_1 _20864_ (.Y(_03542_),
    .A(_10798_),
    .B(_10492_));
 sg13g2_o21ai_1 _20865_ (.B1(_03542_),
    .Y(_03543_),
    .A1(_03535_),
    .A2(_03541_));
 sg13g2_nand2b_1 _20866_ (.Y(_03544_),
    .B(net313),
    .A_N(_10430_));
 sg13g2_o21ai_1 _20867_ (.B1(_03544_),
    .Y(_03545_),
    .A1(_10398_),
    .A2(net236));
 sg13g2_buf_1 _20868_ (.A(_03545_),
    .X(_03546_));
 sg13g2_a22oi_1 _20869_ (.Y(_03547_),
    .B1(_03537_),
    .B2(_03538_),
    .A2(_10456_),
    .A1(net313));
 sg13g2_buf_1 _20870_ (.A(_03547_),
    .X(_03548_));
 sg13g2_buf_1 _20871_ (.A(_03548_),
    .X(_03549_));
 sg13g2_o21ai_1 _20872_ (.B1(_03536_),
    .Y(_03550_),
    .A1(_11442_),
    .A2(net178));
 sg13g2_a221oi_1 _20873_ (.B2(_03550_),
    .C1(net211),
    .B1(_03541_),
    .A1(net179),
    .Y(_03551_),
    .A2(_10976_));
 sg13g2_o21ai_1 _20874_ (.B1(_03551_),
    .Y(_03552_),
    .A1(_03532_),
    .A2(_03543_));
 sg13g2_inv_1 _20875_ (.Y(_03553_),
    .A(_10675_));
 sg13g2_nor2_1 _20876_ (.A(_10651_),
    .B(net236),
    .Y(_03554_));
 sg13g2_a21o_1 _20877_ (.A2(_03553_),
    .A1(net201),
    .B1(_03554_),
    .X(_03555_));
 sg13g2_buf_1 _20878_ (.A(_03555_),
    .X(_03556_));
 sg13g2_nand2_1 _20879_ (.Y(_03557_),
    .A(net319),
    .B(_03556_));
 sg13g2_nand2_1 _20880_ (.Y(_03558_),
    .A(net186),
    .B(_03557_));
 sg13g2_buf_1 _20881_ (.A(_10647_),
    .X(_03559_));
 sg13g2_nand2_1 _20882_ (.Y(_03560_),
    .A(net198),
    .B(_03557_));
 sg13g2_nor2_1 _20883_ (.A(_03535_),
    .B(_03550_),
    .Y(_03561_));
 sg13g2_nor2_1 _20884_ (.A(_11003_),
    .B(_03504_),
    .Y(_03562_));
 sg13g2_nand2_1 _20885_ (.Y(_03563_),
    .A(net341),
    .B(net317));
 sg13g2_buf_1 _20886_ (.A(_03563_),
    .X(_03564_));
 sg13g2_a221oi_1 _20887_ (.B2(_03564_),
    .C1(_03527_),
    .B1(_03506_),
    .A1(net322),
    .Y(_03565_),
    .A2(_03504_));
 sg13g2_nand2b_1 _20888_ (.Y(_03566_),
    .B(_03451_),
    .A_N(_11669_));
 sg13g2_o21ai_1 _20889_ (.B1(_03566_),
    .Y(_03567_),
    .A1(_10394_),
    .A2(net313));
 sg13g2_buf_1 _20890_ (.A(_03567_),
    .X(_03568_));
 sg13g2_o21ai_1 _20891_ (.B1(_03493_),
    .Y(_03569_),
    .A1(_10883_),
    .A2(net200));
 sg13g2_nor3_1 _20892_ (.A(_03568_),
    .B(_03527_),
    .C(_03569_),
    .Y(_03570_));
 sg13g2_or4_1 _20893_ (.A(_03562_),
    .B(_03502_),
    .C(_03565_),
    .D(_03570_),
    .X(_03571_));
 sg13g2_buf_2 _20894_ (.A(_03571_),
    .X(_03572_));
 sg13g2_nor2_1 _20895_ (.A(_03535_),
    .B(_03541_),
    .Y(_03573_));
 sg13g2_a221oi_1 _20896_ (.B2(_03572_),
    .C1(_03573_),
    .B1(_03561_),
    .A1(_11075_),
    .Y(_03574_),
    .A2(_11093_));
 sg13g2_buf_1 _20897_ (.A(_03574_),
    .X(_03575_));
 sg13g2_a221oi_1 _20898_ (.B2(_03560_),
    .C1(_03575_),
    .B1(_03558_),
    .A1(_03488_),
    .Y(_03576_),
    .A2(_03552_));
 sg13g2_buf_1 _20899_ (.A(_03576_),
    .X(_03577_));
 sg13g2_buf_1 _20900_ (.A(_03556_),
    .X(_03578_));
 sg13g2_nand2_1 _20901_ (.Y(_03579_),
    .A(net198),
    .B(net186));
 sg13g2_nand2b_1 _20902_ (.Y(_03580_),
    .B(_03557_),
    .A_N(_03579_));
 sg13g2_o21ai_1 _20903_ (.B1(_03580_),
    .Y(_03581_),
    .A1(net319),
    .A2(net140));
 sg13g2_buf_1 _20904_ (.A(_03581_),
    .X(_03582_));
 sg13g2_nor2_1 _20905_ (.A(_03577_),
    .B(_03582_),
    .Y(_03583_));
 sg13g2_buf_1 _20906_ (.A(_03583_),
    .X(_03584_));
 sg13g2_nor2_1 _20907_ (.A(net119),
    .B(_03584_),
    .Y(_03585_));
 sg13g2_a21oi_1 _20908_ (.A1(net119),
    .A2(_03584_),
    .Y(_03586_),
    .B1(_11139_));
 sg13g2_nor3_1 _20909_ (.A(_03479_),
    .B(_03585_),
    .C(_03586_),
    .Y(_03587_));
 sg13g2_or2_1 _20910_ (.X(_03588_),
    .B(_03587_),
    .A(_03472_));
 sg13g2_mux2_1 _20911_ (.A0(_10621_),
    .A1(_10573_),
    .S(net201),
    .X(_03589_));
 sg13g2_buf_1 _20912_ (.A(_03589_),
    .X(_03590_));
 sg13g2_buf_1 _20913_ (.A(_03590_),
    .X(_03591_));
 sg13g2_buf_1 _20914_ (.A(_03483_),
    .X(_03592_));
 sg13g2_nor4_1 _20915_ (.A(net138),
    .B(_03479_),
    .C(_03577_),
    .D(_03582_),
    .Y(_03593_));
 sg13g2_nor4_1 _20916_ (.A(net208),
    .B(_03479_),
    .C(_03577_),
    .D(_03582_),
    .Y(_03594_));
 sg13g2_nor2_1 _20917_ (.A(_10169_),
    .B(net138),
    .Y(_03595_));
 sg13g2_and2_1 _20918_ (.A(_03478_),
    .B(_03595_),
    .X(_03596_));
 sg13g2_nor4_2 _20919_ (.A(_03472_),
    .B(_03593_),
    .C(_03594_),
    .Y(_03597_),
    .D(_03596_));
 sg13g2_a21oi_1 _20920_ (.A1(net139),
    .A2(_03597_),
    .Y(_03598_),
    .B1(net163));
 sg13g2_a221oi_1 _20921_ (.B2(_03588_),
    .C1(_03598_),
    .B1(_03461_),
    .A1(net188),
    .Y(_03599_),
    .A2(_03456_));
 sg13g2_o21ai_1 _20922_ (.B1(net901),
    .Y(_03600_),
    .A1(net188),
    .A2(_03456_));
 sg13g2_nor2_1 _20923_ (.A(_03457_),
    .B(_10619_),
    .Y(_03601_));
 sg13g2_a21oi_1 _20924_ (.A1(_03449_),
    .A2(_03457_),
    .Y(_03602_),
    .B1(_03601_));
 sg13g2_buf_1 _20925_ (.A(_03602_),
    .X(_03603_));
 sg13g2_nand2_1 _20926_ (.Y(_03604_),
    .A(net188),
    .B(net157));
 sg13g2_inv_1 _20927_ (.Y(_03605_),
    .A(_03604_));
 sg13g2_nor2_2 _20928_ (.A(net162),
    .B(net139),
    .Y(_03606_));
 sg13g2_nor2_1 _20929_ (.A(net163),
    .B(net159),
    .Y(_03607_));
 sg13g2_buf_1 _20930_ (.A(_03468_),
    .X(_03608_));
 sg13g2_or2_1 _20931_ (.X(_03609_),
    .B(net137),
    .A(net187));
 sg13g2_inv_1 _20932_ (.Y(_03610_),
    .A(_03609_));
 sg13g2_nand4_1 _20933_ (.B(_10848_),
    .C(_10354_),
    .A(_10813_),
    .Y(_03611_),
    .D(_10392_));
 sg13g2_nand3b_1 _20934_ (.B(_10813_),
    .C(_10848_),
    .Y(_03612_),
    .A_N(_10394_));
 sg13g2_mux2_1 _20935_ (.A0(_03611_),
    .A1(_03612_),
    .S(net235),
    .X(_03613_));
 sg13g2_buf_1 _20936_ (.A(_03613_),
    .X(_03614_));
 sg13g2_nor2_1 _20937_ (.A(net200),
    .B(_03614_),
    .Y(_03615_));
 sg13g2_a21oi_1 _20938_ (.A1(_03491_),
    .A2(_03614_),
    .Y(_03616_),
    .B1(net340));
 sg13g2_nand2_1 _20939_ (.Y(_03617_),
    .A(_11003_),
    .B(_10492_));
 sg13g2_o21ai_1 _20940_ (.B1(_03617_),
    .Y(_03618_),
    .A1(_03615_),
    .A2(_03616_));
 sg13g2_a221oi_1 _20941_ (.B2(_03510_),
    .C1(_10918_),
    .B1(_03515_),
    .A1(_10925_),
    .Y(_03619_),
    .A2(_10945_));
 sg13g2_a221oi_1 _20942_ (.B2(net426),
    .C1(_03520_),
    .B1(net427),
    .A1(net1056),
    .Y(_03620_),
    .A2(net1009));
 sg13g2_a221oi_1 _20943_ (.B2(net426),
    .C1(_10206_),
    .B1(net427),
    .A1(net1056),
    .Y(_03621_),
    .A2(net1009));
 sg13g2_mux2_1 _20944_ (.A0(_03620_),
    .A1(_03621_),
    .S(net235),
    .X(_03622_));
 sg13g2_buf_1 _20945_ (.A(_03622_),
    .X(_03623_));
 sg13g2_a21o_1 _20946_ (.A2(_10945_),
    .A1(_10925_),
    .B1(_03520_),
    .X(_03624_));
 sg13g2_a221oi_1 _20947_ (.B2(_03510_),
    .C1(_03624_),
    .B1(_11672_),
    .A1(_10176_),
    .Y(_03625_),
    .A2(_03538_));
 sg13g2_nor4_1 _20948_ (.A(_10206_),
    .B(_03510_),
    .C(net313),
    .D(_10947_),
    .Y(_03626_));
 sg13g2_or4_1 _20949_ (.A(_03619_),
    .B(_03623_),
    .C(_03625_),
    .D(_03626_),
    .X(_03627_));
 sg13g2_buf_1 _20950_ (.A(_03627_),
    .X(_03628_));
 sg13g2_nor3_1 _20951_ (.A(_10798_),
    .B(_10488_),
    .C(_10490_),
    .Y(_03629_));
 sg13g2_a221oi_1 _20952_ (.B2(net340),
    .C1(_03629_),
    .B1(net200),
    .A1(_10850_),
    .Y(_03630_),
    .A2(net180));
 sg13g2_nor2_1 _20953_ (.A(net322),
    .B(_10492_),
    .Y(_03631_));
 sg13g2_a21oi_1 _20954_ (.A1(_03628_),
    .A2(_03630_),
    .Y(_03632_),
    .B1(_03631_));
 sg13g2_nor2_2 _20955_ (.A(_10801_),
    .B(_03548_),
    .Y(_03633_));
 sg13g2_nor2_2 _20956_ (.A(net247),
    .B(net321),
    .Y(_03634_));
 sg13g2_nand2_1 _20957_ (.Y(_03635_),
    .A(net247),
    .B(net321));
 sg13g2_o21ai_1 _20958_ (.B1(_03635_),
    .Y(_03636_),
    .A1(_03633_),
    .A2(_03634_));
 sg13g2_nand2_1 _20959_ (.Y(_03637_),
    .A(net179),
    .B(_11488_));
 sg13g2_nand4_1 _20960_ (.B(_03632_),
    .C(_03636_),
    .A(_03618_),
    .Y(_03638_),
    .D(_03637_));
 sg13g2_nor2_1 _20961_ (.A(net179),
    .B(net184),
    .Y(_03639_));
 sg13g2_a22oi_1 _20962_ (.Y(_03640_),
    .B1(net321),
    .B2(net247),
    .A2(_03548_),
    .A1(net243));
 sg13g2_nor2_1 _20963_ (.A(_03634_),
    .B(_03640_),
    .Y(_03641_));
 sg13g2_o21ai_1 _20964_ (.B1(_03637_),
    .Y(_03642_),
    .A1(_03639_),
    .A2(_03641_));
 sg13g2_nand2b_1 _20965_ (.Y(_03643_),
    .B(net235),
    .A_N(_10626_));
 sg13g2_o21ai_1 _20966_ (.B1(_03643_),
    .Y(_03644_),
    .A1(net235),
    .A2(_10645_));
 sg13g2_buf_2 _20967_ (.A(_03644_),
    .X(_03645_));
 sg13g2_nand2_2 _20968_ (.Y(_03646_),
    .A(_03645_),
    .B(_11073_));
 sg13g2_nand2_1 _20969_ (.Y(_03647_),
    .A(net211),
    .B(_03646_));
 sg13g2_nand2_1 _20970_ (.Y(_03648_),
    .A(_10717_),
    .B(_03646_));
 sg13g2_a22oi_1 _20971_ (.Y(_03649_),
    .B1(_03647_),
    .B2(_03648_),
    .A2(_03642_),
    .A1(_03638_));
 sg13g2_buf_2 _20972_ (.A(_03649_),
    .X(_03650_));
 sg13g2_nand2_1 _20973_ (.Y(_03651_),
    .A(_03559_),
    .B(_11513_));
 sg13g2_nand3_1 _20974_ (.B(net211),
    .C(_03646_),
    .A(_10717_),
    .Y(_03652_));
 sg13g2_nand2_1 _20975_ (.Y(_03653_),
    .A(_03651_),
    .B(_03652_));
 sg13g2_buf_1 _20976_ (.A(_03465_),
    .X(_03654_));
 sg13g2_nor2_2 _20977_ (.A(_11139_),
    .B(_03483_),
    .Y(_03655_));
 sg13g2_nor3_1 _20978_ (.A(net140),
    .B(net136),
    .C(_03655_),
    .Y(_03656_));
 sg13g2_o21ai_1 _20979_ (.B1(_03656_),
    .Y(_03657_),
    .A1(_03650_),
    .A2(_03653_));
 sg13g2_nor3_1 _20980_ (.A(net320),
    .B(net136),
    .C(_03655_),
    .Y(_03658_));
 sg13g2_o21ai_1 _20981_ (.B1(_03658_),
    .Y(_03659_),
    .A1(_03650_),
    .A2(_03653_));
 sg13g2_nor2_1 _20982_ (.A(_10169_),
    .B(_03484_),
    .Y(_03660_));
 sg13g2_buf_2 _20983_ (.A(_03660_),
    .X(_03661_));
 sg13g2_a21oi_1 _20984_ (.A1(net201),
    .A2(_03553_),
    .Y(_03662_),
    .B1(_03554_));
 sg13g2_buf_2 _20985_ (.A(_03662_),
    .X(_03663_));
 sg13g2_a22oi_1 _20986_ (.Y(_03664_),
    .B1(_03658_),
    .B2(_03663_),
    .A2(_03661_),
    .A1(net158));
 sg13g2_and3_1 _20987_ (.X(_03665_),
    .A(_03657_),
    .B(_03659_),
    .C(_03664_));
 sg13g2_buf_1 _20988_ (.A(_03665_),
    .X(_03666_));
 sg13g2_and2_1 _20989_ (.A(_03651_),
    .B(_03652_),
    .X(_03667_));
 sg13g2_nor3_1 _20990_ (.A(_03663_),
    .B(net158),
    .C(_03661_),
    .Y(_03668_));
 sg13g2_nand3b_1 _20991_ (.B(_03667_),
    .C(_03668_),
    .Y(_03669_),
    .A_N(_03650_));
 sg13g2_nor3_1 _20992_ (.A(net319),
    .B(net158),
    .C(_03661_),
    .Y(_03670_));
 sg13g2_nand3b_1 _20993_ (.B(_03667_),
    .C(_03670_),
    .Y(_03671_),
    .A_N(_03650_));
 sg13g2_a22oi_1 _20994_ (.Y(_03672_),
    .B1(_03670_),
    .B2(_03578_),
    .A2(_03655_),
    .A1(net136));
 sg13g2_nand4_1 _20995_ (.B(_03669_),
    .C(_03671_),
    .A(_11572_),
    .Y(_03673_),
    .D(_03672_));
 sg13g2_buf_1 _20996_ (.A(_03673_),
    .X(_03674_));
 sg13g2_and2_1 _20997_ (.A(net187),
    .B(_03468_),
    .X(_03675_));
 sg13g2_buf_1 _20998_ (.A(_03675_),
    .X(_03676_));
 sg13g2_a21oi_1 _20999_ (.A1(_03666_),
    .A2(_03674_),
    .Y(_03677_),
    .B1(_03676_));
 sg13g2_nor3_1 _21000_ (.A(_03607_),
    .B(_03610_),
    .C(_03677_),
    .Y(_03678_));
 sg13g2_nor2_1 _21001_ (.A(_03606_),
    .B(_03678_),
    .Y(_03679_));
 sg13g2_nor2_1 _21002_ (.A(net188),
    .B(net157),
    .Y(_03680_));
 sg13g2_nor2_1 _21003_ (.A(net901),
    .B(_03680_),
    .Y(_03681_));
 sg13g2_o21ai_1 _21004_ (.B1(_03681_),
    .Y(_03682_),
    .A1(_03605_),
    .A2(_03679_));
 sg13g2_o21ai_1 _21005_ (.B1(_03682_),
    .Y(_03683_),
    .A1(_03599_),
    .A2(_03600_));
 sg13g2_nand2_1 _21006_ (.Y(_03684_),
    .A(\cpu.ex.r_cc ),
    .B(_03448_));
 sg13g2_o21ai_1 _21007_ (.B1(_03684_),
    .Y(_00929_),
    .A1(_03448_),
    .A2(_03683_));
 sg13g2_nor2_1 _21008_ (.A(net1096),
    .B(_10057_),
    .Y(_03685_));
 sg13g2_nand4_1 _21009_ (.B(net1010),
    .C(net1097),
    .A(net1011),
    .Y(_03686_),
    .D(_03685_));
 sg13g2_nand2b_1 _21010_ (.Y(_03687_),
    .B(_08738_),
    .A_N(_03686_));
 sg13g2_buf_1 _21011_ (.A(_03687_),
    .X(_03688_));
 sg13g2_buf_1 _21012_ (.A(_03688_),
    .X(_03689_));
 sg13g2_buf_1 _21013_ (.A(_03688_),
    .X(_03690_));
 sg13g2_nand2_1 _21014_ (.Y(_03691_),
    .A(\cpu.ex.r_epc[1] ),
    .B(net587));
 sg13g2_o21ai_1 _21015_ (.B1(_03691_),
    .Y(_00931_),
    .A1(_09976_),
    .A2(net588));
 sg13g2_mux2_1 _21016_ (.A0(net848),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net588),
    .X(_00932_));
 sg13g2_buf_1 _21017_ (.A(_08822_),
    .X(_03692_));
 sg13g2_buf_1 _21018_ (.A(_03692_),
    .X(_03693_));
 sg13g2_nand2_1 _21019_ (.Y(_03694_),
    .A(\cpu.ex.r_epc[12] ),
    .B(net587));
 sg13g2_o21ai_1 _21020_ (.B1(_03694_),
    .Y(_00933_),
    .A1(net640),
    .A2(net588));
 sg13g2_buf_1 _21021_ (.A(net528),
    .X(_03695_));
 sg13g2_mux2_1 _21022_ (.A0(net467),
    .A1(\cpu.ex.r_epc[13] ),
    .S(net588),
    .X(_00934_));
 sg13g2_buf_1 _21023_ (.A(net594),
    .X(_03696_));
 sg13g2_mux2_1 _21024_ (.A0(net520),
    .A1(\cpu.ex.r_epc[14] ),
    .S(net588),
    .X(_00935_));
 sg13g2_buf_1 _21025_ (.A(net717),
    .X(_03697_));
 sg13g2_mux2_1 _21026_ (.A0(net639),
    .A1(\cpu.ex.r_epc[15] ),
    .S(net588),
    .X(_00936_));
 sg13g2_buf_1 _21027_ (.A(net892),
    .X(_03698_));
 sg13g2_buf_2 _21028_ (.A(net713),
    .X(_03699_));
 sg13g2_nand2_1 _21029_ (.Y(_03700_),
    .A(\cpu.ex.r_epc[2] ),
    .B(net587));
 sg13g2_o21ai_1 _21030_ (.B1(_03700_),
    .Y(_00937_),
    .A1(net638),
    .A2(net588));
 sg13g2_nand2_1 _21031_ (.Y(_03701_),
    .A(\cpu.ex.r_epc[3] ),
    .B(net587));
 sg13g2_o21ai_1 _21032_ (.B1(_03701_),
    .Y(_00938_),
    .A1(net780),
    .A2(net588));
 sg13g2_buf_1 _21033_ (.A(net891),
    .X(_03702_));
 sg13g2_buf_1 _21034_ (.A(net712),
    .X(_03703_));
 sg13g2_buf_1 _21035_ (.A(net637),
    .X(_03704_));
 sg13g2_nand2_1 _21036_ (.Y(_03705_),
    .A(\cpu.ex.r_epc[4] ),
    .B(net587));
 sg13g2_o21ai_1 _21037_ (.B1(_03705_),
    .Y(_00939_),
    .A1(net586),
    .A2(_03689_));
 sg13g2_nand2_1 _21038_ (.Y(_03706_),
    .A(\cpu.ex.r_epc[5] ),
    .B(_03688_));
 sg13g2_o21ai_1 _21039_ (.B1(_03706_),
    .Y(_00940_),
    .A1(net729),
    .A2(_03689_));
 sg13g2_mux2_1 _21040_ (.A0(net728),
    .A1(\cpu.ex.r_epc[6] ),
    .S(_03690_),
    .X(_00941_));
 sg13g2_mux2_1 _21041_ (.A0(net727),
    .A1(\cpu.ex.r_epc[7] ),
    .S(net587),
    .X(_00942_));
 sg13g2_mux2_1 _21042_ (.A0(net726),
    .A1(\cpu.ex.r_epc[8] ),
    .S(_03690_),
    .X(_00943_));
 sg13g2_mux2_1 _21043_ (.A0(net850),
    .A1(\cpu.ex.r_epc[9] ),
    .S(net587),
    .X(_00944_));
 sg13g2_mux2_1 _21044_ (.A0(net849),
    .A1(\cpu.ex.r_epc[10] ),
    .S(net587),
    .X(_00945_));
 sg13g2_nand4_1 _21045_ (.B(net1010),
    .C(net1097),
    .A(_03410_),
    .Y(_03707_),
    .D(_03685_));
 sg13g2_buf_1 _21046_ (.A(_03707_),
    .X(_03708_));
 sg13g2_buf_1 _21047_ (.A(_03708_),
    .X(_03709_));
 sg13g2_buf_1 _21048_ (.A(_03708_),
    .X(_03710_));
 sg13g2_nand2_1 _21049_ (.Y(_03711_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net584));
 sg13g2_o21ai_1 _21050_ (.B1(_03711_),
    .Y(_00951_),
    .A1(_09976_),
    .A2(net585));
 sg13g2_mux2_1 _21051_ (.A0(net848),
    .A1(\cpu.ex.r_lr[11] ),
    .S(net585),
    .X(_00952_));
 sg13g2_nand2_1 _21052_ (.Y(_03712_),
    .A(\cpu.ex.r_lr[12] ),
    .B(net584));
 sg13g2_o21ai_1 _21053_ (.B1(_03712_),
    .Y(_00953_),
    .A1(net640),
    .A2(net585));
 sg13g2_mux2_1 _21054_ (.A0(net467),
    .A1(\cpu.ex.r_lr[13] ),
    .S(net585),
    .X(_00954_));
 sg13g2_mux2_1 _21055_ (.A0(net520),
    .A1(\cpu.ex.r_lr[14] ),
    .S(_03709_),
    .X(_00955_));
 sg13g2_mux2_1 _21056_ (.A0(net639),
    .A1(\cpu.ex.r_lr[15] ),
    .S(_03709_),
    .X(_00956_));
 sg13g2_nand2_1 _21057_ (.Y(_03713_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net584));
 sg13g2_o21ai_1 _21058_ (.B1(_03713_),
    .Y(_00957_),
    .A1(net638),
    .A2(net585));
 sg13g2_nand2_1 _21059_ (.Y(_03714_),
    .A(\cpu.ex.r_lr[3] ),
    .B(_03710_));
 sg13g2_o21ai_1 _21060_ (.B1(_03714_),
    .Y(_00958_),
    .A1(net780),
    .A2(net585));
 sg13g2_nand2_1 _21061_ (.Y(_03715_),
    .A(\cpu.ex.r_lr[4] ),
    .B(net584));
 sg13g2_o21ai_1 _21062_ (.B1(_03715_),
    .Y(_00959_),
    .A1(net586),
    .A2(net585));
 sg13g2_nand2_1 _21063_ (.Y(_03716_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03708_));
 sg13g2_o21ai_1 _21064_ (.B1(_03716_),
    .Y(_00960_),
    .A1(net729),
    .A2(net585));
 sg13g2_mux2_1 _21065_ (.A0(net728),
    .A1(\cpu.ex.r_lr[6] ),
    .S(_03710_),
    .X(_00961_));
 sg13g2_mux2_1 _21066_ (.A0(net727),
    .A1(\cpu.ex.r_lr[7] ),
    .S(net584),
    .X(_00962_));
 sg13g2_mux2_1 _21067_ (.A0(net726),
    .A1(\cpu.ex.r_lr[8] ),
    .S(net584),
    .X(_00963_));
 sg13g2_mux2_1 _21068_ (.A0(net850),
    .A1(\cpu.ex.r_lr[9] ),
    .S(net584),
    .X(_00964_));
 sg13g2_mux2_1 _21069_ (.A0(net849),
    .A1(\cpu.ex.r_lr[10] ),
    .S(net584),
    .X(_00965_));
 sg13g2_nor2_2 _21070_ (.A(_09216_),
    .B(net604),
    .Y(_03717_));
 sg13g2_nand2_1 _21071_ (.Y(_03718_),
    .A(net542),
    .B(_03717_));
 sg13g2_buf_1 _21072_ (.A(_03718_),
    .X(_03719_));
 sg13g2_inv_1 _21073_ (.Y(_03720_),
    .A(\cpu.ex.r_mult[15] ));
 sg13g2_inv_1 _21074_ (.Y(_03721_),
    .A(_11640_));
 sg13g2_a22oi_1 _21075_ (.Y(_03722_),
    .B1(_11640_),
    .B2(_11641_),
    .A2(_11622_),
    .A1(_11634_));
 sg13g2_a21oi_1 _21076_ (.A1(_11641_),
    .A2(_11205_),
    .Y(_03723_),
    .B1(_11239_));
 sg13g2_and4_1 _21077_ (.A(_11327_),
    .B(_11618_),
    .C(_11630_),
    .D(_03723_),
    .X(_03724_));
 sg13g2_or4_1 _21078_ (.A(_11634_),
    .B(_10524_),
    .C(_10650_),
    .D(_10720_),
    .X(_03725_));
 sg13g2_a221oi_1 _21079_ (.B2(_11641_),
    .C1(_03725_),
    .B1(_11640_),
    .A1(_11616_),
    .Y(_03726_),
    .A2(_11626_));
 sg13g2_nand2b_1 _21080_ (.Y(_03727_),
    .B(_11270_),
    .A_N(_11634_));
 sg13g2_or4_1 _21081_ (.A(_10524_),
    .B(_10650_),
    .C(_10720_),
    .D(_03727_),
    .X(_03728_));
 sg13g2_a21oi_1 _21082_ (.A1(_11641_),
    .A2(_11640_),
    .Y(_03729_),
    .B1(_03728_));
 sg13g2_or3_1 _21083_ (.A(_03724_),
    .B(_03726_),
    .C(_03729_),
    .X(_03730_));
 sg13g2_a221oi_1 _21084_ (.B2(_11621_),
    .C1(_03730_),
    .B1(_03722_),
    .A1(_11660_),
    .Y(_03731_),
    .A2(_03721_));
 sg13g2_buf_2 _21085_ (.A(_03731_),
    .X(_03732_));
 sg13g2_and2_1 _21086_ (.A(_03720_),
    .B(_03732_),
    .X(_03733_));
 sg13g2_nor2_1 _21087_ (.A(_03720_),
    .B(_03732_),
    .Y(_03734_));
 sg13g2_nor3_1 _21088_ (.A(_03719_),
    .B(_03733_),
    .C(_03734_),
    .Y(_03735_));
 sg13g2_nor2_1 _21089_ (.A(_11279_),
    .B(_11308_),
    .Y(_03736_));
 sg13g2_buf_8 _21090_ (.A(_03736_),
    .X(_03737_));
 sg13g2_o21ai_1 _21091_ (.B1(net88),
    .Y(_03738_),
    .A1(net245),
    .A2(_03737_));
 sg13g2_a21o_1 _21092_ (.A2(_11144_),
    .A1(_11137_),
    .B1(_11277_),
    .X(_03739_));
 sg13g2_inv_1 _21093_ (.Y(_03740_),
    .A(_11276_));
 sg13g2_a21oi_1 _21094_ (.A1(_11281_),
    .A2(_11289_),
    .Y(_03741_),
    .B1(_11292_));
 sg13g2_a221oi_1 _21095_ (.B2(_03741_),
    .C1(_11305_),
    .B1(_03740_),
    .A1(net539),
    .Y(_03742_),
    .A2(_11304_));
 sg13g2_nand2_1 _21096_ (.Y(_03743_),
    .A(_03739_),
    .B(_03742_));
 sg13g2_buf_8 _21097_ (.A(_03743_),
    .X(_03744_));
 sg13g2_nand3_1 _21098_ (.B(net244),
    .C(net28),
    .A(net87),
    .Y(_03745_));
 sg13g2_a21oi_1 _21099_ (.A1(_03738_),
    .A2(_03745_),
    .Y(_03746_),
    .B1(_11533_));
 sg13g2_inv_1 _21100_ (.Y(_03747_),
    .A(net1032));
 sg13g2_nor2_1 _21101_ (.A(_03747_),
    .B(_10061_),
    .Y(_03748_));
 sg13g2_nand3_1 _21102_ (.B(_10062_),
    .C(\cpu.ex.r_cc ),
    .A(_10055_),
    .Y(_03749_));
 sg13g2_and2_1 _21103_ (.A(_09207_),
    .B(_10067_),
    .X(_03750_));
 sg13g2_nand3_1 _21104_ (.B(_10064_),
    .C(_03750_),
    .A(\cpu.ex.r_mult[16] ),
    .Y(_03751_));
 sg13g2_inv_1 _21105_ (.Y(_03752_),
    .A(_10059_));
 sg13g2_nor3_1 _21106_ (.A(_10085_),
    .B(_03400_),
    .C(_03752_),
    .Y(_03753_));
 sg13g2_buf_1 _21107_ (.A(_03753_),
    .X(_03754_));
 sg13g2_buf_1 _21108_ (.A(net583),
    .X(_03755_));
 sg13g2_a21oi_1 _21109_ (.A1(_03749_),
    .A2(_03751_),
    .Y(_03756_),
    .B1(_03755_));
 sg13g2_or4_1 _21110_ (.A(_03735_),
    .B(_03746_),
    .C(_03748_),
    .D(_03756_),
    .X(_00966_));
 sg13g2_inv_1 _21111_ (.Y(_03757_),
    .A(\cpu.ex.r_mult[17] ));
 sg13g2_nor2_1 _21112_ (.A(net538),
    .B(_10068_),
    .Y(_03758_));
 sg13g2_buf_1 _21113_ (.A(_03758_),
    .X(_03759_));
 sg13g2_nor2_1 _21114_ (.A(net88),
    .B(net245),
    .Y(_03760_));
 sg13g2_xnor2_1 _21115_ (.Y(_03761_),
    .A(net318),
    .B(_03760_));
 sg13g2_o21ai_1 _21116_ (.B1(_03761_),
    .Y(_03762_),
    .A1(_11279_),
    .A2(_11308_));
 sg13g2_xnor2_1 _21117_ (.Y(_03763_),
    .A(_10887_),
    .B(_03762_));
 sg13g2_nand2_1 _21118_ (.Y(_03764_),
    .A(net61),
    .B(_03763_));
 sg13g2_xnor2_1 _21119_ (.Y(_03765_),
    .A(_00309_),
    .B(_03734_));
 sg13g2_nand2_2 _21120_ (.Y(_03766_),
    .A(_10064_),
    .B(_03750_));
 sg13g2_nand4_1 _21121_ (.B(_10055_),
    .C(_10062_),
    .A(_08842_),
    .Y(_03767_),
    .D(\cpu.ex.r_cc ));
 sg13g2_a21oi_1 _21122_ (.A1(_03766_),
    .A2(_03767_),
    .Y(_03768_),
    .B1(net583));
 sg13g2_buf_1 _21123_ (.A(_03768_),
    .X(_03769_));
 sg13g2_buf_1 _21124_ (.A(_03769_),
    .X(_03770_));
 sg13g2_a221oi_1 _21125_ (.B2(_03765_),
    .C1(net334),
    .B1(net338),
    .A1(net609),
    .Y(_03771_),
    .A2(net519));
 sg13g2_a22oi_1 _21126_ (.Y(_00967_),
    .B1(_03764_),
    .B2(_03771_),
    .A2(net404),
    .A1(_03757_));
 sg13g2_inv_1 _21127_ (.Y(_03772_),
    .A(\cpu.ex.r_mult[18] ));
 sg13g2_a21oi_1 _21128_ (.A1(net469),
    .A2(net519),
    .Y(_03773_),
    .B1(net334));
 sg13g2_nand2_1 _21129_ (.Y(_03774_),
    .A(_10887_),
    .B(_10918_));
 sg13g2_nand3_1 _21130_ (.B(net122),
    .C(_11331_),
    .A(_03774_),
    .Y(_03775_));
 sg13g2_buf_1 _21131_ (.A(_03775_),
    .X(_03776_));
 sg13g2_and2_1 _21132_ (.A(_11019_),
    .B(_03776_),
    .X(_03777_));
 sg13g2_xnor2_1 _21133_ (.Y(_03778_),
    .A(net209),
    .B(_03777_));
 sg13g2_a21oi_1 _21134_ (.A1(_03739_),
    .A2(_03742_),
    .Y(_03779_),
    .B1(_03778_));
 sg13g2_nand2_1 _21135_ (.Y(_03780_),
    .A(net539),
    .B(net77));
 sg13g2_or3_1 _21136_ (.A(_00309_),
    .B(_03720_),
    .C(_11372_),
    .X(_03781_));
 sg13g2_buf_1 _21137_ (.A(_03781_),
    .X(_03782_));
 sg13g2_o21ai_1 _21138_ (.B1(_03717_),
    .Y(_03783_),
    .A1(_03732_),
    .A2(_03782_));
 sg13g2_and2_1 _21139_ (.A(_10810_),
    .B(_03783_),
    .X(_03784_));
 sg13g2_o21ai_1 _21140_ (.B1(_03784_),
    .Y(_03785_),
    .A1(_03779_),
    .A2(_03780_));
 sg13g2_nor2_1 _21141_ (.A(_03732_),
    .B(_03782_),
    .Y(_03786_));
 sg13g2_buf_2 _21142_ (.A(_03786_),
    .X(_03787_));
 sg13g2_a21o_1 _21143_ (.A2(_03787_),
    .A1(_03717_),
    .B1(_10810_),
    .X(_03788_));
 sg13g2_a21o_1 _21144_ (.A2(_03779_),
    .A1(_11324_),
    .B1(_03788_),
    .X(_03789_));
 sg13g2_nand3_1 _21145_ (.B(_03785_),
    .C(_03789_),
    .A(net542),
    .Y(_03790_));
 sg13g2_a22oi_1 _21146_ (.Y(_00968_),
    .B1(_03773_),
    .B2(_03790_),
    .A2(net404),
    .A1(_03772_));
 sg13g2_inv_1 _21147_ (.Y(_03791_),
    .A(\cpu.ex.r_mult[19] ));
 sg13g2_nand3_1 _21148_ (.B(_11019_),
    .C(_03776_),
    .A(net209),
    .Y(_03792_));
 sg13g2_nand2_1 _21149_ (.Y(_03793_),
    .A(_10810_),
    .B(net606));
 sg13g2_a21oi_1 _21150_ (.A1(_11019_),
    .A2(_03776_),
    .Y(_03794_),
    .B1(net209));
 sg13g2_a21o_1 _21151_ (.A2(_03793_),
    .A1(_03792_),
    .B1(_03794_),
    .X(_03795_));
 sg13g2_xnor2_1 _21152_ (.Y(_03796_),
    .A(net316),
    .B(_03795_));
 sg13g2_a221oi_1 _21153_ (.B2(_03796_),
    .C1(_10851_),
    .B1(net28),
    .A1(_09202_),
    .Y(_03797_),
    .A2(net737));
 sg13g2_buf_1 _21154_ (.A(_10883_),
    .X(_03798_));
 sg13g2_xnor2_1 _21155_ (.Y(_03799_),
    .A(net312),
    .B(_03795_));
 sg13g2_nor3_1 _21156_ (.A(_11015_),
    .B(_03737_),
    .C(_03799_),
    .Y(_03800_));
 sg13g2_o21ai_1 _21157_ (.B1(net61),
    .Y(_03801_),
    .A1(_03797_),
    .A2(_03800_));
 sg13g2_nor2_1 _21158_ (.A(_10851_),
    .B(_10809_),
    .Y(_03802_));
 sg13g2_inv_1 _21159_ (.Y(_03803_),
    .A(_10851_));
 sg13g2_a21oi_1 _21160_ (.A1(_10810_),
    .A2(_03787_),
    .Y(_03804_),
    .B1(_03803_));
 sg13g2_a21oi_1 _21161_ (.A1(_03787_),
    .A2(_03802_),
    .Y(_03805_),
    .B1(_03804_));
 sg13g2_a221oi_1 _21162_ (.B2(_03805_),
    .C1(net334),
    .B1(net338),
    .A1(_03396_),
    .Y(_03806_),
    .A2(net519));
 sg13g2_a22oi_1 _21163_ (.Y(_00969_),
    .B1(_03801_),
    .B2(_03806_),
    .A2(net404),
    .A1(_03791_));
 sg13g2_nor2_1 _21164_ (.A(net1088),
    .B(net616),
    .Y(_03807_));
 sg13g2_buf_1 _21165_ (.A(_09213_),
    .X(_03808_));
 sg13g2_nor2_1 _21166_ (.A(net518),
    .B(_10885_),
    .Y(_03809_));
 sg13g2_nor2_1 _21167_ (.A(_03776_),
    .B(_03809_),
    .Y(_03810_));
 sg13g2_or2_1 _21168_ (.X(_03811_),
    .B(_03810_),
    .A(_11024_));
 sg13g2_xnor2_1 _21169_ (.Y(_03812_),
    .A(net322),
    .B(_03811_));
 sg13g2_o21ai_1 _21170_ (.B1(_03812_),
    .Y(_03813_),
    .A1(_11279_),
    .A2(_11308_));
 sg13g2_xnor2_1 _21171_ (.Y(_03814_),
    .A(_03807_),
    .B(_03813_));
 sg13g2_nand2_1 _21172_ (.Y(_03815_),
    .A(net77),
    .B(_03814_));
 sg13g2_nor2_1 _21173_ (.A(net1088),
    .B(net604),
    .Y(_03816_));
 sg13g2_nand2_1 _21174_ (.Y(_03817_),
    .A(_03787_),
    .B(_03802_));
 sg13g2_mux2_1 _21175_ (.A0(net1088),
    .A1(_03816_),
    .S(_03817_),
    .X(_03818_));
 sg13g2_a221oi_1 _21176_ (.B2(net1103),
    .C1(net334),
    .B1(_03818_),
    .A1(net366),
    .Y(_03819_),
    .A2(net519));
 sg13g2_nor2_1 _21177_ (.A(\cpu.ex.r_mult[20] ),
    .B(_03766_),
    .Y(_03820_));
 sg13g2_nor2_1 _21178_ (.A(_10064_),
    .B(_03769_),
    .Y(_03821_));
 sg13g2_o21ai_1 _21179_ (.B1(_10061_),
    .Y(_03822_),
    .A1(_03820_),
    .A2(_03821_));
 sg13g2_o21ai_1 _21180_ (.B1(_03822_),
    .Y(_03823_),
    .A1(net335),
    .A2(_10061_));
 sg13g2_a21oi_1 _21181_ (.A1(_03815_),
    .A2(_03819_),
    .Y(_00970_),
    .B1(_03823_));
 sg13g2_inv_1 _21182_ (.Y(_03824_),
    .A(\cpu.ex.r_mult[21] ));
 sg13g2_inv_1 _21183_ (.Y(_03825_),
    .A(_10807_));
 sg13g2_nor3_1 _21184_ (.A(net1088),
    .B(_10851_),
    .C(_10809_),
    .Y(_03826_));
 sg13g2_nand2_1 _21185_ (.Y(_03827_),
    .A(_03787_),
    .B(_03826_));
 sg13g2_xnor2_1 _21186_ (.Y(_03828_),
    .A(_03825_),
    .B(_03827_));
 sg13g2_a221oi_1 _21187_ (.B2(_03828_),
    .C1(net334),
    .B1(net338),
    .A1(net643),
    .Y(_03829_),
    .A2(net519));
 sg13g2_mux2_1 _21188_ (.A0(_10851_),
    .A1(_11015_),
    .S(net312),
    .X(_03830_));
 sg13g2_a22oi_1 _21189_ (.Y(_03831_),
    .B1(_03830_),
    .B2(net1088),
    .A2(net340),
    .A1(net616));
 sg13g2_or2_1 _21190_ (.X(_03832_),
    .B(_03831_),
    .A(net373));
 sg13g2_xnor2_1 _21191_ (.Y(_03833_),
    .A(_03803_),
    .B(net312));
 sg13g2_nand3_1 _21192_ (.B(_03807_),
    .C(_03833_),
    .A(net373),
    .Y(_03834_));
 sg13g2_a221oi_1 _21193_ (.B2(_03834_),
    .C1(_03794_),
    .B1(_03832_),
    .A1(_03792_),
    .Y(_03835_),
    .A2(_03793_));
 sg13g2_buf_1 _21194_ (.A(_03835_),
    .X(_03836_));
 sg13g2_nand2_1 _21195_ (.Y(_03837_),
    .A(_10884_),
    .B(net322));
 sg13g2_nor2_1 _21196_ (.A(_10884_),
    .B(net322),
    .Y(_03838_));
 sg13g2_a21oi_2 _21197_ (.B1(_03838_),
    .Y(_03839_),
    .A2(_03837_),
    .A1(_10764_));
 sg13g2_nor2_1 _21198_ (.A(_03836_),
    .B(_03839_),
    .Y(_03840_));
 sg13g2_xnor2_1 _21199_ (.Y(_03841_),
    .A(net242),
    .B(_03840_));
 sg13g2_o21ai_1 _21200_ (.B1(_11026_),
    .Y(_03842_),
    .A1(_03737_),
    .A2(_03841_));
 sg13g2_a21o_1 _21201_ (.A2(_03839_),
    .A1(net539),
    .B1(_03836_),
    .X(_03843_));
 sg13g2_mux2_1 _21202_ (.A0(_03840_),
    .A1(_03843_),
    .S(net242),
    .X(_03844_));
 sg13g2_xnor2_1 _21203_ (.Y(_03845_),
    .A(net242),
    .B(_03836_));
 sg13g2_a22oi_1 _21204_ (.Y(_03846_),
    .B1(_03845_),
    .B2(net518),
    .A2(_03844_),
    .A1(_10807_));
 sg13g2_or2_1 _21205_ (.X(_03847_),
    .B(_03846_),
    .A(_03737_));
 sg13g2_a21o_1 _21206_ (.A2(_03847_),
    .A1(_03842_),
    .B1(_11533_),
    .X(_03848_));
 sg13g2_a22oi_1 _21207_ (.Y(_00971_),
    .B1(_03829_),
    .B2(_03848_),
    .A2(net404),
    .A1(_03824_));
 sg13g2_a21oi_1 _21208_ (.A1(net87),
    .A2(_10949_),
    .Y(_03849_),
    .B1(_11031_));
 sg13g2_xnor2_1 _21209_ (.Y(_03850_),
    .A(_03849_),
    .B(net323));
 sg13g2_o21ai_1 _21210_ (.B1(_03850_),
    .Y(_03851_),
    .A1(_11279_),
    .A2(_11308_));
 sg13g2_xnor2_1 _21211_ (.Y(_03852_),
    .A(_10978_),
    .B(_03851_));
 sg13g2_nand2_1 _21212_ (.Y(_03853_),
    .A(net77),
    .B(_03852_));
 sg13g2_nor2_1 _21213_ (.A(_10977_),
    .B(net604),
    .Y(_03854_));
 sg13g2_nor2_1 _21214_ (.A(_10807_),
    .B(_03827_),
    .Y(_03855_));
 sg13g2_mux2_1 _21215_ (.A0(_03854_),
    .A1(_10977_),
    .S(_03855_),
    .X(_03856_));
 sg13g2_a221oi_1 _21216_ (.B2(net1103),
    .C1(net334),
    .B1(_03856_),
    .A1(net953),
    .Y(_03857_),
    .A2(net583));
 sg13g2_nor2_1 _21217_ (.A(_10501_),
    .B(_03766_),
    .Y(_03858_));
 sg13g2_o21ai_1 _21218_ (.B1(_10061_),
    .Y(_03859_),
    .A1(_03821_),
    .A2(_03858_));
 sg13g2_o21ai_1 _21219_ (.B1(_03859_),
    .Y(_03860_),
    .A1(net853),
    .A2(_10061_));
 sg13g2_a21oi_1 _21220_ (.A1(_03853_),
    .A2(_03857_),
    .Y(_00972_),
    .B1(_03860_));
 sg13g2_inv_1 _21221_ (.Y(_03861_),
    .A(\cpu.ex.r_mult[23] ));
 sg13g2_inv_1 _21222_ (.Y(_03862_),
    .A(_10977_));
 sg13g2_and3_1 _21223_ (.X(_03863_),
    .A(_03862_),
    .B(_03825_),
    .C(_03826_));
 sg13g2_nand2_1 _21224_ (.Y(_03864_),
    .A(_03787_),
    .B(_03863_));
 sg13g2_xnor2_1 _21225_ (.Y(_03865_),
    .A(_10501_),
    .B(_03864_));
 sg13g2_a221oi_1 _21226_ (.B2(_03865_),
    .C1(net334),
    .B1(net338),
    .A1(net1037),
    .Y(_03866_),
    .A2(net519));
 sg13g2_nand2_1 _21227_ (.Y(_03867_),
    .A(net242),
    .B(_11026_));
 sg13g2_o21ai_1 _21228_ (.B1(_03867_),
    .Y(_03868_),
    .A1(_03825_),
    .A2(net242));
 sg13g2_a22oi_1 _21229_ (.Y(_03869_),
    .B1(_03868_),
    .B2(_10977_),
    .A2(net243),
    .A1(net616));
 sg13g2_xnor2_1 _21230_ (.Y(_03870_),
    .A(_10807_),
    .B(net243));
 sg13g2_nand3_1 _21231_ (.B(net323),
    .C(_03870_),
    .A(_10978_),
    .Y(_03871_));
 sg13g2_o21ai_1 _21232_ (.B1(_03871_),
    .Y(_03872_),
    .A1(net323),
    .A2(_03869_));
 sg13g2_o21ai_1 _21233_ (.B1(_03825_),
    .Y(_03873_),
    .A1(net243),
    .A2(_03839_));
 sg13g2_nand2_1 _21234_ (.Y(_03874_),
    .A(net243),
    .B(_03839_));
 sg13g2_a22oi_1 _21235_ (.Y(_03875_),
    .B1(_03873_),
    .B2(_03874_),
    .A2(net323),
    .A1(_10977_));
 sg13g2_a21oi_1 _21236_ (.A1(_03862_),
    .A2(net321),
    .Y(_03876_),
    .B1(_03875_));
 sg13g2_nor2_1 _21237_ (.A(net616),
    .B(_03876_),
    .Y(_03877_));
 sg13g2_a21oi_1 _21238_ (.A1(_03836_),
    .A2(_03872_),
    .Y(_03878_),
    .B1(_03877_));
 sg13g2_buf_2 _21239_ (.A(_03878_),
    .X(_03879_));
 sg13g2_xnor2_1 _21240_ (.Y(_03880_),
    .A(_10976_),
    .B(_03879_));
 sg13g2_a21oi_1 _21241_ (.A1(net28),
    .A2(_03880_),
    .Y(_03881_),
    .B1(_11001_));
 sg13g2_and3_1 _21242_ (.X(_03882_),
    .A(_11001_),
    .B(net28),
    .C(_03880_));
 sg13g2_o21ai_1 _21243_ (.B1(_11659_),
    .Y(_03883_),
    .A1(_03881_),
    .A2(_03882_));
 sg13g2_a22oi_1 _21244_ (.Y(_00973_),
    .B1(_03866_),
    .B2(_03883_),
    .A2(net404),
    .A1(_03861_));
 sg13g2_inv_1 _21245_ (.Y(_03884_),
    .A(\cpu.ex.r_mult[24] ));
 sg13g2_nor2_1 _21246_ (.A(net1087),
    .B(_03808_),
    .Y(_03885_));
 sg13g2_xnor2_1 _21247_ (.Y(_03886_),
    .A(_11047_),
    .B(net211));
 sg13g2_o21ai_1 _21248_ (.B1(_03886_),
    .Y(_03887_),
    .A1(_11279_),
    .A2(_11308_));
 sg13g2_xnor2_1 _21249_ (.Y(_03888_),
    .A(_03885_),
    .B(_03887_));
 sg13g2_nand2_1 _21250_ (.Y(_03889_),
    .A(net61),
    .B(_03888_));
 sg13g2_nand2_1 _21251_ (.Y(_03890_),
    .A(_10501_),
    .B(_03863_));
 sg13g2_nor3_1 _21252_ (.A(_03732_),
    .B(_03782_),
    .C(_03890_),
    .Y(_03891_));
 sg13g2_xnor2_1 _21253_ (.Y(_03892_),
    .A(net1087),
    .B(_03891_));
 sg13g2_a221oi_1 _21254_ (.B2(_03892_),
    .C1(net334),
    .B1(net338),
    .A1(net1038),
    .Y(_03893_),
    .A2(net519));
 sg13g2_a22oi_1 _21255_ (.Y(_00974_),
    .B1(_03889_),
    .B2(_03893_),
    .A2(_03759_),
    .A1(_03884_));
 sg13g2_nand2_1 _21256_ (.Y(_03894_),
    .A(_10627_),
    .B(net583));
 sg13g2_nor2_1 _21257_ (.A(_03754_),
    .B(_03821_),
    .Y(_03895_));
 sg13g2_o21ai_1 _21258_ (.B1(_03895_),
    .Y(_03896_),
    .A1(\cpu.ex.r_mult[25] ),
    .A2(_03766_));
 sg13g2_nand2_1 _21259_ (.Y(_03897_),
    .A(_03894_),
    .B(_03896_));
 sg13g2_nor2b_1 _21260_ (.A(net1087),
    .B_N(_03891_),
    .Y(_03898_));
 sg13g2_xnor2_1 _21261_ (.Y(_03899_),
    .A(_11123_),
    .B(_03898_));
 sg13g2_nand2b_1 _21262_ (.Y(_03900_),
    .B(_03894_),
    .A_N(_03769_));
 sg13g2_a21o_1 _21263_ (.A2(_03899_),
    .A1(_03717_),
    .B1(_03900_),
    .X(_03901_));
 sg13g2_and4_1 _21264_ (.A(_11284_),
    .B(_03744_),
    .C(net77),
    .D(_03897_),
    .X(_03902_));
 sg13g2_nor3_1 _21265_ (.A(net184),
    .B(net183),
    .C(_03879_),
    .Y(_03903_));
 sg13g2_nand3b_1 _21266_ (.B(_11513_),
    .C(net518),
    .Y(_03904_),
    .A_N(_03903_));
 sg13g2_o21ai_1 _21267_ (.B1(net183),
    .Y(_03905_),
    .A1(net184),
    .A2(_03879_));
 sg13g2_nand3_1 _21268_ (.B(_03885_),
    .C(_03905_),
    .A(net186),
    .Y(_03906_));
 sg13g2_inv_1 _21269_ (.Y(_03907_),
    .A(_10501_));
 sg13g2_o21ai_1 _21270_ (.B1(_03907_),
    .Y(_03908_),
    .A1(net184),
    .A2(_03879_));
 sg13g2_a22oi_1 _21271_ (.Y(_03909_),
    .B1(_03879_),
    .B2(net184),
    .A2(net183),
    .A1(net1087));
 sg13g2_o21ai_1 _21272_ (.B1(_11513_),
    .Y(_03910_),
    .A1(net1087),
    .A2(net183));
 sg13g2_a21o_1 _21273_ (.A2(_03909_),
    .A1(_03908_),
    .B1(_03910_),
    .X(_03911_));
 sg13g2_a221oi_1 _21274_ (.B2(net184),
    .C1(_11001_),
    .B1(_03879_),
    .A1(_11128_),
    .Y(_03912_),
    .A2(net183));
 sg13g2_o21ai_1 _21275_ (.B1(net186),
    .Y(_03913_),
    .A1(_03903_),
    .A2(_03912_));
 sg13g2_nand4_1 _21276_ (.B(_03906_),
    .C(_03911_),
    .A(_03904_),
    .Y(_03914_),
    .D(_03913_));
 sg13g2_a22oi_1 _21277_ (.Y(_03915_),
    .B1(_03902_),
    .B2(_03914_),
    .A2(_03901_),
    .A1(_03897_));
 sg13g2_nand3_1 _21278_ (.B(_11324_),
    .C(_03897_),
    .A(_11283_),
    .Y(_03916_));
 sg13g2_a21o_1 _21279_ (.A2(_03914_),
    .A1(net28),
    .B1(_03916_),
    .X(_03917_));
 sg13g2_nand2_1 _21280_ (.Y(_00975_),
    .A(_03915_),
    .B(_03917_));
 sg13g2_nand2_1 _21281_ (.Y(_03918_),
    .A(_11133_),
    .B(_03898_));
 sg13g2_nand2_1 _21282_ (.Y(_03919_),
    .A(_10170_),
    .B(_03918_));
 sg13g2_or3_1 _21283_ (.A(_11123_),
    .B(net1087),
    .C(_03890_),
    .X(_03920_));
 sg13g2_nor4_1 _21284_ (.A(_10170_),
    .B(_03732_),
    .C(_03782_),
    .D(_03920_),
    .Y(_03921_));
 sg13g2_buf_2 _21285_ (.A(_03921_),
    .X(_03922_));
 sg13g2_nor2_1 _21286_ (.A(_03719_),
    .B(_03922_),
    .Y(_03923_));
 sg13g2_a221oi_1 _21287_ (.B2(_03923_),
    .C1(_03770_),
    .B1(_03919_),
    .A1(net1089),
    .Y(_03924_),
    .A2(_03755_));
 sg13g2_nor2_1 _21288_ (.A(_11047_),
    .B(_11097_),
    .Y(_03925_));
 sg13g2_a21oi_1 _21289_ (.A1(_11121_),
    .A2(_11136_),
    .Y(_03926_),
    .B1(_03925_));
 sg13g2_xnor2_1 _21290_ (.Y(_03927_),
    .A(_03926_),
    .B(net319));
 sg13g2_o21ai_1 _21291_ (.B1(_03927_),
    .Y(_03928_),
    .A1(_11279_),
    .A2(_11308_));
 sg13g2_nor2_1 _21292_ (.A(_10170_),
    .B(net518),
    .Y(_03929_));
 sg13g2_xnor2_1 _21293_ (.Y(_03930_),
    .A(_03928_),
    .B(_03929_));
 sg13g2_nand2_1 _21294_ (.Y(_03931_),
    .A(net61),
    .B(_03930_));
 sg13g2_a22oi_1 _21295_ (.Y(_00976_),
    .B1(_03924_),
    .B2(_03931_),
    .A2(_03759_),
    .A1(_10073_));
 sg13g2_inv_1 _21296_ (.Y(_03932_),
    .A(\cpu.ex.r_mult[27] ));
 sg13g2_xnor2_1 _21297_ (.Y(_03933_),
    .A(_10073_),
    .B(_03922_));
 sg13g2_a221oi_1 _21298_ (.B2(_03933_),
    .C1(_03770_),
    .B1(net338),
    .A1(net1094),
    .Y(_03934_),
    .A2(net519));
 sg13g2_o21ai_1 _21299_ (.B1(_10170_),
    .Y(_03935_),
    .A1(_11047_),
    .A2(_11097_));
 sg13g2_a21oi_2 _21300_ (.B1(_11136_),
    .Y(_03936_),
    .A2(_03935_),
    .A1(_11120_));
 sg13g2_o21ai_1 _21301_ (.B1(net320),
    .Y(_03937_),
    .A1(_10170_),
    .A2(net616));
 sg13g2_o21ai_1 _21302_ (.B1(_03937_),
    .Y(_03938_),
    .A1(_11121_),
    .A2(_03925_));
 sg13g2_buf_2 _21303_ (.A(_03938_),
    .X(_03939_));
 sg13g2_nor2_1 _21304_ (.A(_03936_),
    .B(_03939_),
    .Y(_03940_));
 sg13g2_xnor2_1 _21305_ (.Y(_03941_),
    .A(net246),
    .B(_03940_));
 sg13g2_nor2_1 _21306_ (.A(_10073_),
    .B(net616),
    .Y(_03942_));
 sg13g2_o21ai_1 _21307_ (.B1(_03942_),
    .Y(_03943_),
    .A1(_03737_),
    .A2(_03941_));
 sg13g2_nand3b_1 _21308_ (.B(_03744_),
    .C(_11140_),
    .Y(_03944_),
    .A_N(_03941_));
 sg13g2_a21o_1 _21309_ (.A2(_03944_),
    .A1(_03943_),
    .B1(_11533_),
    .X(_03945_));
 sg13g2_a22oi_1 _21310_ (.Y(_00977_),
    .B1(_03934_),
    .B2(_03945_),
    .A2(net404),
    .A1(_03932_));
 sg13g2_nand2_1 _21311_ (.Y(_03946_),
    .A(net675),
    .B(net583));
 sg13g2_o21ai_1 _21312_ (.B1(_03895_),
    .Y(_03947_),
    .A1(net1086),
    .A2(_03766_));
 sg13g2_nand2_1 _21313_ (.Y(_03948_),
    .A(_03946_),
    .B(_03947_));
 sg13g2_nor2_1 _21314_ (.A(_10073_),
    .B(_11174_),
    .Y(_03949_));
 sg13g2_nand2_1 _21315_ (.Y(_03950_),
    .A(_03922_),
    .B(_03949_));
 sg13g2_a21o_1 _21316_ (.A2(_03922_),
    .A1(_10072_),
    .B1(_11175_),
    .X(_03951_));
 sg13g2_nand3_1 _21317_ (.B(_03950_),
    .C(_03951_),
    .A(_03717_),
    .Y(_03952_));
 sg13g2_nand3b_1 _21318_ (.B(_03946_),
    .C(_03952_),
    .Y(_03953_),
    .A_N(_03769_));
 sg13g2_nand2_1 _21319_ (.Y(_03954_),
    .A(_03948_),
    .B(_03953_));
 sg13g2_buf_1 _21320_ (.A(_11177_),
    .X(_03955_));
 sg13g2_a21oi_1 _21321_ (.A1(_11137_),
    .A2(_11144_),
    .Y(_03956_),
    .B1(_03808_));
 sg13g2_or2_1 _21322_ (.X(_03957_),
    .B(_03956_),
    .A(_03741_));
 sg13g2_xnor2_1 _21323_ (.Y(_03958_),
    .A(net177),
    .B(_03957_));
 sg13g2_nand3_1 _21324_ (.B(net77),
    .C(_03948_),
    .A(_11178_),
    .Y(_03959_));
 sg13g2_a21o_1 _21325_ (.A2(_03958_),
    .A1(net28),
    .B1(_03959_),
    .X(_03960_));
 sg13g2_a21oi_1 _21326_ (.A1(_03946_),
    .A2(_03947_),
    .Y(_03961_),
    .B1(_11175_));
 sg13g2_nand4_1 _21327_ (.B(net77),
    .C(_03958_),
    .A(net28),
    .Y(_03962_),
    .D(_03961_));
 sg13g2_nand3_1 _21328_ (.B(_03960_),
    .C(_03962_),
    .A(_03954_),
    .Y(_00978_));
 sg13g2_nor4_1 _21329_ (.A(net177),
    .B(net208),
    .C(_03936_),
    .D(_03939_),
    .Y(_03963_));
 sg13g2_nand2_1 _21330_ (.Y(_03964_),
    .A(_11178_),
    .B(net246));
 sg13g2_nor3_1 _21331_ (.A(_03936_),
    .B(_03939_),
    .C(_03964_),
    .Y(_03965_));
 sg13g2_o21ai_1 _21332_ (.B1(_10072_),
    .Y(_03966_),
    .A1(_11175_),
    .A2(net182));
 sg13g2_nor4_1 _21333_ (.A(net518),
    .B(_03936_),
    .C(_03939_),
    .D(_03966_),
    .Y(_03967_));
 sg13g2_nor3_1 _21334_ (.A(net518),
    .B(net208),
    .C(_03966_),
    .Y(_03968_));
 sg13g2_a21o_1 _21335_ (.A2(_11178_),
    .A1(net182),
    .B1(_03968_),
    .X(_03969_));
 sg13g2_nor4_1 _21336_ (.A(_03963_),
    .B(_03965_),
    .C(_03967_),
    .D(_03969_),
    .Y(_03970_));
 sg13g2_xnor2_1 _21337_ (.Y(_03971_),
    .A(net187),
    .B(_03970_));
 sg13g2_a21o_1 _21338_ (.A2(net583),
    .A1(net611),
    .B1(_03769_),
    .X(_03972_));
 sg13g2_inv_1 _21339_ (.Y(_03973_),
    .A(net1086));
 sg13g2_and4_1 _21340_ (.A(_03973_),
    .B(net338),
    .C(_03922_),
    .D(_03949_),
    .X(_03974_));
 sg13g2_nor3_1 _21341_ (.A(_03973_),
    .B(_03719_),
    .C(_03922_),
    .Y(_03975_));
 sg13g2_nor3_1 _21342_ (.A(_03973_),
    .B(_03719_),
    .C(_03949_),
    .Y(_03976_));
 sg13g2_or4_1 _21343_ (.A(_03972_),
    .B(_03974_),
    .C(_03975_),
    .D(_03976_),
    .X(_03977_));
 sg13g2_buf_1 _21344_ (.A(_03977_),
    .X(_03978_));
 sg13g2_nand2_1 _21345_ (.Y(_03979_),
    .A(net1086),
    .B(net539));
 sg13g2_nor2b_1 _21346_ (.A(_03978_),
    .B_N(_03979_),
    .Y(_03980_));
 sg13g2_o21ai_1 _21347_ (.B1(_03980_),
    .Y(_03981_),
    .A1(_03737_),
    .A2(_03971_));
 sg13g2_or4_1 _21348_ (.A(_03737_),
    .B(_03978_),
    .C(_03971_),
    .D(_03979_),
    .X(_03982_));
 sg13g2_nor2_1 _21349_ (.A(_11659_),
    .B(_03978_),
    .Y(_03983_));
 sg13g2_a21oi_1 _21350_ (.A1(_11249_),
    .A2(net404),
    .Y(_03984_),
    .B1(_03983_));
 sg13g2_and3_1 _21351_ (.X(_00979_),
    .A(_03981_),
    .B(_03982_),
    .C(_03984_));
 sg13g2_nor3_1 _21352_ (.A(\cpu.ex.r_mult[30] ),
    .B(net538),
    .C(_10068_),
    .Y(_03985_));
 sg13g2_nor2_1 _21353_ (.A(_10585_),
    .B(_03719_),
    .Y(_03986_));
 sg13g2_nor2_1 _21354_ (.A(_11249_),
    .B(_03719_),
    .Y(_03987_));
 sg13g2_nand3_1 _21355_ (.B(_03922_),
    .C(_03949_),
    .A(net1086),
    .Y(_03988_));
 sg13g2_mux2_1 _21356_ (.A0(_03986_),
    .A1(_03987_),
    .S(_03988_),
    .X(_03989_));
 sg13g2_a21o_1 _21357_ (.A2(net583),
    .A1(net672),
    .B1(_03769_),
    .X(_03990_));
 sg13g2_buf_1 _21358_ (.A(_03990_),
    .X(_03991_));
 sg13g2_nor4_1 _21359_ (.A(_11249_),
    .B(net518),
    .C(_03989_),
    .D(_03991_),
    .Y(_03992_));
 sg13g2_nor2_1 _21360_ (.A(_11249_),
    .B(net518),
    .Y(_03993_));
 sg13g2_nor3_1 _21361_ (.A(_03989_),
    .B(_03991_),
    .C(_03993_),
    .Y(_03994_));
 sg13g2_a21oi_1 _21362_ (.A1(net246),
    .A2(_03942_),
    .Y(_03995_),
    .B1(_11299_));
 sg13g2_o21ai_1 _21363_ (.B1(_03995_),
    .Y(_03996_),
    .A1(_03936_),
    .A2(_03939_));
 sg13g2_a21oi_1 _21364_ (.A1(_10169_),
    .A2(_11140_),
    .Y(_03997_),
    .B1(net177));
 sg13g2_nand3_1 _21365_ (.B(net208),
    .C(_11140_),
    .A(net177),
    .Y(_03998_));
 sg13g2_a21oi_1 _21366_ (.A1(_03973_),
    .A2(net187),
    .Y(_03999_),
    .B1(_11174_));
 sg13g2_nand2_1 _21367_ (.Y(_04000_),
    .A(_03998_),
    .B(_03999_));
 sg13g2_o21ai_1 _21368_ (.B1(_11150_),
    .Y(_04001_),
    .A1(net210),
    .A2(_03997_));
 sg13g2_a21oi_1 _21369_ (.A1(_04000_),
    .A2(_04001_),
    .Y(_04002_),
    .B1(_09213_));
 sg13g2_a21o_1 _21370_ (.A2(_03997_),
    .A1(net210),
    .B1(_04002_),
    .X(_04003_));
 sg13g2_buf_1 _21371_ (.A(_04003_),
    .X(_04004_));
 sg13g2_nand3_1 _21372_ (.B(_03996_),
    .C(_04004_),
    .A(net162),
    .Y(_04005_));
 sg13g2_a21o_1 _21373_ (.A2(_04004_),
    .A1(_03996_),
    .B1(net162),
    .X(_04006_));
 sg13g2_nand3_1 _21374_ (.B(_04005_),
    .C(_04006_),
    .A(net28),
    .Y(_04007_));
 sg13g2_mux2_1 _21375_ (.A0(_03992_),
    .A1(_03994_),
    .S(_04007_),
    .X(_04008_));
 sg13g2_nor3_1 _21376_ (.A(net61),
    .B(_03989_),
    .C(_03991_),
    .Y(_04009_));
 sg13g2_nor3_1 _21377_ (.A(_03985_),
    .B(_04008_),
    .C(_04009_),
    .Y(_00980_));
 sg13g2_inv_1 _21378_ (.Y(_04010_),
    .A(\cpu.ex.r_mult[31] ));
 sg13g2_nor2_1 _21379_ (.A(_11249_),
    .B(_03988_),
    .Y(_04011_));
 sg13g2_xnor2_1 _21380_ (.Y(_04012_),
    .A(_11181_),
    .B(_04011_));
 sg13g2_nand2_1 _21381_ (.Y(_04013_),
    .A(net338),
    .B(_04012_));
 sg13g2_and2_1 _21382_ (.A(_11210_),
    .B(net61),
    .X(_04014_));
 sg13g2_nand2_1 _21383_ (.Y(_04015_),
    .A(net162),
    .B(_03993_));
 sg13g2_nand3_1 _21384_ (.B(_04004_),
    .C(_03993_),
    .A(_03996_),
    .Y(_04016_));
 sg13g2_nand3_1 _21385_ (.B(_04015_),
    .C(_04016_),
    .A(_04005_),
    .Y(_04017_));
 sg13g2_and2_1 _21386_ (.A(net188),
    .B(_04014_),
    .X(_04018_));
 sg13g2_a21o_1 _21387_ (.A2(net583),
    .A1(net890),
    .B1(_03769_),
    .X(_04019_));
 sg13g2_a221oi_1 _21388_ (.B2(_04018_),
    .C1(_04019_),
    .B1(_04017_),
    .A1(_03737_),
    .Y(_04020_),
    .A2(_04014_));
 sg13g2_a22oi_1 _21389_ (.Y(_00981_),
    .B1(_04013_),
    .B2(_04020_),
    .A2(net404),
    .A1(_04010_));
 sg13g2_nand2b_1 _21390_ (.Y(_04021_),
    .B(_08769_),
    .A_N(_11345_));
 sg13g2_mux2_1 _21391_ (.A0(net1111),
    .A1(_04021_),
    .S(_11678_),
    .X(_04022_));
 sg13g2_nor3_1 _21392_ (.A(_11343_),
    .B(_10183_),
    .C(_04022_),
    .Y(_04023_));
 sg13g2_buf_1 _21393_ (.A(_04023_),
    .X(_04024_));
 sg13g2_buf_1 _21394_ (.A(_11354_),
    .X(_04025_));
 sg13g2_nand2_2 _21395_ (.Y(_04026_),
    .A(_08357_),
    .B(_03455_));
 sg13g2_nor3_1 _21396_ (.A(net318),
    .B(_03564_),
    .C(_04026_),
    .Y(_04027_));
 sg13g2_buf_1 _21397_ (.A(_03488_),
    .X(_04028_));
 sg13g2_nor2_1 _21398_ (.A(net209),
    .B(net318),
    .Y(_04029_));
 sg13g2_nor2_1 _21399_ (.A(net317),
    .B(net339),
    .Y(_04030_));
 sg13g2_a21oi_1 _21400_ (.A1(net135),
    .A2(_04029_),
    .Y(_04031_),
    .B1(_04030_));
 sg13g2_nor2_1 _21401_ (.A(net312),
    .B(_04031_),
    .Y(_04032_));
 sg13g2_o21ai_1 _21402_ (.B1(net244),
    .Y(_04033_),
    .A1(_04027_),
    .A2(_04032_));
 sg13g2_nor3_1 _21403_ (.A(net339),
    .B(_11315_),
    .C(_04026_),
    .Y(_04034_));
 sg13g2_nand2_1 _21404_ (.Y(_04035_),
    .A(net201),
    .B(_11668_));
 sg13g2_o21ai_1 _21405_ (.B1(_04035_),
    .Y(_04036_),
    .A1(_00191_),
    .A2(net201));
 sg13g2_buf_1 _21406_ (.A(_04036_),
    .X(_04037_));
 sg13g2_nand2_1 _21407_ (.Y(_04038_),
    .A(net339),
    .B(net245));
 sg13g2_buf_1 _21408_ (.A(_04038_),
    .X(_04039_));
 sg13g2_nor2_1 _21409_ (.A(_11315_),
    .B(_04039_),
    .Y(_04040_));
 sg13g2_buf_1 _21410_ (.A(_04040_),
    .X(_04041_));
 sg13g2_nand2_1 _21411_ (.Y(_04042_),
    .A(net134),
    .B(net133));
 sg13g2_inv_2 _21412_ (.Y(_04043_),
    .A(net247));
 sg13g2_nand2_1 _21413_ (.Y(_04044_),
    .A(_10918_),
    .B(_11331_));
 sg13g2_buf_2 _21414_ (.A(_04044_),
    .X(_04045_));
 sg13g2_nand2_1 _21415_ (.Y(_04046_),
    .A(_11313_),
    .B(net317));
 sg13g2_buf_2 _21416_ (.A(_04046_),
    .X(_04047_));
 sg13g2_nor2_1 _21417_ (.A(_04045_),
    .B(_04047_),
    .Y(_04048_));
 sg13g2_nand2_1 _21418_ (.Y(_04049_),
    .A(_04043_),
    .B(_04048_));
 sg13g2_nand2_1 _21419_ (.Y(_04050_),
    .A(net312),
    .B(_10850_));
 sg13g2_buf_2 _21420_ (.A(_04050_),
    .X(_04051_));
 sg13g2_nor2_1 _21421_ (.A(net185),
    .B(_04051_),
    .Y(_04052_));
 sg13g2_buf_1 _21422_ (.A(_04052_),
    .X(_04053_));
 sg13g2_buf_1 _21423_ (.A(_04053_),
    .X(_04054_));
 sg13g2_nor2_1 _21424_ (.A(_03564_),
    .B(_04039_),
    .Y(_04055_));
 sg13g2_a22oi_1 _21425_ (.Y(_04056_),
    .B1(_04055_),
    .B2(_03455_),
    .A2(net118),
    .A1(_03645_));
 sg13g2_nor2_1 _21426_ (.A(_03564_),
    .B(_04045_),
    .Y(_04057_));
 sg13g2_nor2_1 _21427_ (.A(net185),
    .B(_03564_),
    .Y(_04058_));
 sg13g2_buf_2 _21428_ (.A(_04058_),
    .X(_04059_));
 sg13g2_or2_1 _21429_ (.X(_04060_),
    .B(_04051_),
    .A(_04039_));
 sg13g2_buf_1 _21430_ (.A(_04060_),
    .X(_04061_));
 sg13g2_nand2_1 _21431_ (.Y(_04062_),
    .A(net201),
    .B(_10456_));
 sg13g2_o21ai_1 _21432_ (.B1(_04062_),
    .Y(_04063_),
    .A1(_10399_),
    .A2(net201));
 sg13g2_buf_2 _21433_ (.A(_04063_),
    .X(_04064_));
 sg13g2_nor2_1 _21434_ (.A(net185),
    .B(_04047_),
    .Y(_04065_));
 sg13g2_buf_2 _21435_ (.A(_04065_),
    .X(_04066_));
 sg13g2_nand2_1 _21436_ (.Y(_04067_),
    .A(_04064_),
    .B(_04066_));
 sg13g2_o21ai_1 _21437_ (.B1(_04067_),
    .Y(_04068_),
    .A1(_03483_),
    .A2(_04061_));
 sg13g2_a221oi_1 _21438_ (.B2(net137),
    .C1(_04068_),
    .B1(_04059_),
    .A1(net159),
    .Y(_04069_),
    .A2(_04057_));
 sg13g2_nand4_1 _21439_ (.B(_04049_),
    .C(_04056_),
    .A(_04042_),
    .Y(_04070_),
    .D(_04069_));
 sg13g2_nand2_1 _21440_ (.Y(_04071_),
    .A(net339),
    .B(_11331_));
 sg13g2_buf_1 _21441_ (.A(_04071_),
    .X(_04072_));
 sg13g2_or2_1 _21442_ (.X(_04073_),
    .B(_04051_),
    .A(_04072_));
 sg13g2_buf_1 _21443_ (.A(_04073_),
    .X(_04074_));
 sg13g2_nor2_1 _21444_ (.A(_04045_),
    .B(_04051_),
    .Y(_04075_));
 sg13g2_buf_1 _21445_ (.A(_04075_),
    .X(_04076_));
 sg13g2_nand2_1 _21446_ (.Y(_04077_),
    .A(net140),
    .B(net132));
 sg13g2_o21ai_1 _21447_ (.B1(_04077_),
    .Y(_04078_),
    .A1(_03476_),
    .A2(_04074_));
 sg13g2_nand2_1 _21448_ (.Y(_04079_),
    .A(_11021_),
    .B(_03518_));
 sg13g2_nor2_1 _21449_ (.A(_04039_),
    .B(_04047_),
    .Y(_04080_));
 sg13g2_buf_2 _21450_ (.A(_04080_),
    .X(_04081_));
 sg13g2_buf_1 _21451_ (.A(_04081_),
    .X(_04082_));
 sg13g2_nand2_1 _21452_ (.Y(_04083_),
    .A(net179),
    .B(net117));
 sg13g2_o21ai_1 _21453_ (.B1(_04083_),
    .Y(_04084_),
    .A1(_10492_),
    .A2(_04079_));
 sg13g2_nor4_1 _21454_ (.A(_04034_),
    .B(_04070_),
    .C(_04078_),
    .D(_04084_),
    .Y(_04085_));
 sg13g2_nor2_1 _21455_ (.A(_11315_),
    .B(_04045_),
    .Y(_04086_));
 sg13g2_buf_1 _21456_ (.A(_04086_),
    .X(_04087_));
 sg13g2_buf_1 _21457_ (.A(_04087_),
    .X(_04088_));
 sg13g2_buf_1 _21458_ (.A(net116),
    .X(_04089_));
 sg13g2_buf_1 _21459_ (.A(_04089_),
    .X(_04090_));
 sg13g2_nor2_1 _21460_ (.A(_08357_),
    .B(_09714_),
    .Y(_04091_));
 sg13g2_buf_2 _21461_ (.A(_04091_),
    .X(_04092_));
 sg13g2_a221oi_1 _21462_ (.B2(net180),
    .C1(_04092_),
    .B1(net84),
    .A1(_04033_),
    .Y(_04093_),
    .A2(_04085_));
 sg13g2_nand2_1 _21463_ (.Y(_04094_),
    .A(_11368_),
    .B(_03521_));
 sg13g2_nand2b_1 _21464_ (.Y(_04095_),
    .B(_04094_),
    .A_N(_03623_));
 sg13g2_buf_1 _21465_ (.A(_04095_),
    .X(_04096_));
 sg13g2_o21ai_1 _21466_ (.B1(net244),
    .Y(_04097_),
    .A1(_09716_),
    .A2(_03517_));
 sg13g2_nand2_1 _21467_ (.Y(_04098_),
    .A(_03517_),
    .B(_04096_));
 sg13g2_nand2_1 _21468_ (.Y(_04099_),
    .A(_09716_),
    .B(_04098_));
 sg13g2_inv_1 _21469_ (.Y(_04100_),
    .A(_08842_));
 sg13g2_nand2_1 _21470_ (.Y(_04101_),
    .A(_09716_),
    .B(_03517_));
 sg13g2_o21ai_1 _21471_ (.B1(_04101_),
    .Y(_04102_),
    .A1(_04100_),
    .A2(_03517_));
 sg13g2_nor3_1 _21472_ (.A(net245),
    .B(_04096_),
    .C(_04102_),
    .Y(_04103_));
 sg13g2_a221oi_1 _21473_ (.B2(_04100_),
    .C1(_04103_),
    .B1(_04099_),
    .A1(_04096_),
    .Y(_04104_),
    .A2(_04097_));
 sg13g2_mux2_1 _21474_ (.A0(net1039),
    .A1(net1021),
    .S(_03623_),
    .X(_04105_));
 sg13g2_o21ai_1 _21475_ (.B1(_04094_),
    .Y(_04106_),
    .A1(net1022),
    .A2(_04105_));
 sg13g2_nand2_1 _21476_ (.Y(_04107_),
    .A(_03510_),
    .B(_03515_));
 sg13g2_buf_2 _21477_ (.A(_04107_),
    .X(_04108_));
 sg13g2_buf_1 _21478_ (.A(_04108_),
    .X(_04109_));
 sg13g2_nand3_1 _21479_ (.B(net176),
    .C(net84),
    .A(net1100),
    .Y(_04110_));
 sg13g2_a21oi_1 _21480_ (.A1(net1040),
    .A2(net186),
    .Y(_04111_),
    .B1(net234));
 sg13g2_nor4_1 _21481_ (.A(net1109),
    .B(_09735_),
    .C(\cpu.dec.r_op[8] ),
    .D(_09748_),
    .Y(_04112_));
 sg13g2_nor4_1 _21482_ (.A(_08842_),
    .B(net1108),
    .C(_09716_),
    .D(_09767_),
    .Y(_04113_));
 sg13g2_and3_1 _21483_ (.X(_04114_),
    .A(_04092_),
    .B(_04112_),
    .C(_04113_));
 sg13g2_buf_1 _21484_ (.A(_04114_),
    .X(_04115_));
 sg13g2_buf_1 _21485_ (.A(_04115_),
    .X(_04116_));
 sg13g2_nand2_1 _21486_ (.Y(_04117_),
    .A(net244),
    .B(_04108_));
 sg13g2_xor2_1 _21487_ (.B(_04096_),
    .A(_04117_),
    .X(_04118_));
 sg13g2_o21ai_1 _21488_ (.B1(_04118_),
    .Y(_04119_),
    .A1(_09767_),
    .A2(net582));
 sg13g2_nand4_1 _21489_ (.B(_04110_),
    .C(_04111_),
    .A(_04106_),
    .Y(_04120_),
    .D(_04119_));
 sg13g2_nor3_1 _21490_ (.A(_04093_),
    .B(_04104_),
    .C(_04120_),
    .Y(_04121_));
 sg13g2_a21oi_1 _21491_ (.A1(net234),
    .A2(_11378_),
    .Y(_04122_),
    .B1(_04121_));
 sg13g2_nand2_1 _21492_ (.Y(_04123_),
    .A(net85),
    .B(_04122_));
 sg13g2_and2_1 _21493_ (.A(net379),
    .B(_10181_),
    .X(_04124_));
 sg13g2_buf_2 _21494_ (.A(_04124_),
    .X(_04125_));
 sg13g2_and4_1 _21495_ (.A(_08769_),
    .B(net737),
    .C(_04125_),
    .D(_11679_),
    .X(_04126_));
 sg13g2_buf_1 _21496_ (.A(_04126_),
    .X(_04127_));
 sg13g2_and2_1 _21497_ (.A(_09018_),
    .B(net379),
    .X(_04128_));
 sg13g2_buf_1 _21498_ (.A(_04128_),
    .X(_04129_));
 sg13g2_nand2_1 _21499_ (.Y(_04130_),
    .A(_11342_),
    .B(_04129_));
 sg13g2_nand2_1 _21500_ (.Y(_04131_),
    .A(_09028_),
    .B(_09200_));
 sg13g2_a21oi_1 _21501_ (.A1(_04130_),
    .A2(_04131_),
    .Y(_04132_),
    .B1(net1111));
 sg13g2_nand4_1 _21502_ (.B(_09029_),
    .C(_09075_),
    .A(net1110),
    .Y(_04133_),
    .D(net737));
 sg13g2_nand2_1 _21503_ (.Y(_04134_),
    .A(_09127_),
    .B(_04133_));
 sg13g2_nor4_1 _21504_ (.A(_04023_),
    .B(net83),
    .C(_04132_),
    .D(_04134_),
    .Y(_04135_));
 sg13g2_buf_1 _21505_ (.A(_04135_),
    .X(_04136_));
 sg13g2_buf_1 _21506_ (.A(_04136_),
    .X(_04137_));
 sg13g2_a22oi_1 _21507_ (.Y(_04138_),
    .B1(_04137_),
    .B2(net919),
    .A2(net83),
    .A1(_10206_));
 sg13g2_nand2_1 _21508_ (.Y(_00982_),
    .A(_04123_),
    .B(_04138_));
 sg13g2_or2_1 _21509_ (.X(_04139_),
    .B(_03661_),
    .A(_03655_));
 sg13g2_buf_1 _21510_ (.A(_04139_),
    .X(_04140_));
 sg13g2_xor2_1 _21511_ (.B(_04140_),
    .A(_03584_),
    .X(_04141_));
 sg13g2_inv_1 _21512_ (.Y(_04142_),
    .A(_03639_));
 sg13g2_and2_1 _21513_ (.A(_03637_),
    .B(_04142_),
    .X(_04143_));
 sg13g2_buf_1 _21514_ (.A(_04143_),
    .X(_04144_));
 sg13g2_or2_1 _21515_ (.X(_04145_),
    .B(_03634_),
    .A(_03633_));
 sg13g2_nand2_1 _21516_ (.Y(_04146_),
    .A(_03618_),
    .B(_03632_));
 sg13g2_a22oi_1 _21517_ (.Y(_04147_),
    .B1(_03640_),
    .B2(_04146_),
    .A2(_04145_),
    .A1(_03635_));
 sg13g2_xnor2_1 _21518_ (.Y(_04148_),
    .A(_04144_),
    .B(_04147_));
 sg13g2_a21oi_1 _21519_ (.A1(_09716_),
    .A2(_04148_),
    .Y(_04149_),
    .B1(net582));
 sg13g2_buf_1 _21520_ (.A(_03654_),
    .X(_04150_));
 sg13g2_nand3_1 _21521_ (.B(_11331_),
    .C(_11021_),
    .A(net318),
    .Y(_04151_));
 sg13g2_buf_1 _21522_ (.A(_04151_),
    .X(_04152_));
 sg13g2_inv_1 _21523_ (.Y(_04153_),
    .A(_09714_));
 sg13g2_buf_1 _21524_ (.A(_04066_),
    .X(_04154_));
 sg13g2_nor2_1 _21525_ (.A(_10918_),
    .B(_11331_),
    .Y(_04155_));
 sg13g2_nand2_1 _21526_ (.Y(_04156_),
    .A(net339),
    .B(_03590_));
 sg13g2_a22oi_1 _21527_ (.Y(_04157_),
    .B1(_04156_),
    .B2(net244),
    .A2(_04155_),
    .A1(net137));
 sg13g2_nor2_1 _21528_ (.A(_11315_),
    .B(_04157_),
    .Y(_04158_));
 sg13g2_a21oi_1 _21529_ (.A1(net142),
    .A2(net114),
    .Y(_04159_),
    .B1(_04158_));
 sg13g2_a21oi_1 _21530_ (.A1(_11021_),
    .A2(_11318_),
    .Y(_04160_),
    .B1(net157));
 sg13g2_o21ai_1 _21531_ (.B1(net1055),
    .Y(_04161_),
    .A1(_04158_),
    .A2(_04160_));
 sg13g2_o21ai_1 _21532_ (.B1(_04161_),
    .Y(_04162_),
    .A1(_04153_),
    .A2(_04159_));
 sg13g2_o21ai_1 _21533_ (.B1(_04162_),
    .Y(_04163_),
    .A1(net115),
    .A2(net175));
 sg13g2_nor2_1 _21534_ (.A(_11315_),
    .B(_04072_),
    .Y(_04164_));
 sg13g2_buf_1 _21535_ (.A(_04164_),
    .X(_04165_));
 sg13g2_a21oi_1 _21536_ (.A1(net135),
    .A2(net131),
    .Y(_04166_),
    .B1(net116));
 sg13g2_nor2_2 _21537_ (.A(_04072_),
    .B(_04051_),
    .Y(_04167_));
 sg13g2_nand2_1 _21538_ (.Y(_04168_),
    .A(net176),
    .B(_04167_));
 sg13g2_or2_1 _21539_ (.X(_04169_),
    .B(_04051_),
    .A(_04045_));
 sg13g2_nand2_1 _21540_ (.Y(_04170_),
    .A(_03453_),
    .B(_10325_));
 sg13g2_o21ai_1 _21541_ (.B1(_04170_),
    .Y(_04171_),
    .A1(_10206_),
    .A2(_03453_));
 sg13g2_buf_1 _21542_ (.A(_04171_),
    .X(_04172_));
 sg13g2_nor2_1 _21543_ (.A(_04039_),
    .B(_04051_),
    .Y(_04173_));
 sg13g2_buf_1 _21544_ (.A(_04173_),
    .X(_04174_));
 sg13g2_a22oi_1 _21545_ (.Y(_04175_),
    .B1(_04081_),
    .B2(_04064_),
    .A2(net130),
    .A1(_04172_));
 sg13g2_o21ai_1 _21546_ (.B1(_04175_),
    .Y(_04176_),
    .A1(net180),
    .A2(_04169_));
 sg13g2_or2_1 _21547_ (.X(_04177_),
    .B(_04047_),
    .A(net185));
 sg13g2_buf_1 _21548_ (.A(_04177_),
    .X(_04178_));
 sg13g2_nor2_1 _21549_ (.A(_03534_),
    .B(_04178_),
    .Y(_04179_));
 sg13g2_nand2_2 _21550_ (.Y(_04180_),
    .A(_11021_),
    .B(_04155_));
 sg13g2_nor2_1 _21551_ (.A(net198),
    .B(_04180_),
    .Y(_04181_));
 sg13g2_buf_1 _21552_ (.A(net200),
    .X(_04182_));
 sg13g2_or2_1 _21553_ (.X(_04183_),
    .B(_04051_),
    .A(net185));
 sg13g2_buf_1 _21554_ (.A(_04183_),
    .X(_04184_));
 sg13g2_nor2_1 _21555_ (.A(_04072_),
    .B(_04047_),
    .Y(_04185_));
 sg13g2_buf_1 _21556_ (.A(_04185_),
    .X(_04186_));
 sg13g2_nand2_1 _21557_ (.Y(_04187_),
    .A(_03505_),
    .B(_04186_));
 sg13g2_o21ai_1 _21558_ (.B1(_04187_),
    .Y(_04188_),
    .A1(_04182_),
    .A2(_04184_));
 sg13g2_nor4_1 _21559_ (.A(_04176_),
    .B(_04179_),
    .C(_04181_),
    .D(_04188_),
    .Y(_04189_));
 sg13g2_nand4_1 _21560_ (.B(_04166_),
    .C(_04168_),
    .A(_04049_),
    .Y(_04190_),
    .D(_04189_));
 sg13g2_nand2_1 _21561_ (.Y(_04191_),
    .A(_03663_),
    .B(net97));
 sg13g2_nand3_1 _21562_ (.B(_04190_),
    .C(_04191_),
    .A(net1100),
    .Y(_04192_));
 sg13g2_inv_1 _21563_ (.Y(_04193_),
    .A(_09735_));
 sg13g2_nand2_1 _21564_ (.Y(_04194_),
    .A(_10169_),
    .B(net119));
 sg13g2_or2_1 _21565_ (.X(_04195_),
    .B(_03655_),
    .A(net1108));
 sg13g2_o21ai_1 _21566_ (.B1(_04195_),
    .Y(_04196_),
    .A1(net1099),
    .A2(_04194_));
 sg13g2_a21oi_1 _21567_ (.A1(_04193_),
    .A2(_04196_),
    .Y(_04197_),
    .B1(_03661_));
 sg13g2_a21oi_1 _21568_ (.A1(net1040),
    .A2(net312),
    .Y(_04198_),
    .B1(_04197_));
 sg13g2_nand4_1 _21569_ (.B(_04163_),
    .C(_04192_),
    .A(_04149_),
    .Y(_04199_),
    .D(_04198_));
 sg13g2_a21oi_1 _21570_ (.A1(net901),
    .A2(_04141_),
    .Y(_04200_),
    .B1(_04199_));
 sg13g2_nand3_1 _21571_ (.B(_04112_),
    .C(_04113_),
    .A(_04092_),
    .Y(_04201_));
 sg13g2_buf_1 _21572_ (.A(_04201_),
    .X(_04202_));
 sg13g2_nand2_1 _21573_ (.Y(_04203_),
    .A(net319),
    .B(_03663_));
 sg13g2_nand2_1 _21574_ (.Y(_04204_),
    .A(net320),
    .B(_03578_));
 sg13g2_o21ai_1 _21575_ (.B1(_04204_),
    .Y(_04205_),
    .A1(_03650_),
    .A2(_03653_));
 sg13g2_nand2_2 _21576_ (.Y(_04206_),
    .A(_04203_),
    .B(_04205_));
 sg13g2_xor2_1 _21577_ (.B(_04140_),
    .A(_04206_),
    .X(_04207_));
 sg13g2_nor2_1 _21578_ (.A(_04202_),
    .B(_04207_),
    .Y(_04208_));
 sg13g2_nor3_1 _21579_ (.A(net234),
    .B(_04200_),
    .C(_04208_),
    .Y(_04209_));
 sg13g2_a21o_1 _21580_ (.A2(\cpu.ex.c_mult[11] ),
    .A1(net234),
    .B1(_04209_),
    .X(_04210_));
 sg13g2_nand2_1 _21581_ (.Y(_04211_),
    .A(net85),
    .B(_04210_));
 sg13g2_buf_1 _21582_ (.A(_11074_),
    .X(_04212_));
 sg13g2_nand2_2 _21583_ (.Y(_04213_),
    .A(_08147_),
    .B(net1117));
 sg13g2_nor2_1 _21584_ (.A(net918),
    .B(_04213_),
    .Y(_04214_));
 sg13g2_and2_1 _21585_ (.A(net1116),
    .B(_04214_),
    .X(_04215_));
 sg13g2_buf_1 _21586_ (.A(_04215_),
    .X(_04216_));
 sg13g2_nand3_1 _21587_ (.B(_08669_),
    .C(_04216_),
    .A(_08701_),
    .Y(_04217_));
 sg13g2_or2_1 _21588_ (.X(_04218_),
    .B(_04217_),
    .A(_08680_));
 sg13g2_buf_1 _21589_ (.A(_04218_),
    .X(_04219_));
 sg13g2_nor2_1 _21590_ (.A(net948),
    .B(_04219_),
    .Y(_04220_));
 sg13g2_nand3_1 _21591_ (.B(_08710_),
    .C(_04220_),
    .A(_08719_),
    .Y(_04221_));
 sg13g2_xor2_1 _21592_ (.B(_04221_),
    .A(_10676_),
    .X(_04222_));
 sg13g2_buf_1 _21593_ (.A(net83),
    .X(_04223_));
 sg13g2_a22oi_1 _21594_ (.Y(_04224_),
    .B1(_04222_),
    .B2(net76),
    .A2(net33),
    .A1(\cpu.ex.pc[11] ));
 sg13g2_nand2_1 _21595_ (.Y(_00983_),
    .A(_04211_),
    .B(_04224_));
 sg13g2_nor2_1 _21596_ (.A(_08659_),
    .B(_04221_),
    .Y(_04225_));
 sg13g2_xnor2_1 _21597_ (.Y(_04226_),
    .A(_00289_),
    .B(_04225_));
 sg13g2_a22oi_1 _21598_ (.Y(_04227_),
    .B1(_04226_),
    .B2(_04223_),
    .A2(net33),
    .A1(net688));
 sg13g2_or3_1 _21599_ (.A(_03477_),
    .B(_03585_),
    .C(_03586_),
    .X(_04228_));
 sg13g2_o21ai_1 _21600_ (.B1(_03477_),
    .Y(_04229_),
    .A1(_03585_),
    .A2(_03586_));
 sg13g2_nand3_1 _21601_ (.B(_04228_),
    .C(_04229_),
    .A(net901),
    .Y(_04230_));
 sg13g2_a21oi_2 _21602_ (.B1(_03661_),
    .Y(_04231_),
    .A2(_04194_),
    .A1(_04206_));
 sg13g2_xor2_1 _21603_ (.B(_03477_),
    .A(_04231_),
    .X(_04232_));
 sg13g2_a21oi_2 _21604_ (.B1(_11354_),
    .Y(_04233_),
    .A2(_04148_),
    .A1(_09716_));
 sg13g2_o21ai_1 _21605_ (.B1(net244),
    .Y(_04234_),
    .A1(net318),
    .A2(_03455_));
 sg13g2_nand2_1 _21606_ (.Y(_04235_),
    .A(net159),
    .B(_04155_));
 sg13g2_a21oi_1 _21607_ (.A1(_04234_),
    .A2(_04235_),
    .Y(_04236_),
    .B1(_11315_));
 sg13g2_nand2b_1 _21608_ (.Y(_04237_),
    .B(_04088_),
    .A_N(net137));
 sg13g2_nand3_1 _21609_ (.B(_04236_),
    .C(_04237_),
    .A(_09714_),
    .Y(_04238_));
 sg13g2_nand2_1 _21610_ (.Y(_04239_),
    .A(_11177_),
    .B(_03654_));
 sg13g2_mux2_1 _21611_ (.A0(net1099),
    .A1(net1108),
    .S(_04239_),
    .X(_04240_));
 sg13g2_nand2_1 _21612_ (.Y(_04241_),
    .A(net182),
    .B(_03476_));
 sg13g2_o21ai_1 _21613_ (.B1(_04241_),
    .Y(_04242_),
    .A1(_09735_),
    .A2(_04240_));
 sg13g2_nand2_1 _21614_ (.Y(_04243_),
    .A(_04238_),
    .B(_04242_));
 sg13g2_a21oi_1 _21615_ (.A1(net1040),
    .A2(net373),
    .Y(_04244_),
    .B1(_04243_));
 sg13g2_and2_1 _21616_ (.A(net1055),
    .B(_04237_),
    .X(_04245_));
 sg13g2_o21ai_1 _21617_ (.B1(_04245_),
    .Y(_04246_),
    .A1(_04160_),
    .A2(_04236_));
 sg13g2_nand2_1 _21618_ (.Y(_04247_),
    .A(net140),
    .B(net133));
 sg13g2_nand2_1 _21619_ (.Y(_04248_),
    .A(_04043_),
    .B(_04081_));
 sg13g2_buf_1 _21620_ (.A(_03568_),
    .X(_04249_));
 sg13g2_a22oi_1 _21621_ (.Y(_04250_),
    .B1(net130),
    .B2(_04249_),
    .A2(_04059_),
    .A1(net176));
 sg13g2_nand3_1 _21622_ (.B(_04248_),
    .C(_04250_),
    .A(_04247_),
    .Y(_04251_));
 sg13g2_buf_1 _21623_ (.A(_04048_),
    .X(_04252_));
 sg13g2_buf_1 _21624_ (.A(_04186_),
    .X(_04253_));
 sg13g2_a22oi_1 _21625_ (.Y(_04254_),
    .B1(net129),
    .B2(_04064_),
    .A2(net155),
    .A1(net179));
 sg13g2_a22oi_1 _21626_ (.Y(_04255_),
    .B1(net132),
    .B2(net134),
    .A2(net114),
    .A1(net135));
 sg13g2_a21oi_1 _21627_ (.A1(_03645_),
    .A2(_04165_),
    .Y(_04256_),
    .B1(net116));
 sg13g2_buf_1 _21628_ (.A(_04172_),
    .X(_04257_));
 sg13g2_a22oi_1 _21629_ (.Y(_04258_),
    .B1(_04167_),
    .B2(net113),
    .A2(net118),
    .A1(net199));
 sg13g2_nand4_1 _21630_ (.B(_04255_),
    .C(_04256_),
    .A(_04254_),
    .Y(_04259_),
    .D(_04258_));
 sg13g2_inv_2 _21631_ (.Y(_04260_),
    .A(net1100));
 sg13g2_a21oi_1 _21632_ (.A1(net138),
    .A2(_04090_),
    .Y(_04261_),
    .B1(_04260_));
 sg13g2_o21ai_1 _21633_ (.B1(_04261_),
    .Y(_04262_),
    .A1(_04251_),
    .A2(_04259_));
 sg13g2_nand4_1 _21634_ (.B(_04244_),
    .C(_04246_),
    .A(_04233_),
    .Y(_04263_),
    .D(_04262_));
 sg13g2_a21oi_1 _21635_ (.A1(_04116_),
    .A2(_04232_),
    .Y(_04264_),
    .B1(_04263_));
 sg13g2_or2_1 _21636_ (.X(_04265_),
    .B(_11352_),
    .A(_10067_));
 sg13g2_buf_1 _21637_ (.A(_04265_),
    .X(_04266_));
 sg13g2_nor4_1 _21638_ (.A(_04266_),
    .B(_11571_),
    .C(_11592_),
    .D(_11594_),
    .Y(_04267_));
 sg13g2_a21oi_1 _21639_ (.A1(_04230_),
    .A2(_04264_),
    .Y(_04268_),
    .B1(_04267_));
 sg13g2_nand2_1 _21640_ (.Y(_04269_),
    .A(_04024_),
    .B(_04268_));
 sg13g2_nand2_1 _21641_ (.Y(_00984_),
    .A(_04227_),
    .B(_04269_));
 sg13g2_nor3_1 _21642_ (.A(net120),
    .B(_03577_),
    .C(_03582_),
    .Y(_04270_));
 sg13g2_nand2_1 _21643_ (.Y(_04271_),
    .A(_03592_),
    .B(_04270_));
 sg13g2_o21ai_1 _21644_ (.B1(_04271_),
    .Y(_04272_),
    .A1(net177),
    .A2(net138));
 sg13g2_nand2_1 _21645_ (.Y(_04273_),
    .A(_03592_),
    .B(_03474_));
 sg13g2_nand2_1 _21646_ (.Y(_04274_),
    .A(_03485_),
    .B(_04270_));
 sg13g2_nand3_1 _21647_ (.B(_04273_),
    .C(_04274_),
    .A(net208),
    .Y(_04275_));
 sg13g2_o21ai_1 _21648_ (.B1(_04275_),
    .Y(_04276_),
    .A1(_11564_),
    .A2(_04272_));
 sg13g2_o21ai_1 _21649_ (.B1(net177),
    .Y(_04277_),
    .A1(net208),
    .A2(net138));
 sg13g2_nand2_1 _21650_ (.Y(_04278_),
    .A(net177),
    .B(net158));
 sg13g2_nand2_1 _21651_ (.Y(_04279_),
    .A(_03584_),
    .B(_04278_));
 sg13g2_a221oi_1 _21652_ (.B2(net120),
    .C1(_04100_),
    .B1(_04279_),
    .A1(_04150_),
    .Y(_04280_),
    .A2(_04277_));
 sg13g2_nand2_1 _21653_ (.Y(_04281_),
    .A(_04231_),
    .B(_04241_));
 sg13g2_nand3b_1 _21654_ (.B(net120),
    .C(_04239_),
    .Y(_04282_),
    .A_N(_04231_));
 sg13g2_o21ai_1 _21655_ (.B1(_04282_),
    .Y(_04283_),
    .A1(net120),
    .A2(_04281_));
 sg13g2_or2_1 _21656_ (.X(_04284_),
    .B(_03676_),
    .A(_03610_));
 sg13g2_or2_1 _21657_ (.X(_04285_),
    .B(_04239_),
    .A(net120));
 sg13g2_o21ai_1 _21658_ (.B1(_04285_),
    .Y(_04286_),
    .A1(_04284_),
    .A2(_04241_));
 sg13g2_nor2_1 _21659_ (.A(net177),
    .B(net158),
    .Y(_04287_));
 sg13g2_a21oi_1 _21660_ (.A1(_03595_),
    .A2(_04278_),
    .Y(_04288_),
    .B1(_04287_));
 sg13g2_or2_1 _21661_ (.X(_04289_),
    .B(_04278_),
    .A(net120));
 sg13g2_o21ai_1 _21662_ (.B1(_04289_),
    .Y(_04290_),
    .A1(_04284_),
    .A2(_04288_));
 sg13g2_a22oi_1 _21663_ (.Y(_04291_),
    .B1(_04290_),
    .B2(_08844_),
    .A2(_04286_),
    .A1(net582));
 sg13g2_a22oi_1 _21664_ (.Y(_04292_),
    .B1(net97),
    .B2(net141),
    .A2(_04041_),
    .A1(net142));
 sg13g2_o21ai_1 _21665_ (.B1(net1055),
    .Y(_04293_),
    .A1(net142),
    .A2(_04088_));
 sg13g2_a21oi_1 _21666_ (.A1(net139),
    .A2(net116),
    .Y(_04294_),
    .B1(_04293_));
 sg13g2_a21oi_1 _21667_ (.A1(net1109),
    .A2(net242),
    .Y(_04295_),
    .B1(_04294_));
 sg13g2_o21ai_1 _21668_ (.B1(_04295_),
    .Y(_04296_),
    .A1(_04153_),
    .A2(_04292_));
 sg13g2_mux2_1 _21669_ (.A0(_08996_),
    .A1(_09749_),
    .S(_03676_),
    .X(_04297_));
 sg13g2_o21ai_1 _21670_ (.B1(_03609_),
    .Y(_04298_),
    .A1(_09736_),
    .A2(_04297_));
 sg13g2_nand2b_1 _21671_ (.Y(_04299_),
    .B(_04298_),
    .A_N(_04296_));
 sg13g2_nand2_1 _21672_ (.Y(_04300_),
    .A(net119),
    .B(net133));
 sg13g2_nor2_1 _21673_ (.A(_03663_),
    .B(_04079_),
    .Y(_04301_));
 sg13g2_a21oi_1 _21674_ (.A1(net113),
    .A2(_04059_),
    .Y(_04302_),
    .B1(_04301_));
 sg13g2_a22oi_1 _21675_ (.Y(_04303_),
    .B1(net132),
    .B2(net199),
    .A2(net130),
    .A1(net134));
 sg13g2_a22oi_1 _21676_ (.Y(_04304_),
    .B1(net114),
    .B2(_03645_),
    .A2(_04057_),
    .A1(net176));
 sg13g2_and4_1 _21677_ (.A(_04300_),
    .B(_04302_),
    .C(_04303_),
    .D(_04304_),
    .X(_04305_));
 sg13g2_or2_1 _21678_ (.X(_04306_),
    .B(_04047_),
    .A(_04045_));
 sg13g2_buf_1 _21679_ (.A(_04306_),
    .X(_04307_));
 sg13g2_nor2_1 _21680_ (.A(_10717_),
    .B(_04307_),
    .Y(_04308_));
 sg13g2_nor2_1 _21681_ (.A(net178),
    .B(_04184_),
    .Y(_04309_));
 sg13g2_or2_1 _21682_ (.X(_04310_),
    .B(_04047_),
    .A(_04072_));
 sg13g2_o21ai_1 _21683_ (.B1(_04083_),
    .Y(_04311_),
    .A1(net247),
    .A2(_04310_));
 sg13g2_o21ai_1 _21684_ (.B1(net175),
    .Y(_04312_),
    .A1(_03498_),
    .A2(_04074_));
 sg13g2_nor4_1 _21685_ (.A(_04308_),
    .B(_04309_),
    .C(_04311_),
    .D(_04312_),
    .Y(_04313_));
 sg13g2_a221oi_1 _21686_ (.B2(_04313_),
    .C1(_04260_),
    .B1(_04305_),
    .A1(net158),
    .Y(_04314_),
    .A2(_04090_));
 sg13g2_nor2_1 _21687_ (.A(_04299_),
    .B(_04314_),
    .Y(_04315_));
 sg13g2_nand3_1 _21688_ (.B(_04291_),
    .C(_04315_),
    .A(_04233_),
    .Y(_04316_));
 sg13g2_a221oi_1 _21689_ (.B2(net582),
    .C1(_04316_),
    .B1(_04283_),
    .A1(_04276_),
    .Y(_04317_),
    .A2(_04280_));
 sg13g2_buf_1 _21690_ (.A(_04266_),
    .X(_04318_));
 sg13g2_nor2_1 _21691_ (.A(net233),
    .B(\cpu.ex.c_mult[13] ),
    .Y(_04319_));
 sg13g2_nor2_1 _21692_ (.A(_04317_),
    .B(_04319_),
    .Y(_04320_));
 sg13g2_nand2_1 _21693_ (.Y(_04321_),
    .A(net688),
    .B(_04225_));
 sg13g2_xor2_1 _21694_ (.B(_04321_),
    .A(_00196_),
    .X(_04322_));
 sg13g2_a22oi_1 _21695_ (.Y(_04323_),
    .B1(_04322_),
    .B2(net83),
    .A2(_04136_),
    .A1(net788));
 sg13g2_inv_1 _21696_ (.Y(_04324_),
    .A(_04323_));
 sg13g2_a21o_1 _21697_ (.A2(_04320_),
    .A1(net85),
    .B1(_04324_),
    .X(_00985_));
 sg13g2_inv_1 _21698_ (.Y(_04325_),
    .A(_04023_));
 sg13g2_nor2_2 _21699_ (.A(_03606_),
    .B(_03607_),
    .Y(_04326_));
 sg13g2_mux2_1 _21700_ (.A0(_03597_),
    .A1(_03587_),
    .S(_04326_),
    .X(_04327_));
 sg13g2_buf_1 _21701_ (.A(net137),
    .X(_04328_));
 sg13g2_nand3b_1 _21702_ (.B(net158),
    .C(net187),
    .Y(_04329_),
    .A_N(net112));
 sg13g2_nand2_1 _21703_ (.Y(_04330_),
    .A(net210),
    .B(net112));
 sg13g2_a221oi_1 _21704_ (.B2(_04330_),
    .C1(_03661_),
    .B1(_04329_),
    .A1(_04206_),
    .Y(_04331_),
    .A2(_04194_));
 sg13g2_and2_1 _21705_ (.A(net112),
    .B(net115),
    .X(_04332_));
 sg13g2_o21ai_1 _21706_ (.B1(_03955_),
    .Y(_04333_),
    .A1(_04331_),
    .A2(_04332_));
 sg13g2_o21ai_1 _21707_ (.B1(_04326_),
    .Y(_04334_),
    .A1(_03610_),
    .A2(_03677_));
 sg13g2_o21ai_1 _21708_ (.B1(_04334_),
    .Y(_04335_),
    .A1(_04326_),
    .A2(_04333_));
 sg13g2_a21o_1 _21709_ (.A2(_03472_),
    .A1(_08843_),
    .B1(net1039),
    .X(_04336_));
 sg13g2_a21oi_1 _21710_ (.A1(net179),
    .A2(net129),
    .Y(_04337_),
    .B1(net116));
 sg13g2_a22oi_1 _21711_ (.Y(_04338_),
    .B1(net132),
    .B2(_04064_),
    .A2(_04059_),
    .A1(net156));
 sg13g2_nand2_1 _21712_ (.Y(_04339_),
    .A(net140),
    .B(_04066_));
 sg13g2_o21ai_1 _21713_ (.B1(_04339_),
    .Y(_04340_),
    .A1(_10492_),
    .A2(_04061_));
 sg13g2_a221oi_1 _21714_ (.B2(net119),
    .C1(_04340_),
    .B1(net131),
    .A1(net115),
    .Y(_04341_),
    .A2(net133));
 sg13g2_nor2_1 _21715_ (.A(_03521_),
    .B(_04045_),
    .Y(_04342_));
 sg13g2_nor2_1 _21716_ (.A(_03517_),
    .B(_04039_),
    .Y(_04343_));
 sg13g2_o21ai_1 _21717_ (.B1(_03500_),
    .Y(_04344_),
    .A1(_04342_),
    .A2(_04343_));
 sg13g2_nor2_1 _21718_ (.A(net198),
    .B(_04307_),
    .Y(_04345_));
 sg13g2_a21oi_1 _21719_ (.A1(net135),
    .A2(_04081_),
    .Y(_04346_),
    .B1(_04345_));
 sg13g2_a22oi_1 _21720_ (.Y(_04347_),
    .B1(_04167_),
    .B2(net134),
    .A2(net118),
    .A1(_04043_));
 sg13g2_and3_1 _21721_ (.X(_04348_),
    .A(_04344_),
    .B(_04346_),
    .C(_04347_));
 sg13g2_nand4_1 _21722_ (.B(_04338_),
    .C(_04341_),
    .A(_04337_),
    .Y(_04349_),
    .D(_04348_));
 sg13g2_nand3_1 _21723_ (.B(_04237_),
    .C(_04349_),
    .A(net1100),
    .Y(_04350_));
 sg13g2_nor2_1 _21724_ (.A(_04153_),
    .B(net157),
    .Y(_04351_));
 sg13g2_a22oi_1 _21725_ (.Y(_04352_),
    .B1(net84),
    .B2(_04351_),
    .A2(_03606_),
    .A1(_09749_));
 sg13g2_nand2_1 _21726_ (.Y(_04353_),
    .A(net162),
    .B(net139));
 sg13g2_a22oi_1 _21727_ (.Y(_04354_),
    .B1(_04353_),
    .B2(net1022),
    .A2(_11000_),
    .A1(_08892_));
 sg13g2_nor2_1 _21728_ (.A(_04202_),
    .B(_04326_),
    .Y(_04355_));
 sg13g2_nand2b_1 _21729_ (.Y(_04356_),
    .B(_04239_),
    .A_N(_04328_));
 sg13g2_nand3_1 _21730_ (.B(_04355_),
    .C(_04356_),
    .A(_11271_),
    .Y(_04357_));
 sg13g2_nand4_1 _21731_ (.B(_04352_),
    .C(_04354_),
    .A(_04350_),
    .Y(_04358_),
    .D(_04357_));
 sg13g2_a21oi_1 _21732_ (.A1(_04326_),
    .A2(_04336_),
    .Y(_04359_),
    .B1(_04358_));
 sg13g2_and2_1 _21733_ (.A(_04026_),
    .B(_04233_),
    .X(_04360_));
 sg13g2_nand4_1 _21734_ (.B(_04287_),
    .C(net120),
    .A(_04231_),
    .Y(_04361_),
    .D(_04355_));
 sg13g2_nand3_1 _21735_ (.B(_04360_),
    .C(_04361_),
    .A(_04359_),
    .Y(_04362_));
 sg13g2_a221oi_1 _21736_ (.B2(_04116_),
    .C1(_04362_),
    .B1(_04335_),
    .A1(_08844_),
    .Y(_04363_),
    .A2(_04327_));
 sg13g2_a21o_1 _21737_ (.A2(_11638_),
    .A1(net234),
    .B1(_04363_),
    .X(_04364_));
 sg13g2_nand3_1 _21738_ (.B(_08411_),
    .C(_04225_),
    .A(net688),
    .Y(_04365_));
 sg13g2_xor2_1 _21739_ (.B(_04365_),
    .A(_10621_),
    .X(_04366_));
 sg13g2_a22oi_1 _21740_ (.Y(_04367_),
    .B1(_04366_),
    .B2(net76),
    .A2(net33),
    .A1(_08386_));
 sg13g2_o21ai_1 _21741_ (.B1(_04367_),
    .Y(_00986_),
    .A1(_04325_),
    .A2(_04364_));
 sg13g2_a221oi_1 _21742_ (.B2(_11660_),
    .C1(net233),
    .B1(net61),
    .A1(\cpu.ex.r_mult[15] ),
    .Y(_04368_),
    .A2(_10071_));
 sg13g2_xnor2_1 _21743_ (.Y(_04369_),
    .A(_11206_),
    .B(net157));
 sg13g2_buf_1 _21744_ (.A(_04369_),
    .X(_04370_));
 sg13g2_or4_1 _21745_ (.A(_03606_),
    .B(_03678_),
    .C(_04202_),
    .D(_04370_),
    .X(_04371_));
 sg13g2_a21oi_1 _21746_ (.A1(net163),
    .A2(net139),
    .Y(_04372_),
    .B1(_04100_));
 sg13g2_nand2b_1 _21747_ (.Y(_04373_),
    .B(_04372_),
    .A_N(_04370_));
 sg13g2_nand3_1 _21748_ (.B(net163),
    .C(_04370_),
    .A(net1041),
    .Y(_04374_));
 sg13g2_mux2_1 _21749_ (.A0(_04373_),
    .A1(_04374_),
    .S(_03597_),
    .X(_04375_));
 sg13g2_nand3_1 _21750_ (.B(net139),
    .C(_04370_),
    .A(_08842_),
    .Y(_04376_));
 sg13g2_or4_1 _21751_ (.A(_03472_),
    .B(_03584_),
    .C(_03595_),
    .D(_04376_),
    .X(_04377_));
 sg13g2_nor3_1 _21752_ (.A(_03485_),
    .B(_03472_),
    .C(_04376_),
    .Y(_04378_));
 sg13g2_nand2_1 _21753_ (.Y(_04379_),
    .A(net162),
    .B(_03461_));
 sg13g2_o21ai_1 _21754_ (.B1(_11628_),
    .Y(_04380_),
    .A1(_03472_),
    .A2(_03478_));
 sg13g2_nand3_1 _21755_ (.B(_04370_),
    .C(_04380_),
    .A(net139),
    .Y(_04381_));
 sg13g2_o21ai_1 _21756_ (.B1(_04381_),
    .Y(_04382_),
    .A1(_04370_),
    .A2(_04379_));
 sg13g2_nor3_1 _21757_ (.A(net198),
    .B(_04039_),
    .C(_04047_),
    .Y(_04383_));
 sg13g2_nor2_1 _21758_ (.A(_03483_),
    .B(_04178_),
    .Y(_04384_));
 sg13g2_o21ai_1 _21759_ (.B1(net175),
    .Y(_04385_),
    .A1(net178),
    .A2(_04061_));
 sg13g2_a22oi_1 _21760_ (.Y(_04386_),
    .B1(_04186_),
    .B2(_03488_),
    .A2(_04040_),
    .A1(_03468_));
 sg13g2_a22oi_1 _21761_ (.Y(_04387_),
    .B1(_04167_),
    .B2(net199),
    .A2(_04053_),
    .A1(net179));
 sg13g2_nand2_1 _21762_ (.Y(_04388_),
    .A(_04386_),
    .B(_04387_));
 sg13g2_nor4_1 _21763_ (.A(_04383_),
    .B(_04384_),
    .C(_04385_),
    .D(_04388_),
    .Y(_04389_));
 sg13g2_nor2_1 _21764_ (.A(net339),
    .B(_04037_),
    .Y(_04390_));
 sg13g2_or4_1 _21765_ (.A(net244),
    .B(_03525_),
    .C(_03564_),
    .D(_04390_),
    .X(_04391_));
 sg13g2_a22oi_1 _21766_ (.Y(_04392_),
    .B1(_03500_),
    .B2(_04108_),
    .A2(net136),
    .A1(_11021_));
 sg13g2_nand2b_1 _21767_ (.Y(_04393_),
    .B(_03518_),
    .A_N(_04392_));
 sg13g2_nor2_1 _21768_ (.A(_03663_),
    .B(_04307_),
    .Y(_04394_));
 sg13g2_a221oi_1 _21769_ (.B2(_04043_),
    .C1(_04394_),
    .B1(net132),
    .A1(net156),
    .Y(_04395_),
    .A2(_04057_));
 sg13g2_and4_1 _21770_ (.A(_04389_),
    .B(_04391_),
    .C(_04393_),
    .D(_04395_),
    .X(_04396_));
 sg13g2_o21ai_1 _21771_ (.B1(_09744_),
    .Y(_04397_),
    .A1(net141),
    .A2(net175));
 sg13g2_o21ai_1 _21772_ (.B1(_08995_),
    .Y(_04398_),
    .A1(_11206_),
    .A2(net157));
 sg13g2_nand2_1 _21773_ (.Y(_04399_),
    .A(net1099),
    .B(_03680_));
 sg13g2_nand3_1 _21774_ (.B(_04398_),
    .C(_04399_),
    .A(_04193_),
    .Y(_04400_));
 sg13g2_nand2_1 _21775_ (.Y(_04401_),
    .A(_04115_),
    .B(_04370_));
 sg13g2_o21ai_1 _21776_ (.B1(net163),
    .Y(_04402_),
    .A1(net159),
    .A2(_03676_));
 sg13g2_nor2_1 _21777_ (.A(_04401_),
    .B(_04402_),
    .Y(_04403_));
 sg13g2_a221oi_1 _21778_ (.B2(_04400_),
    .C1(_04403_),
    .B1(_03604_),
    .A1(_08891_),
    .Y(_04404_),
    .A2(_11488_));
 sg13g2_o21ai_1 _21779_ (.B1(_04404_),
    .Y(_04405_),
    .A1(_04396_),
    .A2(_04397_));
 sg13g2_a221oi_1 _21780_ (.B2(net1041),
    .C1(_04405_),
    .B1(_04382_),
    .A1(_11564_),
    .Y(_04406_),
    .A2(_04378_));
 sg13g2_nand3_1 _21781_ (.B(_03591_),
    .C(_03474_),
    .A(_11623_),
    .Y(_04407_));
 sg13g2_nand3_1 _21782_ (.B(net141),
    .C(net112),
    .A(_11272_),
    .Y(_04408_));
 sg13g2_a21oi_1 _21783_ (.A1(_04407_),
    .A2(_04408_),
    .Y(_04409_),
    .B1(_04401_));
 sg13g2_nand3_1 _21784_ (.B(_03674_),
    .C(_04409_),
    .A(_03666_),
    .Y(_04410_));
 sg13g2_and4_1 _21785_ (.A(_04360_),
    .B(_04377_),
    .C(_04406_),
    .D(_04410_),
    .X(_04411_));
 sg13g2_nor3_1 _21786_ (.A(_11295_),
    .B(net139),
    .C(_04401_),
    .Y(_04412_));
 sg13g2_o21ai_1 _21787_ (.B1(_04412_),
    .Y(_04413_),
    .A1(_11628_),
    .A2(_04328_));
 sg13g2_a21o_1 _21788_ (.A2(_03674_),
    .A1(_03666_),
    .B1(net112),
    .X(_04414_));
 sg13g2_nand2b_1 _21789_ (.Y(_04415_),
    .B(_04414_),
    .A_N(_04413_));
 sg13g2_and3_1 _21790_ (.X(_04416_),
    .A(_04375_),
    .B(_04411_),
    .C(_04415_));
 sg13g2_a22oi_1 _21791_ (.Y(_04417_),
    .B1(_04371_),
    .B2(_04416_),
    .A2(_04368_),
    .A1(_11658_));
 sg13g2_nand2_1 _21792_ (.Y(_04418_),
    .A(_04024_),
    .B(_04417_));
 sg13g2_or2_1 _21793_ (.X(_04419_),
    .B(_04365_),
    .A(_08599_));
 sg13g2_xnor2_1 _21794_ (.Y(_04420_),
    .A(_03449_),
    .B(_04419_));
 sg13g2_a22oi_1 _21795_ (.Y(_04421_),
    .B1(_04420_),
    .B2(net76),
    .A2(net33),
    .A1(_08379_));
 sg13g2_nand2_1 _21796_ (.Y(_00987_),
    .A(_04418_),
    .B(_04421_));
 sg13g2_nand2_1 _21797_ (.Y(_04422_),
    .A(net245),
    .B(_04026_));
 sg13g2_a22oi_1 _21798_ (.Y(_04423_),
    .B1(_04422_),
    .B2(net318),
    .A2(_11332_),
    .A1(_04064_));
 sg13g2_a22oi_1 _21799_ (.Y(_04424_),
    .B1(net130),
    .B2(net115),
    .A2(_04059_),
    .A1(net159));
 sg13g2_o21ai_1 _21800_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_03663_),
    .A2(_04184_));
 sg13g2_nand2_1 _21801_ (.Y(_04426_),
    .A(net199),
    .B(net133));
 sg13g2_nand2_1 _21802_ (.Y(_04427_),
    .A(net142),
    .B(_04057_));
 sg13g2_a22oi_1 _21803_ (.Y(_04428_),
    .B1(_04253_),
    .B2(_03645_),
    .A2(_04076_),
    .A1(net119));
 sg13g2_nand3_1 _21804_ (.B(_04427_),
    .C(_04428_),
    .A(_04426_),
    .Y(_04429_));
 sg13g2_nand2_1 _21805_ (.Y(_04430_),
    .A(net135),
    .B(net117));
 sg13g2_nand2_1 _21806_ (.Y(_04431_),
    .A(_04043_),
    .B(_04066_));
 sg13g2_a221oi_1 _21807_ (.B2(net137),
    .C1(_04027_),
    .B1(_04167_),
    .A1(_03546_),
    .Y(_04432_),
    .A2(net155));
 sg13g2_nand3_1 _21808_ (.B(_04431_),
    .C(_04432_),
    .A(_04430_),
    .Y(_04433_));
 sg13g2_nor3_1 _21809_ (.A(_04425_),
    .B(_04429_),
    .C(_04433_),
    .Y(_04434_));
 sg13g2_o21ai_1 _21810_ (.B1(_04434_),
    .Y(_04435_),
    .A1(_11315_),
    .A2(_04423_));
 sg13g2_a21oi_1 _21811_ (.A1(_04182_),
    .A2(net84),
    .Y(_04436_),
    .B1(_04092_));
 sg13g2_nand2_1 _21812_ (.Y(_04437_),
    .A(_04435_),
    .B(_04436_));
 sg13g2_nand2_1 _21813_ (.Y(_04438_),
    .A(net209),
    .B(net180));
 sg13g2_a21o_1 _21814_ (.A2(_03614_),
    .A1(net1039),
    .B1(net1022),
    .X(_04439_));
 sg13g2_a22oi_1 _21815_ (.Y(_04440_),
    .B1(net97),
    .B2(net113),
    .A2(net133),
    .A1(net176));
 sg13g2_nor2_1 _21816_ (.A(net209),
    .B(net180),
    .Y(_04441_));
 sg13g2_a221oi_1 _21817_ (.B2(net1021),
    .C1(_11354_),
    .B1(_04441_),
    .A1(net1109),
    .Y(_04442_),
    .A2(net320));
 sg13g2_o21ai_1 _21818_ (.B1(_04442_),
    .Y(_04443_),
    .A1(_04260_),
    .A2(_04440_));
 sg13g2_a21oi_1 _21819_ (.A1(_04438_),
    .A2(_04439_),
    .Y(_04444_),
    .B1(_04443_));
 sg13g2_nor2_1 _21820_ (.A(_09716_),
    .B(_09767_),
    .Y(_04445_));
 sg13g2_nand2_1 _21821_ (.Y(_04446_),
    .A(_04445_),
    .B(_04202_));
 sg13g2_buf_1 _21822_ (.A(_04446_),
    .X(_04447_));
 sg13g2_nand2_1 _21823_ (.Y(_04448_),
    .A(_03614_),
    .B(_04438_));
 sg13g2_xnor2_1 _21824_ (.Y(_04449_),
    .A(_03628_),
    .B(_04448_));
 sg13g2_xor2_1 _21825_ (.B(_04448_),
    .A(_03527_),
    .X(_04450_));
 sg13g2_a22oi_1 _21826_ (.Y(_04451_),
    .B1(_04450_),
    .B2(net1041),
    .A2(_04449_),
    .A1(_04447_));
 sg13g2_nand3_1 _21827_ (.B(_04444_),
    .C(_04451_),
    .A(_04437_),
    .Y(_04452_));
 sg13g2_o21ai_1 _21828_ (.B1(_04452_),
    .Y(_04453_),
    .A1(net233),
    .A2(\cpu.ex.c_mult[2] ));
 sg13g2_a21oi_1 _21829_ (.A1(net913),
    .A2(net83),
    .Y(_04454_),
    .B1(_04136_));
 sg13g2_a21oi_1 _21830_ (.A1(net919),
    .A2(_04127_),
    .Y(_04455_),
    .B1(net798));
 sg13g2_a21oi_1 _21831_ (.A1(net798),
    .A2(_04454_),
    .Y(_04456_),
    .B1(_04455_));
 sg13g2_a21oi_1 _21832_ (.A1(_11344_),
    .A2(_04129_),
    .Y(_04457_),
    .B1(_04456_));
 sg13g2_o21ai_1 _21833_ (.B1(_04457_),
    .Y(_00988_),
    .A1(_04325_),
    .A2(_04453_));
 sg13g2_a21oi_1 _21834_ (.A1(net185),
    .A2(_03500_),
    .Y(_04458_),
    .B1(_11319_));
 sg13g2_nor2_1 _21835_ (.A(net178),
    .B(_04180_),
    .Y(_04459_));
 sg13g2_nor2_1 _21836_ (.A(_03591_),
    .B(_04074_),
    .Y(_04460_));
 sg13g2_nor4_1 _21837_ (.A(_04308_),
    .B(_04383_),
    .C(_04459_),
    .D(_04460_),
    .Y(_04461_));
 sg13g2_a21oi_1 _21838_ (.A1(_04043_),
    .A2(net131),
    .Y(_04462_),
    .B1(_04087_));
 sg13g2_a21oi_1 _21839_ (.A1(net119),
    .A2(_04053_),
    .Y(_04463_),
    .B1(_04179_));
 sg13g2_a22oi_1 _21840_ (.Y(_04464_),
    .B1(_04186_),
    .B2(net140),
    .A2(_04059_),
    .A1(_03455_));
 sg13g2_a22oi_1 _21841_ (.Y(_04465_),
    .B1(_04075_),
    .B2(net136),
    .A2(net130),
    .A1(_03468_));
 sg13g2_and2_1 _21842_ (.A(_04464_),
    .B(_04465_),
    .X(_04466_));
 sg13g2_and4_1 _21843_ (.A(_04461_),
    .B(_04462_),
    .C(_04463_),
    .D(_04466_),
    .X(_04467_));
 sg13g2_o21ai_1 _21844_ (.B1(_04467_),
    .Y(_04468_),
    .A1(net157),
    .A2(_04458_));
 sg13g2_nor2_1 _21845_ (.A(_04153_),
    .B(_04467_),
    .Y(_04469_));
 sg13g2_a21o_1 _21846_ (.A2(_04468_),
    .A1(net1055),
    .B1(_04469_),
    .X(_04470_));
 sg13g2_o21ai_1 _21847_ (.B1(_04470_),
    .Y(_04471_),
    .A1(net199),
    .A2(net175));
 sg13g2_o21ai_1 _21848_ (.B1(_04438_),
    .Y(_04472_),
    .A1(_04441_),
    .A2(_03628_));
 sg13g2_buf_1 _21849_ (.A(_04472_),
    .X(_04473_));
 sg13g2_xnor2_1 _21850_ (.Y(_04474_),
    .A(net316),
    .B(net174));
 sg13g2_xor2_1 _21851_ (.B(_04474_),
    .A(_04473_),
    .X(_04475_));
 sg13g2_nand2_1 _21852_ (.Y(_04476_),
    .A(net245),
    .B(net113));
 sg13g2_a21o_1 _21853_ (.A2(_04476_),
    .A1(_04117_),
    .B1(_11368_),
    .X(_04477_));
 sg13g2_o21ai_1 _21854_ (.B1(_04477_),
    .Y(_04478_),
    .A1(_03498_),
    .A2(_04045_));
 sg13g2_nand3_1 _21855_ (.B(_11021_),
    .C(_04478_),
    .A(net1100),
    .Y(_04479_));
 sg13g2_nor2_1 _21856_ (.A(net316),
    .B(net174),
    .Y(_04480_));
 sg13g2_mux2_1 _21857_ (.A0(net1108),
    .A1(net1099),
    .S(_04480_),
    .X(_04481_));
 sg13g2_nand2_1 _21858_ (.Y(_04482_),
    .A(net316),
    .B(net174));
 sg13g2_o21ai_1 _21859_ (.B1(_04482_),
    .Y(_04483_),
    .A1(_09735_),
    .A2(_04481_));
 sg13g2_a21oi_1 _21860_ (.A1(net1109),
    .A2(net208),
    .Y(_04484_),
    .B1(_11354_));
 sg13g2_nand3_1 _21861_ (.B(_04483_),
    .C(_04484_),
    .A(_04479_),
    .Y(_04485_));
 sg13g2_a21oi_1 _21862_ (.A1(_04447_),
    .A2(_04475_),
    .Y(_04486_),
    .B1(_04485_));
 sg13g2_nor2_1 _21863_ (.A(_03568_),
    .B(_03527_),
    .Y(_04487_));
 sg13g2_a21oi_1 _21864_ (.A1(_03568_),
    .A2(_03527_),
    .Y(_04488_),
    .B1(_11393_));
 sg13g2_nor2_1 _21865_ (.A(_04487_),
    .B(_04488_),
    .Y(_04489_));
 sg13g2_xor2_1 _21866_ (.B(_04489_),
    .A(_04474_),
    .X(_04490_));
 sg13g2_nand2_1 _21867_ (.Y(_04491_),
    .A(net1041),
    .B(_04490_));
 sg13g2_nand3_1 _21868_ (.B(_04486_),
    .C(_04491_),
    .A(_04471_),
    .Y(_04492_));
 sg13g2_o21ai_1 _21869_ (.B1(_04492_),
    .Y(_04493_),
    .A1(net233),
    .A2(\cpu.ex.c_mult[3] ));
 sg13g2_a21o_1 _21870_ (.A2(_04213_),
    .A1(_04127_),
    .B1(_04136_),
    .X(_04494_));
 sg13g2_nor2_1 _21871_ (.A(net690),
    .B(_04213_),
    .Y(_04495_));
 sg13g2_nand2_1 _21872_ (.Y(_04496_),
    .A(_11344_),
    .B(_04129_));
 sg13g2_o21ai_1 _21873_ (.B1(_04133_),
    .Y(_04497_),
    .A1(_00274_),
    .A2(_04496_));
 sg13g2_a221oi_1 _21874_ (.B2(net83),
    .C1(_04497_),
    .B1(_04495_),
    .A1(net690),
    .Y(_04498_),
    .A2(_04494_));
 sg13g2_o21ai_1 _21875_ (.B1(_04498_),
    .Y(_00989_),
    .A1(_04325_),
    .A2(_04493_));
 sg13g2_nor2b_1 _21876_ (.A(_04214_),
    .B_N(net83),
    .Y(_04499_));
 sg13g2_o21ai_1 _21877_ (.B1(net1116),
    .Y(_04500_),
    .A1(_04136_),
    .A2(_04499_));
 sg13g2_buf_1 _21878_ (.A(_09028_),
    .X(_04501_));
 sg13g2_nor3_1 _21879_ (.A(net1111),
    .B(_09182_),
    .C(_11342_),
    .Y(_04502_));
 sg13g2_nor3_1 _21880_ (.A(net918),
    .B(net1116),
    .C(_04213_),
    .Y(_04503_));
 sg13g2_a22oi_1 _21881_ (.Y(_04504_),
    .B1(_04503_),
    .B2(net83),
    .A2(_04502_),
    .A1(net311));
 sg13g2_nor2_1 _21882_ (.A(_03629_),
    .B(_03631_),
    .Y(_04505_));
 sg13g2_nand2_1 _21883_ (.Y(_04506_),
    .A(net312),
    .B(net174));
 sg13g2_nor2_1 _21884_ (.A(net312),
    .B(net174),
    .Y(_04507_));
 sg13g2_a21oi_1 _21885_ (.A1(_04489_),
    .A2(_04506_),
    .Y(_04508_),
    .B1(_04507_));
 sg13g2_xor2_1 _21886_ (.B(_04508_),
    .A(_04505_),
    .X(_04509_));
 sg13g2_o21ai_1 _21887_ (.B1(net1055),
    .Y(_04510_),
    .A1(_11319_),
    .A2(_03500_));
 sg13g2_a21oi_1 _21888_ (.A1(_04074_),
    .A2(_04510_),
    .Y(_04511_),
    .B1(net157));
 sg13g2_a21oi_1 _21889_ (.A1(_03546_),
    .A2(_04164_),
    .Y(_04512_),
    .B1(_04087_));
 sg13g2_o21ai_1 _21890_ (.B1(_04512_),
    .Y(_04513_),
    .A1(_03483_),
    .A2(_04310_));
 sg13g2_a22oi_1 _21891_ (.Y(_04514_),
    .B1(_04053_),
    .B2(net136),
    .A2(_04075_),
    .A1(_03468_));
 sg13g2_a22oi_1 _21892_ (.Y(_04515_),
    .B1(_04081_),
    .B2(net140),
    .A2(net130),
    .A1(net159));
 sg13g2_nand2_1 _21893_ (.Y(_04516_),
    .A(_04514_),
    .B(_04515_));
 sg13g2_nor3_1 _21894_ (.A(_04511_),
    .B(_04513_),
    .C(_04516_),
    .Y(_04517_));
 sg13g2_a221oi_1 _21895_ (.B2(net135),
    .C1(_04345_),
    .B1(_04066_),
    .A1(_04043_),
    .Y(_04518_),
    .A2(net133));
 sg13g2_nand2_1 _21896_ (.Y(_04519_),
    .A(_04517_),
    .B(_04518_));
 sg13g2_a21oi_1 _21897_ (.A1(_03549_),
    .A2(net116),
    .Y(_04520_),
    .B1(_04092_));
 sg13g2_nand2_1 _21898_ (.Y(_04521_),
    .A(net156),
    .B(_04040_));
 sg13g2_nand2_1 _21899_ (.Y(_04522_),
    .A(_04108_),
    .B(_04066_));
 sg13g2_a21oi_1 _21900_ (.A1(_04172_),
    .A2(_04164_),
    .Y(_04523_),
    .B1(_04087_));
 sg13g2_nand3_1 _21901_ (.B(_04522_),
    .C(_04523_),
    .A(_04521_),
    .Y(_04524_));
 sg13g2_a21oi_1 _21902_ (.A1(net174),
    .A2(_04087_),
    .Y(_04525_),
    .B1(_04260_));
 sg13g2_a221oi_1 _21903_ (.B2(_04525_),
    .C1(_04115_),
    .B1(_04524_),
    .A1(net1109),
    .Y(_04526_),
    .A2(_03955_));
 sg13g2_mux2_1 _21904_ (.A0(net1108),
    .A1(net1099),
    .S(_03631_),
    .X(_04527_));
 sg13g2_o21ai_1 _21905_ (.B1(_03617_),
    .Y(_04528_),
    .A1(_09735_),
    .A2(_04527_));
 sg13g2_nand2_1 _21906_ (.Y(_04529_),
    .A(_04526_),
    .B(_04528_));
 sg13g2_a221oi_1 _21907_ (.B2(_04520_),
    .C1(_04529_),
    .B1(_04519_),
    .A1(net1041),
    .Y(_04530_),
    .A2(_04509_));
 sg13g2_nor2_1 _21908_ (.A(net582),
    .B(_04530_),
    .Y(_04531_));
 sg13g2_o21ai_1 _21909_ (.B1(net316),
    .Y(_04532_),
    .A1(net174),
    .A2(_04473_));
 sg13g2_nand2_1 _21910_ (.Y(_04533_),
    .A(net174),
    .B(_04473_));
 sg13g2_nand2_1 _21911_ (.Y(_04534_),
    .A(_04532_),
    .B(_04533_));
 sg13g2_xor2_1 _21912_ (.B(_04505_),
    .A(_04534_),
    .X(_04535_));
 sg13g2_a21oi_1 _21913_ (.A1(_04445_),
    .A2(_04530_),
    .Y(_04536_),
    .B1(_04535_));
 sg13g2_nor2_1 _21914_ (.A(_04531_),
    .B(_04536_),
    .Y(_04537_));
 sg13g2_nor2_1 _21915_ (.A(_04266_),
    .B(\cpu.ex.c_mult[4] ),
    .Y(_04538_));
 sg13g2_a21oi_1 _21916_ (.A1(_04318_),
    .A2(_04537_),
    .Y(_04539_),
    .B1(_04538_));
 sg13g2_nand2_1 _21917_ (.Y(_04540_),
    .A(net85),
    .B(_04539_));
 sg13g2_nand3_1 _21918_ (.B(_04504_),
    .C(_04540_),
    .A(_04500_),
    .Y(_00990_));
 sg13g2_nand2_1 _21919_ (.Y(_04541_),
    .A(net243),
    .B(net178));
 sg13g2_nand2b_1 _21920_ (.Y(_04542_),
    .B(_04541_),
    .A_N(_03633_));
 sg13g2_xnor2_1 _21921_ (.Y(_04543_),
    .A(_03572_),
    .B(_04542_));
 sg13g2_xnor2_1 _21922_ (.Y(_04544_),
    .A(_04146_),
    .B(_04542_));
 sg13g2_or2_1 _21923_ (.X(_04545_),
    .B(_09714_),
    .A(_08358_));
 sg13g2_buf_1 _21924_ (.A(_04545_),
    .X(_04546_));
 sg13g2_a22oi_1 _21925_ (.Y(_04547_),
    .B1(net117),
    .B2(net119),
    .A2(net132),
    .A1(net141));
 sg13g2_nor2_1 _21926_ (.A(_03534_),
    .B(_04180_),
    .Y(_04548_));
 sg13g2_a21oi_1 _21927_ (.A1(net112),
    .A2(net118),
    .Y(_04549_),
    .B1(_04548_));
 sg13g2_a21oi_1 _21928_ (.A1(_03645_),
    .A2(_04066_),
    .Y(_04550_),
    .B1(_04394_));
 sg13g2_nor2_1 _21929_ (.A(_11313_),
    .B(_04030_),
    .Y(_04551_));
 sg13g2_and2_1 _21930_ (.A(net1055),
    .B(_03455_),
    .X(_04552_));
 sg13g2_o21ai_1 _21931_ (.B1(_04552_),
    .Y(_04553_),
    .A1(_11319_),
    .A2(_04551_));
 sg13g2_a22oi_1 _21932_ (.Y(_04554_),
    .B1(net129),
    .B2(net136),
    .A2(_04174_),
    .A1(_03455_));
 sg13g2_and4_1 _21933_ (.A(_04166_),
    .B(_04550_),
    .C(_04553_),
    .D(_04554_),
    .X(_04555_));
 sg13g2_nand3_1 _21934_ (.B(_04549_),
    .C(_04555_),
    .A(_04547_),
    .Y(_04556_));
 sg13g2_nand2_1 _21935_ (.Y(_04557_),
    .A(_10518_),
    .B(net97));
 sg13g2_nand3_1 _21936_ (.B(_04556_),
    .C(_04557_),
    .A(_04546_),
    .Y(_04558_));
 sg13g2_mux2_1 _21937_ (.A0(net1039),
    .A1(net1021),
    .S(_03633_),
    .X(_04559_));
 sg13g2_o21ai_1 _21938_ (.B1(_04541_),
    .Y(_04560_),
    .A1(net1022),
    .A2(_04559_));
 sg13g2_a22oi_1 _21939_ (.Y(_04561_),
    .B1(_04252_),
    .B2(_04108_),
    .A2(net114),
    .A1(net113));
 sg13g2_a21oi_1 _21940_ (.A1(net156),
    .A2(net131),
    .Y(_04562_),
    .B1(net116));
 sg13g2_nand3_1 _21941_ (.B(_04561_),
    .C(_04562_),
    .A(_04042_),
    .Y(_04563_));
 sg13g2_a21oi_1 _21942_ (.A1(_10492_),
    .A2(net97),
    .Y(_04564_),
    .B1(_04260_));
 sg13g2_a221oi_1 _21943_ (.B2(_04564_),
    .C1(_11354_),
    .B1(_04563_),
    .A1(net1040),
    .Y(_04565_),
    .A2(_11271_));
 sg13g2_nand3_1 _21944_ (.B(_04560_),
    .C(_04565_),
    .A(_04558_),
    .Y(_04566_));
 sg13g2_a221oi_1 _21945_ (.B2(_04447_),
    .C1(_04566_),
    .B1(_04544_),
    .A1(net1041),
    .Y(_04567_),
    .A2(_04543_));
 sg13g2_a21oi_1 _21946_ (.A1(net234),
    .A2(_11455_),
    .Y(_04568_),
    .B1(_04567_));
 sg13g2_nand2_1 _21947_ (.Y(_04569_),
    .A(net85),
    .B(_04568_));
 sg13g2_buf_1 _21948_ (.A(_08701_),
    .X(_04570_));
 sg13g2_xnor2_1 _21949_ (.Y(_04571_),
    .A(_10399_),
    .B(_04216_));
 sg13g2_a22oi_1 _21950_ (.Y(_04572_),
    .B1(_04571_),
    .B2(_04223_),
    .A2(_04137_),
    .A1(net947));
 sg13g2_nand2_1 _21951_ (.Y(_00991_),
    .A(_04569_),
    .B(_04572_));
 sg13g2_nand2_1 _21952_ (.Y(_04573_),
    .A(_11458_),
    .B(_11467_));
 sg13g2_a221oi_1 _21953_ (.B2(net542),
    .C1(_04318_),
    .B1(_04573_),
    .A1(\cpu.ex.r_mult[6] ),
    .Y(_04574_),
    .A2(net374));
 sg13g2_inv_1 _21954_ (.Y(_04575_),
    .A(_03634_));
 sg13g2_nand2_1 _21955_ (.Y(_04576_),
    .A(_03635_),
    .B(_04575_));
 sg13g2_nor2_1 _21956_ (.A(net178),
    .B(_03572_),
    .Y(_04577_));
 sg13g2_a21oi_1 _21957_ (.A1(net178),
    .A2(_03572_),
    .Y(_04578_),
    .B1(_11442_));
 sg13g2_nor2_1 _21958_ (.A(_04577_),
    .B(_04578_),
    .Y(_04579_));
 sg13g2_xnor2_1 _21959_ (.Y(_04580_),
    .A(_04576_),
    .B(_04579_));
 sg13g2_a21oi_1 _21960_ (.A1(_04146_),
    .A2(_04541_),
    .Y(_04581_),
    .B1(_03633_));
 sg13g2_xor2_1 _21961_ (.B(_04576_),
    .A(_04581_),
    .X(_04582_));
 sg13g2_a22oi_1 _21962_ (.Y(_04583_),
    .B1(net132),
    .B2(net142),
    .A2(net133),
    .A1(_04028_));
 sg13g2_a22oi_1 _21963_ (.Y(_04584_),
    .B1(net129),
    .B2(_03608_),
    .A2(_04054_),
    .A1(_03460_));
 sg13g2_o21ai_1 _21964_ (.B1(_04339_),
    .Y(_04585_),
    .A1(net138),
    .A2(_04307_));
 sg13g2_a21oi_1 _21965_ (.A1(net115),
    .A2(net117),
    .Y(_04586_),
    .B1(_04585_));
 sg13g2_nand4_1 _21966_ (.B(_04583_),
    .C(_04584_),
    .A(_04256_),
    .Y(_04587_),
    .D(_04586_));
 sg13g2_nand2_1 _21967_ (.Y(_04588_),
    .A(_04546_),
    .B(_04587_));
 sg13g2_a22oi_1 _21968_ (.Y(_04589_),
    .B1(_04553_),
    .B2(_04588_),
    .A2(net84),
    .A1(_03534_));
 sg13g2_nand2_1 _21969_ (.Y(_04590_),
    .A(net1039),
    .B(_04575_));
 sg13g2_nand2_1 _21970_ (.Y(_04591_),
    .A(net1021),
    .B(_03634_));
 sg13g2_nand3_1 _21971_ (.B(_04590_),
    .C(_04591_),
    .A(_04193_),
    .Y(_04592_));
 sg13g2_nand2_1 _21972_ (.Y(_04593_),
    .A(net134),
    .B(net131));
 sg13g2_a22oi_1 _21973_ (.Y(_04594_),
    .B1(_04252_),
    .B2(net113),
    .A2(_04154_),
    .A1(net156));
 sg13g2_a21oi_1 _21974_ (.A1(net176),
    .A2(net117),
    .Y(_04595_),
    .B1(_04089_));
 sg13g2_nand4_1 _21975_ (.B(_04593_),
    .C(_04594_),
    .A(_04426_),
    .Y(_04596_),
    .D(_04595_));
 sg13g2_a21oi_1 _21976_ (.A1(net178),
    .A2(net84),
    .Y(_04597_),
    .B1(_04260_));
 sg13g2_a22oi_1 _21977_ (.Y(_04598_),
    .B1(_04596_),
    .B2(_04597_),
    .A2(_04592_),
    .A1(_03635_));
 sg13g2_a21oi_1 _21978_ (.A1(net1040),
    .A2(_11623_),
    .Y(_04599_),
    .B1(net234));
 sg13g2_nand3b_1 _21979_ (.B(_04598_),
    .C(_04599_),
    .Y(_04600_),
    .A_N(_04589_));
 sg13g2_a221oi_1 _21980_ (.B2(_04447_),
    .C1(_04600_),
    .B1(_04582_),
    .A1(net901),
    .Y(_04601_),
    .A2(_04580_));
 sg13g2_nor3_1 _21981_ (.A(_04325_),
    .B(_04574_),
    .C(_04601_),
    .Y(_04602_));
 sg13g2_nand2_1 _21982_ (.Y(_04603_),
    .A(_08701_),
    .B(_04216_));
 sg13g2_xor2_1 _21983_ (.B(_04603_),
    .A(_00295_),
    .X(_04604_));
 sg13g2_a22oi_1 _21984_ (.Y(_04605_),
    .B1(_04604_),
    .B2(net76),
    .A2(net33),
    .A1(_08669_));
 sg13g2_nand2b_1 _21985_ (.Y(_00992_),
    .B(_04605_),
    .A_N(_04602_));
 sg13g2_nor2_1 _21986_ (.A(_04043_),
    .B(net321),
    .Y(_04606_));
 sg13g2_o21ai_1 _21987_ (.B1(_03536_),
    .Y(_04607_),
    .A1(_04606_),
    .A2(_04579_));
 sg13g2_xor2_1 _21988_ (.B(_04607_),
    .A(_04144_),
    .X(_04608_));
 sg13g2_nand2_1 _21989_ (.Y(_04609_),
    .A(_10717_),
    .B(net84));
 sg13g2_o21ai_1 _21990_ (.B1(_04026_),
    .Y(_04610_),
    .A1(_03798_),
    .A2(net245));
 sg13g2_o21ai_1 _21991_ (.B1(_04610_),
    .Y(_04611_),
    .A1(_03798_),
    .A2(_04030_));
 sg13g2_nor2_1 _21992_ (.A(_04301_),
    .B(_04384_),
    .Y(_04612_));
 sg13g2_a21oi_1 _21993_ (.A1(net115),
    .A2(_04048_),
    .Y(_04613_),
    .B1(_04181_));
 sg13g2_nand3_1 _21994_ (.B(_04612_),
    .C(_04613_),
    .A(_04611_),
    .Y(_04614_));
 sg13g2_a221oi_1 _21995_ (.B2(net141),
    .C1(_04614_),
    .B1(net129),
    .A1(net112),
    .Y(_04615_),
    .A2(net117));
 sg13g2_nand2_1 _21996_ (.Y(_04616_),
    .A(_04054_),
    .B(_04351_));
 sg13g2_o21ai_1 _21997_ (.B1(_04616_),
    .Y(_04617_),
    .A1(_04092_),
    .A2(_04615_));
 sg13g2_a21oi_1 _21998_ (.A1(net134),
    .A2(net114),
    .Y(_04618_),
    .B1(net116));
 sg13g2_a22oi_1 _21999_ (.Y(_04619_),
    .B1(net129),
    .B2(_04108_),
    .A2(net155),
    .A1(net156));
 sg13g2_a221oi_1 _22000_ (.B2(net199),
    .C1(_04459_),
    .B1(net131),
    .A1(net113),
    .Y(_04620_),
    .A2(_04081_));
 sg13g2_nand3_1 _22001_ (.B(_04619_),
    .C(_04620_),
    .A(_04618_),
    .Y(_04621_));
 sg13g2_nand3_1 _22002_ (.B(_04557_),
    .C(_04621_),
    .A(net1100),
    .Y(_04622_));
 sg13g2_a21oi_1 _22003_ (.A1(net1109),
    .A2(_11207_),
    .Y(_04623_),
    .B1(_11354_));
 sg13g2_mux2_1 _22004_ (.A0(net1099),
    .A1(net1108),
    .S(_03637_),
    .X(_04624_));
 sg13g2_o21ai_1 _22005_ (.B1(_04142_),
    .Y(_04625_),
    .A1(net1022),
    .A2(_04624_));
 sg13g2_nand3_1 _22006_ (.B(_04623_),
    .C(_04625_),
    .A(_04622_),
    .Y(_04626_));
 sg13g2_a221oi_1 _22007_ (.B2(_04617_),
    .C1(_04626_),
    .B1(_04609_),
    .A1(_04148_),
    .Y(_04627_),
    .A2(_04447_));
 sg13g2_o21ai_1 _22008_ (.B1(_04627_),
    .Y(_04628_),
    .A1(_04100_),
    .A2(_04608_));
 sg13g2_o21ai_1 _22009_ (.B1(_04628_),
    .Y(_04629_),
    .A1(net233),
    .A2(\cpu.ex.c_mult[7] ));
 sg13g2_xor2_1 _22010_ (.B(_04217_),
    .A(_10398_),
    .X(_04630_));
 sg13g2_a22oi_1 _22011_ (.Y(_04631_),
    .B1(_04630_),
    .B2(net76),
    .A2(_04136_),
    .A1(\cpu.ex.pc[7] ));
 sg13g2_o21ai_1 _22012_ (.B1(_04631_),
    .Y(_00993_),
    .A1(_04325_),
    .A2(_04629_));
 sg13g2_a22oi_1 _22013_ (.Y(_04632_),
    .B1(net129),
    .B2(net142),
    .A2(net114),
    .A1(net115));
 sg13g2_o21ai_1 _22014_ (.B1(_04247_),
    .Y(_04633_),
    .A1(net138),
    .A2(_04079_));
 sg13g2_a221oi_1 _22015_ (.B2(net141),
    .C1(_04633_),
    .B1(net117),
    .A1(net137),
    .Y(_04634_),
    .A2(net155));
 sg13g2_nand3_1 _22016_ (.B(_04632_),
    .C(_04634_),
    .A(_04611_),
    .Y(_04635_));
 sg13g2_a21oi_1 _22017_ (.A1(net198),
    .A2(net97),
    .Y(_04636_),
    .B1(_04092_));
 sg13g2_a21oi_1 _22018_ (.A1(_03561_),
    .A2(_03572_),
    .Y(_04637_),
    .B1(_03573_));
 sg13g2_nand2_1 _22019_ (.Y(_04638_),
    .A(_10717_),
    .B(net211));
 sg13g2_nand2_1 _22020_ (.Y(_04639_),
    .A(_03488_),
    .B(_11125_));
 sg13g2_nand2_1 _22021_ (.Y(_04640_),
    .A(_04638_),
    .B(_04639_));
 sg13g2_xor2_1 _22022_ (.B(_04640_),
    .A(_04637_),
    .X(_04641_));
 sg13g2_nor2_1 _22023_ (.A(_10492_),
    .B(_04178_),
    .Y(_04642_));
 sg13g2_a221oi_1 _22024_ (.B2(_04108_),
    .C1(_04642_),
    .B1(net118),
    .A1(net156),
    .Y(_04643_),
    .A2(_04081_));
 sg13g2_nand2_1 _22025_ (.Y(_04644_),
    .A(_04172_),
    .B(_04186_));
 sg13g2_o21ai_1 _22026_ (.B1(_04644_),
    .Y(_04645_),
    .A1(_10518_),
    .A2(_04180_));
 sg13g2_a221oi_1 _22027_ (.B2(_04064_),
    .C1(_04645_),
    .B1(net131),
    .A1(net134),
    .Y(_04646_),
    .A2(net155));
 sg13g2_and3_1 _22028_ (.X(_04647_),
    .A(net175),
    .B(_04643_),
    .C(_04646_));
 sg13g2_o21ai_1 _22029_ (.B1(net1100),
    .Y(_04648_),
    .A1(net179),
    .A2(net175));
 sg13g2_nand3_1 _22030_ (.B(net135),
    .C(_11499_),
    .A(net1099),
    .Y(_04649_));
 sg13g2_nand2_1 _22031_ (.Y(_04650_),
    .A(net1108),
    .B(_04639_));
 sg13g2_nand3_1 _22032_ (.B(_04649_),
    .C(_04650_),
    .A(_04193_),
    .Y(_04651_));
 sg13g2_a22oi_1 _22033_ (.Y(_04652_),
    .B1(_04638_),
    .B2(_04651_),
    .A2(_11332_),
    .A1(net1109));
 sg13g2_o21ai_1 _22034_ (.B1(_04652_),
    .Y(_04653_),
    .A1(_04647_),
    .A2(_04648_));
 sg13g2_a221oi_1 _22035_ (.B2(net1041),
    .C1(_04653_),
    .B1(_04641_),
    .A1(_04635_),
    .Y(_04654_),
    .A2(_04636_));
 sg13g2_nand2_1 _22036_ (.Y(_04655_),
    .A(_03638_),
    .B(_03642_));
 sg13g2_xnor2_1 _22037_ (.Y(_04656_),
    .A(_04655_),
    .B(_04640_));
 sg13g2_a22oi_1 _22038_ (.Y(_04657_),
    .B1(_04656_),
    .B2(net582),
    .A2(_04654_),
    .A1(_04149_));
 sg13g2_mux2_1 _22039_ (.A0(\cpu.ex.c_mult[8] ),
    .A1(_04657_),
    .S(_04266_),
    .X(_04658_));
 sg13g2_nand2_1 _22040_ (.Y(_04659_),
    .A(net85),
    .B(_04658_));
 sg13g2_xor2_1 _22041_ (.B(_04219_),
    .A(_10695_),
    .X(_04660_));
 sg13g2_a22oi_1 _22042_ (.Y(_04661_),
    .B1(_04660_),
    .B2(net76),
    .A2(net33),
    .A1(\cpu.ex.pc[8] ));
 sg13g2_nand2_1 _22043_ (.Y(_00994_),
    .A(_04659_),
    .B(_04661_));
 sg13g2_xnor2_1 _22044_ (.Y(_04662_),
    .A(_10626_),
    .B(_04220_));
 sg13g2_a22oi_1 _22045_ (.Y(_04663_),
    .B1(_04662_),
    .B2(net76),
    .A2(net33),
    .A1(_08719_));
 sg13g2_and2_1 _22046_ (.A(net135),
    .B(_03552_),
    .X(_04664_));
 sg13g2_nor2_1 _22047_ (.A(_04664_),
    .B(_03575_),
    .Y(_04665_));
 sg13g2_nand2_1 _22048_ (.Y(_04666_),
    .A(_03651_),
    .B(_03646_));
 sg13g2_xnor2_1 _22049_ (.Y(_04667_),
    .A(_04665_),
    .B(_04666_));
 sg13g2_a22oi_1 _22050_ (.Y(_04668_),
    .B1(_04165_),
    .B2(net115),
    .A2(_04082_),
    .A1(net142));
 sg13g2_a22oi_1 _22051_ (.Y(_04669_),
    .B1(net155),
    .B2(net141),
    .A2(net114),
    .A1(_03608_));
 sg13g2_and2_1 _22052_ (.A(_04668_),
    .B(_04669_),
    .X(_04670_));
 sg13g2_o21ai_1 _22053_ (.B1(_11402_),
    .Y(_04671_),
    .A1(_11383_),
    .A2(net185));
 sg13g2_nor3_1 _22054_ (.A(_11393_),
    .B(net318),
    .C(_11316_),
    .Y(_04672_));
 sg13g2_o21ai_1 _22055_ (.B1(_04552_),
    .Y(_04673_),
    .A1(_04671_),
    .A2(_04672_));
 sg13g2_nand4_1 _22056_ (.B(_04300_),
    .C(_04670_),
    .A(net175),
    .Y(_04674_),
    .D(_04673_));
 sg13g2_nand3_1 _22057_ (.B(_04191_),
    .C(_04674_),
    .A(_04546_),
    .Y(_04675_));
 sg13g2_mux2_1 _22058_ (.A0(net1021),
    .A1(net1039),
    .S(_03646_),
    .X(_04676_));
 sg13g2_o21ai_1 _22059_ (.B1(_03651_),
    .Y(_04677_),
    .A1(net1022),
    .A2(_04676_));
 sg13g2_a21oi_1 _22060_ (.A1(net1040),
    .A2(net339),
    .Y(_04678_),
    .B1(net582));
 sg13g2_a22oi_1 _22061_ (.Y(_04679_),
    .B1(_04253_),
    .B2(net156),
    .A2(net117),
    .A1(_04037_));
 sg13g2_a22oi_1 _22062_ (.Y(_04680_),
    .B1(net118),
    .B2(_04257_),
    .A2(net155),
    .A1(net199));
 sg13g2_a221oi_1 _22063_ (.B2(_04109_),
    .C1(_04548_),
    .B1(_04076_),
    .A1(_04064_),
    .Y(_04681_),
    .A2(_04154_));
 sg13g2_nand4_1 _22064_ (.B(_04679_),
    .C(_04680_),
    .A(_04462_),
    .Y(_04682_),
    .D(_04681_));
 sg13g2_nand3_1 _22065_ (.B(_04609_),
    .C(_04682_),
    .A(net1100),
    .Y(_04683_));
 sg13g2_nand4_1 _22066_ (.B(_04677_),
    .C(_04678_),
    .A(_04675_),
    .Y(_04684_),
    .D(_04683_));
 sg13g2_a21oi_1 _22067_ (.A1(net901),
    .A2(_04667_),
    .Y(_04685_),
    .B1(_04684_));
 sg13g2_nand2_1 _22068_ (.Y(_04686_),
    .A(_04025_),
    .B(\cpu.ex.c_mult[9] ));
 sg13g2_nand2_1 _22069_ (.Y(_04687_),
    .A(_11095_),
    .B(_04655_));
 sg13g2_o21ai_1 _22070_ (.B1(_10717_),
    .Y(_04688_),
    .A1(_11095_),
    .A2(_04655_));
 sg13g2_nand2_1 _22071_ (.Y(_04689_),
    .A(_04687_),
    .B(_04688_));
 sg13g2_xor2_1 _22072_ (.B(_04666_),
    .A(_04689_),
    .X(_04690_));
 sg13g2_o21ai_1 _22073_ (.B1(net233),
    .Y(_04691_),
    .A1(_04202_),
    .A2(_04690_));
 sg13g2_a22oi_1 _22074_ (.Y(_04692_),
    .B1(_04686_),
    .B2(_04691_),
    .A2(_04685_),
    .A1(_04233_));
 sg13g2_nand2_1 _22075_ (.Y(_04693_),
    .A(net85),
    .B(_04692_));
 sg13g2_nand2_1 _22076_ (.Y(_00995_),
    .A(_04663_),
    .B(_04693_));
 sg13g2_o21ai_1 _22077_ (.B1(_03579_),
    .Y(_04694_),
    .A1(_04664_),
    .A2(_03575_));
 sg13g2_o21ai_1 _22078_ (.B1(_04694_),
    .Y(_04695_),
    .A1(_03559_),
    .A2(net186));
 sg13g2_and2_1 _22079_ (.A(_04203_),
    .B(_04204_),
    .X(_04696_));
 sg13g2_xnor2_1 _22080_ (.Y(_04697_),
    .A(_04695_),
    .B(_04696_));
 sg13g2_nor2_1 _22081_ (.A(_03650_),
    .B(_03653_),
    .Y(_04698_));
 sg13g2_xor2_1 _22082_ (.B(_04696_),
    .A(_04698_),
    .X(_04699_));
 sg13g2_a22oi_1 _22083_ (.Y(_04700_),
    .B1(net155),
    .B2(_04064_),
    .A2(net132),
    .A1(_04257_));
 sg13g2_o21ai_1 _22084_ (.B1(_04431_),
    .Y(_04701_),
    .A1(_10717_),
    .A2(_04180_));
 sg13g2_a221oi_1 _22085_ (.B2(net134),
    .C1(_04701_),
    .B1(net129),
    .A1(_04109_),
    .Y(_04702_),
    .A2(net130));
 sg13g2_a22oi_1 _22086_ (.Y(_04703_),
    .B1(net118),
    .B2(_04249_),
    .A2(_04082_),
    .A1(_03505_));
 sg13g2_nand4_1 _22087_ (.B(_04700_),
    .C(_04702_),
    .A(_04512_),
    .Y(_04704_),
    .D(_04703_));
 sg13g2_a21oi_1 _22088_ (.A1(net198),
    .A2(net84),
    .Y(_04705_),
    .B1(_04260_));
 sg13g2_nand2_1 _22089_ (.Y(_04706_),
    .A(_04704_),
    .B(_04705_));
 sg13g2_mux2_1 _22090_ (.A0(net1021),
    .A1(net1039),
    .S(_04204_),
    .X(_04707_));
 sg13g2_o21ai_1 _22091_ (.B1(_04203_),
    .Y(_04708_),
    .A1(net1022),
    .A2(_04707_));
 sg13g2_o21ai_1 _22092_ (.B1(net1055),
    .Y(_04709_),
    .A1(_04029_),
    .A2(_04671_));
 sg13g2_a21o_1 _22093_ (.A2(_04709_),
    .A1(_04307_),
    .B1(_03603_),
    .X(_04710_));
 sg13g2_a22oi_1 _22094_ (.Y(_04711_),
    .B1(net114),
    .B2(net141),
    .A2(_04041_),
    .A1(_04150_));
 sg13g2_a21oi_1 _22095_ (.A1(net112),
    .A2(net131),
    .Y(_04712_),
    .B1(net97));
 sg13g2_nand3_1 _22096_ (.B(_04711_),
    .C(_04712_),
    .A(_04710_),
    .Y(_04713_));
 sg13g2_a21oi_1 _22097_ (.A1(net138),
    .A2(net97),
    .Y(_04714_),
    .B1(_04092_));
 sg13g2_a22oi_1 _22098_ (.Y(_04715_),
    .B1(_04713_),
    .B2(_04714_),
    .A2(_11383_),
    .A1(net1040));
 sg13g2_nand4_1 _22099_ (.B(_04706_),
    .C(_04708_),
    .A(_04233_),
    .Y(_04716_),
    .D(_04715_));
 sg13g2_a221oi_1 _22100_ (.B2(net582),
    .C1(_04716_),
    .B1(_04699_),
    .A1(net901),
    .Y(_04717_),
    .A2(_04697_));
 sg13g2_a21oi_1 _22101_ (.A1(_04025_),
    .A2(_11551_),
    .Y(_04718_),
    .B1(_04717_));
 sg13g2_nand2_1 _22102_ (.Y(_04719_),
    .A(net85),
    .B(_04718_));
 sg13g2_buf_1 _22103_ (.A(_08710_),
    .X(_04720_));
 sg13g2_nand2_1 _22104_ (.Y(_04721_),
    .A(_08719_),
    .B(_04220_));
 sg13g2_xor2_1 _22105_ (.B(_04721_),
    .A(_10651_),
    .X(_04722_));
 sg13g2_a22oi_1 _22106_ (.Y(_04723_),
    .B1(_04722_),
    .B2(net76),
    .A2(net33),
    .A1(net946));
 sg13g2_nand2_1 _22107_ (.Y(_00996_),
    .A(_04719_),
    .B(_04723_));
 sg13g2_mux2_1 _22108_ (.A0(\cpu.dec.r_set_cc ),
    .A1(_10062_),
    .S(_03448_),
    .X(_00999_));
 sg13g2_buf_1 _22109_ (.A(_00256_),
    .X(_04724_));
 sg13g2_nor4_1 _22110_ (.A(net1096),
    .B(_10057_),
    .C(_04724_),
    .D(_03380_),
    .Y(_04725_));
 sg13g2_buf_2 _22111_ (.A(_04725_),
    .X(_04726_));
 sg13g2_buf_1 _22112_ (.A(_04726_),
    .X(_04727_));
 sg13g2_mux2_1 _22113_ (.A0(_10318_),
    .A1(net544),
    .S(net517),
    .X(_01000_));
 sg13g2_mux2_1 _22114_ (.A0(_10118_),
    .A1(net949),
    .S(net517),
    .X(_01001_));
 sg13g2_mux2_1 _22115_ (.A0(_10527_),
    .A1(net529),
    .S(net517),
    .X(_01002_));
 sg13g2_mux2_1 _22116_ (.A0(_10579_),
    .A1(net468),
    .S(_04727_),
    .X(_01003_));
 sg13g2_mux2_1 _22117_ (.A0(_10554_),
    .A1(net524),
    .S(net517),
    .X(_01004_));
 sg13g2_mux2_1 _22118_ (.A0(_10602_),
    .A1(net641),
    .S(net517),
    .X(_01005_));
 sg13g2_mux2_1 _22119_ (.A0(_10386_),
    .A1(net406),
    .S(_04727_),
    .X(_01006_));
 sg13g2_mux2_1 _22120_ (.A0(_10246_),
    .A1(net405),
    .S(net517),
    .X(_01007_));
 sg13g2_mux2_1 _22121_ (.A0(_10462_),
    .A1(net314),
    .S(net517),
    .X(_01008_));
 sg13g2_mux2_1 _22122_ (.A0(_10448_),
    .A1(net591),
    .S(net517),
    .X(_01009_));
 sg13g2_mux2_1 _22123_ (.A0(_10511_),
    .A1(net840),
    .S(_04726_),
    .X(_01010_));
 sg13g2_mux2_1 _22124_ (.A0(_10406_),
    .A1(net716),
    .S(_04726_),
    .X(_01011_));
 sg13g2_mux2_1 _22125_ (.A0(_10697_),
    .A1(net715),
    .S(_04726_),
    .X(_01012_));
 sg13g2_mux2_1 _22126_ (.A0(_10629_),
    .A1(net839),
    .S(_04726_),
    .X(_01013_));
 sg13g2_mux2_1 _22127_ (.A0(_10662_),
    .A1(net838),
    .S(_04726_),
    .X(_01014_));
 sg13g2_or2_1 _22128_ (.X(_04728_),
    .B(_03380_),
    .A(_03752_));
 sg13g2_buf_1 _22129_ (.A(_04728_),
    .X(_04729_));
 sg13g2_buf_1 _22130_ (.A(_04729_),
    .X(_04730_));
 sg13g2_nor2b_1 _22131_ (.A(_04724_),
    .B_N(net911),
    .Y(_04731_));
 sg13g2_nand2_1 _22132_ (.Y(_04732_),
    .A(_03378_),
    .B(_04731_));
 sg13g2_and2_1 _22133_ (.A(net911),
    .B(_10057_),
    .X(_04733_));
 sg13g2_a21oi_1 _22134_ (.A1(_10058_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04734_),
    .B1(_04733_));
 sg13g2_or4_1 _22135_ (.A(net1096),
    .B(_04724_),
    .C(_03380_),
    .D(_04734_),
    .X(_04735_));
 sg13g2_buf_1 _22136_ (.A(_04735_),
    .X(_04736_));
 sg13g2_buf_1 _22137_ (.A(_04736_),
    .X(_04737_));
 sg13g2_nand2_1 _22138_ (.Y(_04738_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net466));
 sg13g2_o21ai_1 _22139_ (.B1(_04738_),
    .Y(_01015_),
    .A1(_04730_),
    .A2(_04732_));
 sg13g2_mux2_1 _22140_ (.A0(net1089),
    .A1(_10662_),
    .S(net516),
    .X(_04739_));
 sg13g2_buf_1 _22141_ (.A(_04736_),
    .X(_04740_));
 sg13g2_mux2_1 _22142_ (.A0(_04739_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net465),
    .X(_01016_));
 sg13g2_mux2_1 _22143_ (.A0(net1094),
    .A1(_10118_),
    .S(net516),
    .X(_04741_));
 sg13g2_mux2_1 _22144_ (.A0(_04741_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net465),
    .X(_01017_));
 sg13g2_buf_1 _22145_ (.A(_04729_),
    .X(_04742_));
 sg13g2_nor2_1 _22146_ (.A(_08822_),
    .B(net515),
    .Y(_04743_));
 sg13g2_a21oi_1 _22147_ (.A1(_10527_),
    .A2(net516),
    .Y(_04744_),
    .B1(_04743_));
 sg13g2_nand2_1 _22148_ (.Y(_04745_),
    .A(\cpu.ex.r_stmp[12] ),
    .B(net466));
 sg13g2_o21ai_1 _22149_ (.B1(_04745_),
    .Y(_01018_),
    .A1(net465),
    .A2(_04744_));
 sg13g2_mux2_1 _22150_ (.A0(net611),
    .A1(_10579_),
    .S(net516),
    .X(_04746_));
 sg13g2_mux2_1 _22151_ (.A0(_04746_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net465),
    .X(_01019_));
 sg13g2_mux2_1 _22152_ (.A0(net672),
    .A1(_10554_),
    .S(net515),
    .X(_04747_));
 sg13g2_mux2_1 _22153_ (.A0(_04747_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(_04740_),
    .X(_01020_));
 sg13g2_mux2_1 _22154_ (.A0(net890),
    .A1(_10602_),
    .S(net515),
    .X(_04748_));
 sg13g2_mux2_1 _22155_ (.A0(_04748_),
    .A1(\cpu.ex.r_stmp[15] ),
    .S(net466),
    .X(_01021_));
 sg13g2_nor2_1 _22156_ (.A(_09975_),
    .B(net515),
    .Y(_04749_));
 sg13g2_a21oi_1 _22157_ (.A1(_10318_),
    .A2(net516),
    .Y(_04750_),
    .B1(_04749_));
 sg13g2_nand2_1 _22158_ (.Y(_04751_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net466));
 sg13g2_o21ai_1 _22159_ (.B1(_04751_),
    .Y(_01022_),
    .A1(net465),
    .A2(_04750_));
 sg13g2_nor2_1 _22160_ (.A(net638),
    .B(net515),
    .Y(_04752_));
 sg13g2_a21oi_1 _22161_ (.A1(_10386_),
    .A2(net516),
    .Y(_04753_),
    .B1(_04752_));
 sg13g2_nand2_1 _22162_ (.Y(_04754_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net466));
 sg13g2_o21ai_1 _22163_ (.B1(_04754_),
    .Y(_01023_),
    .A1(net465),
    .A2(_04753_));
 sg13g2_nor2_1 _22164_ (.A(_09131_),
    .B(_04742_),
    .Y(_04755_));
 sg13g2_a21oi_1 _22165_ (.A1(_10246_),
    .A2(net516),
    .Y(_04756_),
    .B1(_04755_));
 sg13g2_nand2_1 _22166_ (.Y(_04757_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(_04737_));
 sg13g2_o21ai_1 _22167_ (.B1(_04757_),
    .Y(_01024_),
    .A1(net465),
    .A2(_04756_));
 sg13g2_nor2_1 _22168_ (.A(net712),
    .B(_04729_),
    .Y(_04758_));
 sg13g2_a21oi_1 _22169_ (.A1(_10462_),
    .A2(_04730_),
    .Y(_04759_),
    .B1(_04758_));
 sg13g2_nand2_1 _22170_ (.Y(_04760_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_04736_));
 sg13g2_o21ai_1 _22171_ (.B1(_04760_),
    .Y(_01025_),
    .A1(_04740_),
    .A2(_04759_));
 sg13g2_nor2_1 _22172_ (.A(net865),
    .B(_04729_),
    .Y(_04761_));
 sg13g2_a21oi_1 _22173_ (.A1(_10448_),
    .A2(net516),
    .Y(_04762_),
    .B1(_04761_));
 sg13g2_nand2_1 _22174_ (.Y(_04763_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_04736_));
 sg13g2_o21ai_1 _22175_ (.B1(_04763_),
    .Y(_01026_),
    .A1(net465),
    .A2(_04762_));
 sg13g2_mux2_1 _22176_ (.A0(net953),
    .A1(_10511_),
    .S(_04742_),
    .X(_04764_));
 sg13g2_mux2_1 _22177_ (.A0(_04764_),
    .A1(\cpu.ex.r_stmp[6] ),
    .S(_04737_),
    .X(_01027_));
 sg13g2_mux2_1 _22178_ (.A0(net1037),
    .A1(_10406_),
    .S(net515),
    .X(_04765_));
 sg13g2_mux2_1 _22179_ (.A0(_04765_),
    .A1(\cpu.ex.r_stmp[7] ),
    .S(net466),
    .X(_01028_));
 sg13g2_mux2_1 _22180_ (.A0(net1038),
    .A1(_10697_),
    .S(net515),
    .X(_04766_));
 sg13g2_mux2_1 _22181_ (.A0(_04766_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net466),
    .X(_01029_));
 sg13g2_mux2_1 _22182_ (.A0(_10627_),
    .A1(_10629_),
    .S(net515),
    .X(_04767_));
 sg13g2_mux2_1 _22183_ (.A0(_04767_),
    .A1(\cpu.ex.r_stmp[9] ),
    .S(net466),
    .X(_01030_));
 sg13g2_a21o_1 _22184_ (.A2(net374),
    .A1(_10050_),
    .B1(net233),
    .X(_04768_));
 sg13g2_nor2_1 _22185_ (.A(_11336_),
    .B(_04768_),
    .Y(_04769_));
 sg13g2_nor2_1 _22186_ (.A(net113),
    .B(_04152_),
    .Y(_04770_));
 sg13g2_o21ai_1 _22187_ (.B1(_03500_),
    .Y(_04771_),
    .A1(_11389_),
    .A2(net137));
 sg13g2_or2_1 _22188_ (.X(_04772_),
    .B(_04771_),
    .A(_04234_));
 sg13g2_nor2_1 _22189_ (.A(_03483_),
    .B(_04074_),
    .Y(_04773_));
 sg13g2_a221oi_1 _22190_ (.B2(_04028_),
    .C1(_04773_),
    .B1(net118),
    .A1(net140),
    .Y(_04774_),
    .A2(net130));
 sg13g2_o21ai_1 _22191_ (.B1(_04248_),
    .Y(_04775_),
    .A1(_03549_),
    .A2(_04307_));
 sg13g2_a221oi_1 _22192_ (.B2(net159),
    .C1(_04775_),
    .B1(_04055_),
    .A1(net136),
    .Y(_04776_),
    .A2(_04059_));
 sg13g2_nand3_1 _22193_ (.B(_04774_),
    .C(_04776_),
    .A(_04772_),
    .Y(_04777_));
 sg13g2_o21ai_1 _22194_ (.B1(_04521_),
    .Y(_04778_),
    .A1(net198),
    .A2(_04169_));
 sg13g2_nand2_1 _22195_ (.Y(_04779_),
    .A(_04337_),
    .B(_04593_));
 sg13g2_or4_1 _22196_ (.A(_04642_),
    .B(_04777_),
    .C(_04778_),
    .D(_04779_),
    .X(_04780_));
 sg13g2_a21oi_1 _22197_ (.A1(_11319_),
    .A2(net142),
    .Y(_04781_),
    .B1(_04780_));
 sg13g2_a21oi_1 _22198_ (.A1(_09714_),
    .A2(_04780_),
    .Y(_04782_),
    .B1(net1055));
 sg13g2_nor3_1 _22199_ (.A(_04770_),
    .B(_04781_),
    .C(_04782_),
    .Y(_04783_));
 sg13g2_or3_1 _22200_ (.A(net1041),
    .B(net1039),
    .C(_04447_),
    .X(_04784_));
 sg13g2_or2_1 _22201_ (.X(_04785_),
    .B(_04117_),
    .A(net1021));
 sg13g2_o21ai_1 _22202_ (.B1(_04785_),
    .Y(_04786_),
    .A1(net176),
    .A2(_04784_));
 sg13g2_o21ai_1 _22203_ (.B1(net176),
    .Y(_04787_),
    .A1(net1022),
    .A2(_04784_));
 sg13g2_a22oi_1 _22204_ (.Y(_04788_),
    .B1(_04787_),
    .B2(_11316_),
    .A2(_04786_),
    .A1(_04193_));
 sg13g2_and2_1 _22205_ (.A(net1040),
    .B(net183),
    .X(_04789_));
 sg13g2_nor4_2 _22206_ (.A(net234),
    .B(_04783_),
    .C(_04788_),
    .Y(_04790_),
    .D(_04789_));
 sg13g2_a21oi_1 _22207_ (.A1(_11345_),
    .A2(_11346_),
    .Y(_04791_),
    .B1(_09097_));
 sg13g2_buf_1 _22208_ (.A(_04791_),
    .X(_04792_));
 sg13g2_nand2_1 _22209_ (.Y(_04793_),
    .A(_04125_),
    .B(_11357_));
 sg13g2_nor2_1 _22210_ (.A(net711),
    .B(_04793_),
    .Y(_04794_));
 sg13g2_nand2b_1 _22211_ (.Y(_04795_),
    .B(_04794_),
    .A_N(_04790_));
 sg13g2_buf_1 _22212_ (.A(_11360_),
    .X(_04796_));
 sg13g2_buf_1 _22213_ (.A(_03446_),
    .X(_04797_));
 sg13g2_buf_1 _22214_ (.A(_11790_),
    .X(_04798_));
 sg13g2_buf_1 _22215_ (.A(net546),
    .X(_04799_));
 sg13g2_a22oi_1 _22216_ (.Y(_04800_),
    .B1(net464),
    .B2(\cpu.dcache.r_data[3][0] ),
    .A2(net416),
    .A1(\cpu.dcache.r_data[1][0] ));
 sg13g2_a22oi_1 _22217_ (.Y(_04801_),
    .B1(net532),
    .B2(\cpu.dcache.r_data[6][0] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][0] ));
 sg13g2_buf_1 _22218_ (.A(_09092_),
    .X(_04802_));
 sg13g2_mux2_1 _22219_ (.A0(\cpu.dcache.r_data[5][0] ),
    .A1(\cpu.dcache.r_data[7][0] ),
    .S(net514),
    .X(_04803_));
 sg13g2_a22oi_1 _22220_ (.Y(_04804_),
    .B1(_04803_),
    .B2(net682),
    .A2(net673),
    .A1(\cpu.dcache.r_data[4][0] ));
 sg13g2_nand2b_1 _22221_ (.Y(_04805_),
    .B(net670),
    .A_N(_04804_));
 sg13g2_nand3_1 _22222_ (.B(_04801_),
    .C(_04805_),
    .A(_04800_),
    .Y(_04806_));
 sg13g2_buf_1 _22223_ (.A(net494),
    .X(_04807_));
 sg13g2_buf_1 _22224_ (.A(net403),
    .X(_04808_));
 sg13g2_mux2_1 _22225_ (.A0(\cpu.dcache.r_data[0][0] ),
    .A1(_04806_),
    .S(net365),
    .X(_04809_));
 sg13g2_a22oi_1 _22226_ (.Y(_04810_),
    .B1(net476),
    .B2(\cpu.dcache.r_data[5][16] ),
    .A2(net416),
    .A1(\cpu.dcache.r_data[1][16] ));
 sg13g2_a22oi_1 _22227_ (.Y(_04811_),
    .B1(net464),
    .B2(\cpu.dcache.r_data[3][16] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][16] ));
 sg13g2_mux2_1 _22228_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(\cpu.dcache.r_data[6][16] ),
    .S(net619),
    .X(_04812_));
 sg13g2_a22oi_1 _22229_ (.Y(_04813_),
    .B1(_04812_),
    .B2(net713),
    .A2(net669),
    .A1(\cpu.dcache.r_data[7][16] ));
 sg13g2_nand2b_1 _22230_ (.Y(_04814_),
    .B(net670),
    .A_N(_04813_));
 sg13g2_nand4_1 _22231_ (.B(_04810_),
    .C(_04811_),
    .A(net403),
    .Y(_04815_),
    .D(_04814_));
 sg13g2_o21ai_1 _22232_ (.B1(_04815_),
    .Y(_04816_),
    .A1(\cpu.dcache.r_data[0][16] ),
    .A2(net365));
 sg13g2_or2_1 _22233_ (.X(_04817_),
    .B(_04816_),
    .A(net885));
 sg13g2_nor2_1 _22234_ (.A(_11790_),
    .B(_04817_),
    .Y(_04818_));
 sg13g2_a21oi_1 _22235_ (.A1(net945),
    .A2(_04809_),
    .Y(_04819_),
    .B1(_04818_));
 sg13g2_nand3b_1 _22236_ (.B(net1111),
    .C(_09656_),
    .Y(_04820_),
    .A_N(_08772_));
 sg13g2_buf_1 _22237_ (.A(_04820_),
    .X(_04821_));
 sg13g2_buf_1 _22238_ (.A(net636),
    .X(_04822_));
 sg13g2_buf_1 _22239_ (.A(net550),
    .X(_04823_));
 sg13g2_buf_1 _22240_ (.A(net416),
    .X(_04824_));
 sg13g2_a22oi_1 _22241_ (.Y(_04825_),
    .B1(net476),
    .B2(\cpu.dcache.r_data[5][8] ),
    .A2(net364),
    .A1(\cpu.dcache.r_data[1][8] ));
 sg13g2_a22oi_1 _22242_ (.Y(_04826_),
    .B1(net464),
    .B2(\cpu.dcache.r_data[3][8] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][8] ));
 sg13g2_mux2_1 _22243_ (.A0(\cpu.dcache.r_data[4][8] ),
    .A1(\cpu.dcache.r_data[6][8] ),
    .S(net514),
    .X(_04827_));
 sg13g2_a22oi_1 _22244_ (.Y(_04828_),
    .B1(_04827_),
    .B2(_03698_),
    .A2(net669),
    .A1(\cpu.dcache.r_data[7][8] ));
 sg13g2_nand2b_1 _22245_ (.Y(_04829_),
    .B(net603),
    .A_N(_04828_));
 sg13g2_and4_1 _22246_ (.A(net365),
    .B(_04825_),
    .C(_04826_),
    .D(_04829_),
    .X(_04830_));
 sg13g2_a21oi_1 _22247_ (.A1(_00312_),
    .A2(net463),
    .Y(_04831_),
    .B1(_04830_));
 sg13g2_nand2_1 _22248_ (.Y(_04832_),
    .A(\cpu.dcache.r_data[3][24] ),
    .B(net464));
 sg13g2_a22oi_1 _22249_ (.Y(_04833_),
    .B1(_09394_),
    .B2(\cpu.dcache.r_data[4][24] ),
    .A2(net548),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_a22oi_1 _22250_ (.Y(_04834_),
    .B1(_02905_),
    .B2(\cpu.dcache.r_data[7][24] ),
    .A2(_09286_),
    .A1(\cpu.dcache.r_data[6][24] ));
 sg13g2_a22oi_1 _22251_ (.Y(_04835_),
    .B1(_09346_),
    .B2(\cpu.dcache.r_data[5][24] ),
    .A2(_02887_),
    .A1(\cpu.dcache.r_data[1][24] ));
 sg13g2_nand4_1 _22252_ (.B(_04833_),
    .C(_04834_),
    .A(_04832_),
    .Y(_04836_),
    .D(_04835_));
 sg13g2_nor2_1 _22253_ (.A(net550),
    .B(_04836_),
    .Y(_04837_));
 sg13g2_a21oi_1 _22254_ (.A1(_00311_),
    .A2(_04823_),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_a221oi_1 _22255_ (.B2(net991),
    .C1(net636),
    .B1(_04838_),
    .A1(net759),
    .Y(_04839_),
    .A2(_04831_));
 sg13g2_a21oi_1 _22256_ (.A1(_04819_),
    .A2(net581),
    .Y(_04840_),
    .B1(_04839_));
 sg13g2_nor2_1 _22257_ (.A(_08771_),
    .B(net636),
    .Y(_04841_));
 sg13g2_buf_1 _22258_ (.A(_04841_),
    .X(_04842_));
 sg13g2_nand2_1 _22259_ (.Y(_04843_),
    .A(net759),
    .B(_04809_));
 sg13g2_nand3_1 _22260_ (.B(net513),
    .C(_04843_),
    .A(_04817_),
    .Y(_04844_));
 sg13g2_o21ai_1 _22261_ (.B1(_04844_),
    .Y(_04845_),
    .A1(_04840_),
    .A2(net513));
 sg13g2_and2_1 _22262_ (.A(net953),
    .B(_09819_),
    .X(_04846_));
 sg13g2_buf_1 _22263_ (.A(_04846_),
    .X(_04847_));
 sg13g2_mux2_1 _22264_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(\cpu.intr.r_timer_reload[16] ),
    .S(net730),
    .X(_04848_));
 sg13g2_and2_1 _22265_ (.A(net898),
    .B(\cpu.intr.r_clock_cmp[16] ),
    .X(_04849_));
 sg13g2_a21oi_1 _22266_ (.A1(net759),
    .A2(\cpu.intr.r_clock_cmp[0] ),
    .Y(_04850_),
    .B1(_04849_));
 sg13g2_nor2_1 _22267_ (.A(net772),
    .B(net681),
    .Y(_04851_));
 sg13g2_nor2b_1 _22268_ (.A(net666),
    .B_N(_04851_),
    .Y(_04852_));
 sg13g2_buf_1 _22269_ (.A(_04852_),
    .X(_04853_));
 sg13g2_buf_1 _22270_ (.A(_04853_),
    .X(_04854_));
 sg13g2_o21ai_1 _22271_ (.B1(net402),
    .Y(_04855_),
    .A1(_09033_),
    .A2(_09034_));
 sg13g2_o21ai_1 _22272_ (.B1(_04855_),
    .Y(_04856_),
    .A1(net597),
    .A2(_04850_));
 sg13g2_a21oi_1 _22273_ (.A1(net474),
    .A2(_04848_),
    .Y(_04857_),
    .B1(_04856_));
 sg13g2_nor2_1 _22274_ (.A(net1036),
    .B(_09947_),
    .Y(_04858_));
 sg13g2_buf_2 _22275_ (.A(_04858_),
    .X(_04859_));
 sg13g2_buf_1 _22276_ (.A(_04859_),
    .X(_04860_));
 sg13g2_nand2_1 _22277_ (.Y(_04861_),
    .A(_09967_),
    .B(net462));
 sg13g2_buf_1 _22278_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04862_));
 sg13g2_nand2_1 _22279_ (.Y(_04863_),
    .A(net782),
    .B(_09841_));
 sg13g2_o21ai_1 _22280_ (.B1(_04863_),
    .Y(_04864_),
    .A1(net730),
    .A2(_00285_));
 sg13g2_a22oi_1 _22281_ (.Y(_04865_),
    .B1(_04864_),
    .B2(net475),
    .A2(net429),
    .A1(_04862_));
 sg13g2_nand2_1 _22282_ (.Y(_04866_),
    .A(_09811_),
    .B(net784));
 sg13g2_buf_1 _22283_ (.A(_04866_),
    .X(_04867_));
 sg13g2_nor3_1 _22284_ (.A(net772),
    .B(net619),
    .C(_04867_),
    .Y(_04868_));
 sg13g2_buf_2 _22285_ (.A(_04868_),
    .X(_04869_));
 sg13g2_buf_1 _22286_ (.A(_04869_),
    .X(_04870_));
 sg13g2_and2_1 _22287_ (.A(net666),
    .B(_04867_),
    .X(_04871_));
 sg13g2_buf_1 _22288_ (.A(_04871_),
    .X(_04872_));
 sg13g2_nor2_1 _22289_ (.A(_04802_),
    .B(_04872_),
    .Y(_04873_));
 sg13g2_nor2_1 _22290_ (.A(net670),
    .B(_04873_),
    .Y(_04874_));
 sg13g2_buf_1 _22291_ (.A(_04874_),
    .X(_04875_));
 sg13g2_o21ai_1 _22292_ (.B1(net333),
    .Y(_04876_),
    .A1(_09033_),
    .A2(_09034_));
 sg13g2_nand2b_1 _22293_ (.Y(_04877_),
    .B(_04876_),
    .A_N(net401));
 sg13g2_nand2_1 _22294_ (.Y(_04878_),
    .A(\cpu.intr.r_enable[0] ),
    .B(_04877_));
 sg13g2_nand4_1 _22295_ (.B(_04861_),
    .C(_04865_),
    .A(_04857_),
    .Y(_04879_),
    .D(_04878_));
 sg13g2_nand2b_1 _22296_ (.Y(_04880_),
    .B(_09821_),
    .A_N(_09016_));
 sg13g2_buf_1 _22297_ (.A(_04880_),
    .X(_04881_));
 sg13g2_o21ai_1 _22298_ (.B1(net712),
    .Y(_04882_),
    .A1(net894),
    .A2(net773));
 sg13g2_buf_2 _22299_ (.A(_04882_),
    .X(_04883_));
 sg13g2_nand2_1 _22300_ (.Y(_04884_),
    .A(net1106),
    .B(net784));
 sg13g2_buf_2 _22301_ (.A(_04884_),
    .X(_04885_));
 sg13g2_nor3_1 _22302_ (.A(net772),
    .B(net681),
    .C(_04885_),
    .Y(_04886_));
 sg13g2_buf_1 _22303_ (.A(_04886_),
    .X(_04887_));
 sg13g2_nand2_1 _22304_ (.Y(_04888_),
    .A(net891),
    .B(net681));
 sg13g2_buf_2 _22305_ (.A(_04888_),
    .X(_04889_));
 sg13g2_nor3_1 _22306_ (.A(net1106),
    .B(net682),
    .C(_04889_),
    .Y(_04890_));
 sg13g2_buf_1 _22307_ (.A(_04890_),
    .X(_04891_));
 sg13g2_a22oi_1 _22308_ (.Y(_04892_),
    .B1(net400),
    .B2(\cpu.uart.r_div_value[0] ),
    .A2(net461),
    .A1(\cpu.uart.r_x_invert ));
 sg13g2_nor2_1 _22309_ (.A(net666),
    .B(_04889_),
    .Y(_04893_));
 sg13g2_buf_1 _22310_ (.A(_04893_),
    .X(_04894_));
 sg13g2_a22oi_1 _22311_ (.Y(_04895_),
    .B1(net399),
    .B2(\cpu.uart.r_div_value[8] ),
    .A2(_04869_),
    .A1(_09033_));
 sg13g2_nand2_1 _22312_ (.Y(_04896_),
    .A(_04892_),
    .B(_04895_));
 sg13g2_a21oi_1 _22313_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04883_),
    .Y(_04897_),
    .B1(_04896_));
 sg13g2_o21ai_1 _22314_ (.B1(net1031),
    .Y(_04898_),
    .A1(net512),
    .A2(_04897_));
 sg13g2_a21oi_1 _22315_ (.A1(_04847_),
    .A2(_04879_),
    .Y(_04899_),
    .B1(_04898_));
 sg13g2_nor2b_1 _22316_ (.A(_09010_),
    .B_N(_09016_),
    .Y(_04900_));
 sg13g2_buf_2 _22317_ (.A(_04900_),
    .X(_04901_));
 sg13g2_o21ai_1 _22318_ (.B1(_09253_),
    .Y(_04902_),
    .A1(net892),
    .A2(_09389_));
 sg13g2_nand2_1 _22319_ (.Y(_04903_),
    .A(net682),
    .B(_09389_));
 sg13g2_a22oi_1 _22320_ (.Y(_04904_),
    .B1(_04903_),
    .B2(net619),
    .A2(net773),
    .A1(_09811_));
 sg13g2_nor2_1 _22321_ (.A(_11724_),
    .B(_04904_),
    .Y(_04905_));
 sg13g2_a21oi_1 _22322_ (.A1(_11724_),
    .A2(_04902_),
    .Y(_04906_),
    .B1(_04905_));
 sg13g2_inv_1 _22323_ (.Y(_04907_),
    .A(_09389_));
 sg13g2_nor2_1 _22324_ (.A(net514),
    .B(_04907_),
    .Y(_04908_));
 sg13g2_nand2_1 _22325_ (.Y(_04909_),
    .A(net885),
    .B(net712));
 sg13g2_nor2_1 _22326_ (.A(net995),
    .B(net1036),
    .Y(_04910_));
 sg13g2_a22oi_1 _22327_ (.Y(_04911_),
    .B1(_04910_),
    .B2(net894),
    .A2(_04909_),
    .A1(_04908_));
 sg13g2_o21ai_1 _22328_ (.B1(_04911_),
    .Y(_04912_),
    .A1(net670),
    .A2(_04906_));
 sg13g2_buf_1 _22329_ (.A(_04912_),
    .X(_04913_));
 sg13g2_inv_1 _22330_ (.Y(_04914_),
    .A(_04913_));
 sg13g2_nand3_1 _22331_ (.B(_09051_),
    .C(_04914_),
    .A(_09050_),
    .Y(_04915_));
 sg13g2_buf_2 _22332_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04916_));
 sg13g2_nor3_1 _22333_ (.A(_09818_),
    .B(net1106),
    .C(_12544_),
    .Y(_04917_));
 sg13g2_buf_1 _22334_ (.A(_04917_),
    .X(_04918_));
 sg13g2_buf_2 _22335_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04919_));
 sg13g2_nor3_1 _22336_ (.A(_09389_),
    .B(_04867_),
    .C(_04889_),
    .Y(_04920_));
 sg13g2_buf_1 _22337_ (.A(_04920_),
    .X(_04921_));
 sg13g2_and2_1 _22338_ (.A(_10431_),
    .B(net400),
    .X(_04922_));
 sg13g2_buf_2 _22339_ (.A(_04922_),
    .X(_04923_));
 sg13g2_a22oi_1 _22340_ (.Y(_04924_),
    .B1(_04923_),
    .B2(_09050_),
    .A2(net398),
    .A1(_04919_));
 sg13g2_buf_2 _22341_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04925_));
 sg13g2_buf_1 _22342_ (.A(_09389_),
    .X(_04926_));
 sg13g2_nor3_1 _22343_ (.A(net944),
    .B(_04885_),
    .C(_04889_),
    .Y(_04927_));
 sg13g2_buf_1 _22344_ (.A(_04927_),
    .X(_04928_));
 sg13g2_and2_1 _22345_ (.A(_10431_),
    .B(_04869_),
    .X(_04929_));
 sg13g2_buf_2 _22346_ (.A(_04929_),
    .X(_04930_));
 sg13g2_a22oi_1 _22347_ (.Y(_04931_),
    .B1(_04930_),
    .B2(_09051_),
    .A2(net397),
    .A1(_04925_));
 sg13g2_buf_1 _22348_ (.A(net944),
    .X(_04932_));
 sg13g2_buf_2 _22349_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04933_));
 sg13g2_nor2_1 _22350_ (.A(net885),
    .B(net597),
    .Y(_04934_));
 sg13g2_buf_2 _22351_ (.A(_04934_),
    .X(_04935_));
 sg13g2_nand3_1 _22352_ (.B(_04933_),
    .C(_04935_),
    .A(net837),
    .Y(_04936_));
 sg13g2_buf_2 _22353_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04937_));
 sg13g2_nand2_1 _22354_ (.Y(_04938_),
    .A(net995),
    .B(_04887_));
 sg13g2_buf_2 _22355_ (.A(_04938_),
    .X(_04939_));
 sg13g2_inv_1 _22356_ (.Y(_04940_),
    .A(_04939_));
 sg13g2_and2_1 _22357_ (.A(_04907_),
    .B(_04869_),
    .X(_04941_));
 sg13g2_buf_1 _22358_ (.A(_04941_),
    .X(_04942_));
 sg13g2_buf_2 _22359_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04943_));
 sg13g2_a22oi_1 _22360_ (.Y(_04944_),
    .B1(_04942_),
    .B2(_04943_),
    .A2(_04940_),
    .A1(_04937_));
 sg13g2_nand4_1 _22361_ (.B(_04931_),
    .C(_04936_),
    .A(_04924_),
    .Y(_04945_),
    .D(_04944_));
 sg13g2_a21oi_1 _22362_ (.A1(_04916_),
    .A2(_04918_),
    .Y(_04946_),
    .B1(_04945_));
 sg13g2_nand2_1 _22363_ (.Y(_04947_),
    .A(_04915_),
    .B(_04946_));
 sg13g2_buf_1 _22364_ (.A(net400),
    .X(_04948_));
 sg13g2_nor2_1 _22365_ (.A(net898),
    .B(net533),
    .Y(_04949_));
 sg13g2_buf_1 _22366_ (.A(_04949_),
    .X(_04950_));
 sg13g2_buf_1 _22367_ (.A(_04950_),
    .X(_04951_));
 sg13g2_nor3_1 _22368_ (.A(_00314_),
    .B(net666),
    .C(_04889_),
    .Y(_04952_));
 sg13g2_a221oi_1 _22369_ (.B2(\cpu.spi.r_mode[1][0] ),
    .C1(_04952_),
    .B1(net362),
    .A1(_11743_),
    .Y(_04953_),
    .A2(net363));
 sg13g2_o21ai_1 _22370_ (.B1(net619),
    .Y(_04954_),
    .A1(net712),
    .A2(_09389_));
 sg13g2_inv_1 _22371_ (.Y(_04955_),
    .A(_00228_));
 sg13g2_nor2_1 _22372_ (.A(net784),
    .B(net772),
    .Y(_04956_));
 sg13g2_a22oi_1 _22373_ (.Y(_04957_),
    .B1(_04956_),
    .B2(_09389_),
    .A2(_04955_),
    .A1(_09130_));
 sg13g2_nor3_1 _22374_ (.A(net1106),
    .B(net765),
    .C(_09283_),
    .Y(_04958_));
 sg13g2_a21oi_1 _22375_ (.A1(net1106),
    .A2(_04957_),
    .Y(_04959_),
    .B1(_04958_));
 sg13g2_a21oi_1 _22376_ (.A1(net892),
    .A2(_04954_),
    .Y(_04960_),
    .B1(_04959_));
 sg13g2_nor3_2 _22377_ (.A(_09818_),
    .B(net666),
    .C(_04889_),
    .Y(_04961_));
 sg13g2_nor3_1 _22378_ (.A(_04918_),
    .B(_04960_),
    .C(_04961_),
    .Y(_04962_));
 sg13g2_buf_2 _22379_ (.A(_04962_),
    .X(_04963_));
 sg13g2_a22oi_1 _22380_ (.Y(_04964_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net496),
    .A2(_00228_),
    .A1(_09038_));
 sg13g2_nand3_1 _22381_ (.B(net780),
    .C(\cpu.spi.r_ready ),
    .A(net759),
    .Y(_04965_));
 sg13g2_o21ai_1 _22382_ (.B1(_04965_),
    .Y(_04966_),
    .A1(net759),
    .A2(_04964_));
 sg13g2_nand3_1 _22383_ (.B(net944),
    .C(net612),
    .A(_09080_),
    .Y(_04967_));
 sg13g2_buf_2 _22384_ (.A(_04967_),
    .X(_04968_));
 sg13g2_buf_1 _22385_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04969_));
 sg13g2_nor3_1 _22386_ (.A(net944),
    .B(net666),
    .C(_04889_),
    .Y(_04970_));
 sg13g2_buf_2 _22387_ (.A(_04970_),
    .X(_04971_));
 sg13g2_and2_1 _22388_ (.A(net995),
    .B(\cpu.spi.r_mode[2][0] ),
    .X(_04972_));
 sg13g2_a22oi_1 _22389_ (.Y(_04973_),
    .B1(_04972_),
    .B2(net400),
    .A2(_04971_),
    .A1(_04969_));
 sg13g2_o21ai_1 _22390_ (.B1(_04973_),
    .Y(_04974_),
    .A1(_00313_),
    .A2(_04968_));
 sg13g2_a221oi_1 _22391_ (.B2(net551),
    .C1(_04974_),
    .B1(_04966_),
    .A1(_09163_),
    .Y(_04975_),
    .A2(_04963_));
 sg13g2_o21ai_1 _22392_ (.B1(_04975_),
    .Y(_04976_),
    .A1(net864),
    .A2(_04953_));
 sg13g2_and2_1 _22393_ (.A(_09010_),
    .B(_09016_),
    .X(_04977_));
 sg13g2_buf_2 _22394_ (.A(_04977_),
    .X(_04978_));
 sg13g2_a22oi_1 _22395_ (.Y(_04979_),
    .B1(_04976_),
    .B2(_04978_),
    .A2(_04947_),
    .A1(_04901_));
 sg13g2_a22oi_1 _22396_ (.Y(_04980_),
    .B1(_04899_),
    .B2(_04979_),
    .A2(_04845_),
    .A1(net886));
 sg13g2_nand2_1 _22397_ (.Y(_04981_),
    .A(_03446_),
    .B(_04980_));
 sg13g2_o21ai_1 _22398_ (.B1(_04981_),
    .Y(_04982_),
    .A1(_03747_),
    .A2(net32));
 sg13g2_buf_1 _22399_ (.A(_11360_),
    .X(_04983_));
 sg13g2_buf_1 _22400_ (.A(_04791_),
    .X(_04984_));
 sg13g2_o21ai_1 _22401_ (.B1(net719),
    .Y(_04985_),
    .A1(_10183_),
    .A2(net710));
 sg13g2_nor2_1 _22402_ (.A(net153),
    .B(_04985_),
    .Y(_04986_));
 sg13g2_a21oi_1 _22403_ (.A1(_04796_),
    .A2(_04982_),
    .Y(_04987_),
    .B1(_04986_));
 sg13g2_o21ai_1 _22404_ (.B1(_04987_),
    .Y(_01031_),
    .A1(_04769_),
    .A2(_04795_));
 sg13g2_buf_1 _22405_ (.A(_10183_),
    .X(_04988_));
 sg13g2_nor2_1 _22406_ (.A(net232),
    .B(_11360_),
    .Y(_04989_));
 sg13g2_nand2b_1 _22407_ (.Y(_04990_),
    .B(net711),
    .A_N(_04722_));
 sg13g2_o21ai_1 _22408_ (.B1(_04990_),
    .Y(_04991_),
    .A1(_04792_),
    .A2(_04718_));
 sg13g2_buf_1 _22409_ (.A(_03446_),
    .X(_04992_));
 sg13g2_nor2_1 _22410_ (.A(_09064_),
    .B(_04913_),
    .Y(_04993_));
 sg13g2_nor2b_1 _22411_ (.A(_00160_),
    .B_N(_04869_),
    .Y(_04994_));
 sg13g2_a22oi_1 _22412_ (.Y(_04995_),
    .B1(net461),
    .B2(_09048_),
    .A2(_09961_),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_a221oi_1 _22413_ (.B2(net10),
    .C1(net1036),
    .B1(net545),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .Y(_04996_),
    .A2(_09394_));
 sg13g2_o21ai_1 _22414_ (.B1(_09080_),
    .Y(_04997_),
    .A1(_00162_),
    .A2(net597));
 sg13g2_nand2b_1 _22415_ (.Y(_04998_),
    .B(_04997_),
    .A_N(_04996_));
 sg13g2_nand3_1 _22416_ (.B(_04995_),
    .C(_04998_),
    .A(net944),
    .Y(_04999_));
 sg13g2_o21ai_1 _22417_ (.B1(_04999_),
    .Y(_05000_),
    .A1(net944),
    .A2(_04994_));
 sg13g2_and3_1 _22418_ (.X(_05001_),
    .A(_09048_),
    .B(net944),
    .C(_04853_));
 sg13g2_o21ai_1 _22419_ (.B1(\cpu.gpio.r_enable_io[7] ),
    .Y(_05002_),
    .A1(_04961_),
    .A2(_05001_));
 sg13g2_buf_1 _22420_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05003_));
 sg13g2_nand3b_1 _22421_ (.B(_04853_),
    .C(net995),
    .Y(_05004_),
    .A_N(_00161_));
 sg13g2_o21ai_1 _22422_ (.B1(_05004_),
    .Y(_05005_),
    .A1(_00159_),
    .A2(_04939_));
 sg13g2_a221oi_1 _22423_ (.B2(_09063_),
    .C1(_05005_),
    .B1(_04930_),
    .A1(_05003_),
    .Y(_05006_),
    .A2(_04921_));
 sg13g2_inv_1 _22424_ (.Y(_05007_),
    .A(_00158_));
 sg13g2_a22oi_1 _22425_ (.Y(_05008_),
    .B1(net397),
    .B2(_05007_),
    .A2(_04923_),
    .A1(\cpu.gpio.r_enable_in[7] ));
 sg13g2_nand4_1 _22426_ (.B(_05002_),
    .C(_05006_),
    .A(_05000_),
    .Y(_05009_),
    .D(_05008_));
 sg13g2_o21ai_1 _22427_ (.B1(_04901_),
    .Y(_05010_),
    .A1(_04993_),
    .A2(_05009_));
 sg13g2_nor2b_1 _22428_ (.A(_00222_),
    .B_N(_04963_),
    .Y(_05011_));
 sg13g2_buf_1 _22429_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05012_));
 sg13g2_nor2_1 _22430_ (.A(_09130_),
    .B(_04885_),
    .Y(_05013_));
 sg13g2_buf_2 _22431_ (.A(_05013_),
    .X(_05014_));
 sg13g2_nand2_1 _22432_ (.Y(_05015_),
    .A(_10431_),
    .B(net399));
 sg13g2_buf_1 _22433_ (.A(_05015_),
    .X(_05016_));
 sg13g2_nor2_1 _22434_ (.A(_00157_),
    .B(_05016_),
    .Y(_05017_));
 sg13g2_a221oi_1 _22435_ (.B2(\cpu.spi.r_timeout[7] ),
    .C1(_05017_),
    .B1(_05014_),
    .A1(_05012_),
    .Y(_05018_),
    .A2(_04971_));
 sg13g2_o21ai_1 _22436_ (.B1(_05018_),
    .Y(_05019_),
    .A1(_00156_),
    .A2(_04968_));
 sg13g2_o21ai_1 _22437_ (.B1(_04978_),
    .Y(_05020_),
    .A1(_05011_),
    .A2(_05019_));
 sg13g2_nor2_1 _22438_ (.A(_09821_),
    .B(net333),
    .Y(_05021_));
 sg13g2_a22oi_1 _22439_ (.Y(_05022_),
    .B1(net476),
    .B2(\cpu.intr.r_clock_cmp[7] ),
    .A2(net598),
    .A1(_09996_));
 sg13g2_and2_1 _22440_ (.A(net1036),
    .B(_09849_),
    .X(_05023_));
 sg13g2_a21oi_1 _22441_ (.A1(net885),
    .A2(_09825_),
    .Y(_05024_),
    .B1(_05023_));
 sg13g2_buf_2 _22442_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05025_));
 sg13g2_mux2_1 _22443_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(\cpu.intr.r_timer_reload[23] ),
    .S(net1106),
    .X(_05026_));
 sg13g2_a22oi_1 _22444_ (.Y(_05027_),
    .B1(_05026_),
    .B2(net531),
    .A2(_09961_),
    .A1(_05025_));
 sg13g2_o21ai_1 _22445_ (.B1(_05027_),
    .Y(_05028_),
    .A1(net533),
    .A2(_05024_));
 sg13g2_a21oi_1 _22446_ (.A1(\cpu.intr.r_clock_cmp[23] ),
    .A2(_04935_),
    .Y(_05029_),
    .B1(_05028_));
 sg13g2_o21ai_1 _22447_ (.B1(_05029_),
    .Y(_05030_),
    .A1(net898),
    .A2(_05022_));
 sg13g2_a22oi_1 _22448_ (.Y(_05031_),
    .B1(_04883_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(_04891_),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_nor2_1 _22449_ (.A(_04881_),
    .B(_05031_),
    .Y(_05032_));
 sg13g2_a21oi_1 _22450_ (.A1(_05021_),
    .A2(_05030_),
    .Y(_05033_),
    .B1(_05032_));
 sg13g2_nand3_1 _22451_ (.B(_05020_),
    .C(_05033_),
    .A(_05010_),
    .Y(_05034_));
 sg13g2_a22oi_1 _22452_ (.Y(_05035_),
    .B1(_02905_),
    .B2(\cpu.dcache.r_data[7][15] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[6][15] ));
 sg13g2_a22oi_1 _22453_ (.Y(_05036_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[5][15] ),
    .A2(_09394_),
    .A1(\cpu.dcache.r_data[4][15] ));
 sg13g2_mux2_1 _22454_ (.A0(\cpu.dcache.r_data[1][15] ),
    .A1(\cpu.dcache.r_data[3][15] ),
    .S(net681),
    .X(_05037_));
 sg13g2_a22oi_1 _22455_ (.Y(_05038_),
    .B1(_05037_),
    .B2(net784),
    .A2(_09264_),
    .A1(\cpu.dcache.r_data[2][15] ));
 sg13g2_nand2b_1 _22456_ (.Y(_05039_),
    .B(net1025),
    .A_N(_05038_));
 sg13g2_and4_1 _22457_ (.A(_04807_),
    .B(_05035_),
    .C(_05036_),
    .D(_05039_),
    .X(_05040_));
 sg13g2_a21oi_1 _22458_ (.A1(_00155_),
    .A2(net550),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_nand2_1 _22459_ (.Y(_05042_),
    .A(net885),
    .B(_05041_));
 sg13g2_a21oi_2 _22460_ (.B1(net1110),
    .Y(_05043_),
    .A2(_08768_),
    .A1(net1032));
 sg13g2_nor2_1 _22461_ (.A(_05043_),
    .B(_04821_),
    .Y(_05044_));
 sg13g2_inv_1 _22462_ (.Y(_05045_),
    .A(_00154_));
 sg13g2_a22oi_1 _22463_ (.Y(_05046_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[1][31] ),
    .A2(net548),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_a22oi_1 _22464_ (.Y(_05047_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[7][31] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][31] ));
 sg13g2_mux2_1 _22465_ (.A0(\cpu.dcache.r_data[4][31] ),
    .A1(\cpu.dcache.r_data[6][31] ),
    .S(_09092_),
    .X(_05048_));
 sg13g2_a22oi_1 _22466_ (.Y(_05049_),
    .B1(_05048_),
    .B2(net892),
    .A2(net773),
    .A1(\cpu.dcache.r_data[5][31] ));
 sg13g2_nand2b_1 _22467_ (.Y(_05050_),
    .B(_09814_),
    .A_N(_05049_));
 sg13g2_nand4_1 _22468_ (.B(_05046_),
    .C(_05047_),
    .A(net403),
    .Y(_05051_),
    .D(_05050_));
 sg13g2_o21ai_1 _22469_ (.B1(_05051_),
    .Y(_05052_),
    .A1(_05045_),
    .A2(net403));
 sg13g2_nand3_1 _22470_ (.B(_05044_),
    .C(_05052_),
    .A(_05042_),
    .Y(_05053_));
 sg13g2_nor3_2 _22471_ (.A(_08766_),
    .B(net1031),
    .C(_08772_),
    .Y(_05054_));
 sg13g2_a22oi_1 _22472_ (.Y(_05055_),
    .B1(net493),
    .B2(\cpu.dcache.r_data[1][7] ),
    .A2(net548),
    .A1(\cpu.dcache.r_data[2][7] ));
 sg13g2_a22oi_1 _22473_ (.Y(_05056_),
    .B1(net612),
    .B2(\cpu.dcache.r_data[6][7] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][7] ));
 sg13g2_mux2_1 _22474_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(net681),
    .X(_05057_));
 sg13g2_a22oi_1 _22475_ (.Y(_05058_),
    .B1(_05057_),
    .B2(net682),
    .A2(net673),
    .A1(\cpu.dcache.r_data[4][7] ));
 sg13g2_nand2b_1 _22476_ (.Y(_05059_),
    .B(net772),
    .A_N(_05058_));
 sg13g2_and4_1 _22477_ (.A(net403),
    .B(_05055_),
    .C(_05056_),
    .D(_05059_),
    .X(_05060_));
 sg13g2_a21oi_2 _22478_ (.B1(_05060_),
    .Y(_05061_),
    .A2(net550),
    .A1(_00152_));
 sg13g2_nand2_1 _22479_ (.Y(_05062_),
    .A(_05042_),
    .B(_05044_));
 sg13g2_o21ai_1 _22480_ (.B1(_05062_),
    .Y(_05063_),
    .A1(_05054_),
    .A2(_05061_));
 sg13g2_nand2_1 _22481_ (.Y(_05064_),
    .A(_11790_),
    .B(net636));
 sg13g2_inv_1 _22482_ (.Y(_05065_),
    .A(_05064_));
 sg13g2_a22oi_1 _22483_ (.Y(_05066_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[5][23] ),
    .A2(net493),
    .A1(\cpu.dcache.r_data[1][23] ));
 sg13g2_a22oi_1 _22484_ (.Y(_05067_),
    .B1(net546),
    .B2(\cpu.dcache.r_data[3][23] ),
    .A2(net548),
    .A1(\cpu.dcache.r_data[2][23] ));
 sg13g2_mux2_1 _22485_ (.A0(\cpu.dcache.r_data[4][23] ),
    .A1(\cpu.dcache.r_data[6][23] ),
    .S(net619),
    .X(_05068_));
 sg13g2_a22oi_1 _22486_ (.Y(_05069_),
    .B1(_05068_),
    .B2(net892),
    .A2(net765),
    .A1(\cpu.dcache.r_data[7][23] ));
 sg13g2_nand2b_1 _22487_ (.Y(_05070_),
    .B(net670),
    .A_N(_05069_));
 sg13g2_and4_1 _22488_ (.A(net403),
    .B(_05066_),
    .C(_05067_),
    .D(_05070_),
    .X(_05071_));
 sg13g2_a21oi_1 _22489_ (.A1(_00153_),
    .A2(net550),
    .Y(_05072_),
    .B1(_05071_));
 sg13g2_a21oi_1 _22490_ (.A1(net885),
    .A2(_05061_),
    .Y(_05073_),
    .B1(_08771_));
 sg13g2_nor2_1 _22491_ (.A(net636),
    .B(_05073_),
    .Y(_05074_));
 sg13g2_a221oi_1 _22492_ (.B2(_09117_),
    .C1(_05074_),
    .B1(_05072_),
    .A1(_05061_),
    .Y(_05075_),
    .A2(_05065_));
 sg13g2_a21oi_1 _22493_ (.A1(_11790_),
    .A2(_05063_),
    .Y(_05076_),
    .B1(_05075_));
 sg13g2_and3_1 _22494_ (.X(_05077_),
    .A(net886),
    .B(_05053_),
    .C(_05076_));
 sg13g2_a21oi_2 _22495_ (.B1(_05077_),
    .Y(_05078_),
    .A2(_05034_),
    .A1(net1031));
 sg13g2_inv_1 _22496_ (.Y(_05079_),
    .A(_05078_));
 sg13g2_nor2_1 _22497_ (.A(net1033),
    .B(_05079_),
    .Y(_05080_));
 sg13g2_buf_1 _22498_ (.A(net513),
    .X(_05081_));
 sg13g2_buf_1 _22499_ (.A(net550),
    .X(_05082_));
 sg13g2_buf_1 _22500_ (.A(net365),
    .X(_05083_));
 sg13g2_a22oi_1 _22501_ (.Y(_05084_),
    .B1(net372),
    .B2(\cpu.dcache.r_data[1][10] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][10] ));
 sg13g2_a22oi_1 _22502_ (.Y(_05085_),
    .B1(_02903_),
    .B2(\cpu.dcache.r_data[6][10] ),
    .A2(net414),
    .A1(\cpu.dcache.r_data[3][10] ));
 sg13g2_mux2_1 _22503_ (.A0(\cpu.dcache.r_data[5][10] ),
    .A1(\cpu.dcache.r_data[7][10] ),
    .S(net496),
    .X(_05086_));
 sg13g2_a22oi_1 _22504_ (.Y(_05087_),
    .B1(_05086_),
    .B2(net620),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][10] ));
 sg13g2_nand2b_1 _22505_ (.Y(_05088_),
    .B(net537),
    .A_N(_05087_));
 sg13g2_and4_1 _22506_ (.A(net332),
    .B(_05084_),
    .C(_05085_),
    .D(_05088_),
    .X(_05089_));
 sg13g2_a21oi_1 _22507_ (.A1(_00103_),
    .A2(net459),
    .Y(_05090_),
    .B1(_05089_));
 sg13g2_a22oi_1 _22508_ (.Y(_05091_),
    .B1(net372),
    .B2(\cpu.dcache.r_data[1][26] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][26] ));
 sg13g2_a22oi_1 _22509_ (.Y(_05092_),
    .B1(net475),
    .B2(\cpu.dcache.r_data[6][26] ),
    .A2(net414),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_mux2_1 _22510_ (.A0(\cpu.dcache.r_data[5][26] ),
    .A1(\cpu.dcache.r_data[7][26] ),
    .S(net496),
    .X(_05093_));
 sg13g2_a22oi_1 _22511_ (.Y(_05094_),
    .B1(_05093_),
    .B2(net620),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][26] ));
 sg13g2_nand2b_1 _22512_ (.Y(_05095_),
    .B(_11719_),
    .A_N(_05094_));
 sg13g2_and4_1 _22513_ (.A(_05083_),
    .B(_05091_),
    .C(_05092_),
    .D(_05095_),
    .X(_05096_));
 sg13g2_a21oi_1 _22514_ (.A1(_00102_),
    .A2(net459),
    .Y(_05097_),
    .B1(_05096_));
 sg13g2_buf_1 _22515_ (.A(net668),
    .X(_05098_));
 sg13g2_mux2_1 _22516_ (.A0(_05090_),
    .A1(_05097_),
    .S(net580),
    .X(_05099_));
 sg13g2_nor3_1 _22517_ (.A(net886),
    .B(_09821_),
    .C(_04875_),
    .Y(_05100_));
 sg13g2_buf_2 _22518_ (.A(_05100_),
    .X(_05101_));
 sg13g2_nor2_1 _22519_ (.A(net898),
    .B(_09817_),
    .Y(_05102_));
 sg13g2_buf_1 _22520_ (.A(_05102_),
    .X(_05103_));
 sg13g2_buf_1 _22521_ (.A(_05103_),
    .X(_05104_));
 sg13g2_a22oi_1 _22522_ (.Y(_05105_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_reload[10] ),
    .A2(net362),
    .A1(\cpu.intr.r_timer_count[10] ));
 sg13g2_nor2_1 _22523_ (.A(net1036),
    .B(net597),
    .Y(_05106_));
 sg13g2_buf_1 _22524_ (.A(_05106_),
    .X(_05107_));
 sg13g2_a22oi_1 _22525_ (.Y(_05108_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[10] ),
    .A2(net462),
    .A1(_10015_));
 sg13g2_buf_1 _22526_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05109_));
 sg13g2_buf_1 _22527_ (.A(_04935_),
    .X(_05110_));
 sg13g2_a22oi_1 _22528_ (.Y(_05111_),
    .B1(net396),
    .B2(\cpu.intr.r_clock_cmp[26] ),
    .A2(net375),
    .A1(_05109_));
 sg13g2_nand3_1 _22529_ (.B(_05108_),
    .C(_05111_),
    .A(_05105_),
    .Y(_05112_));
 sg13g2_buf_1 _22530_ (.A(_08768_),
    .X(_05113_));
 sg13g2_a221oi_1 _22531_ (.B2(_05112_),
    .C1(net943),
    .B1(_05101_),
    .A1(net460),
    .Y(_05114_),
    .A2(_05099_));
 sg13g2_o21ai_1 _22532_ (.B1(net32),
    .Y(_05115_),
    .A1(_05080_),
    .A2(_05114_));
 sg13g2_o21ai_1 _22533_ (.B1(_05115_),
    .Y(_05116_),
    .A1(net1089),
    .A2(net31));
 sg13g2_buf_1 _22534_ (.A(net153),
    .X(_05117_));
 sg13g2_nand2_1 _22535_ (.Y(_05118_),
    .A(_10183_),
    .B(_11357_));
 sg13g2_nor2_1 _22536_ (.A(net946),
    .B(_05118_),
    .Y(_05119_));
 sg13g2_a221oi_1 _22537_ (.B2(net128),
    .C1(_05119_),
    .B1(_05116_),
    .A1(_04989_),
    .Y(_01032_),
    .A2(_04991_));
 sg13g2_nand2b_1 _22538_ (.Y(_05120_),
    .B(net711),
    .A_N(_04222_));
 sg13g2_o21ai_1 _22539_ (.B1(_05120_),
    .Y(_05121_),
    .A1(_04792_),
    .A2(_04210_));
 sg13g2_a22oi_1 _22540_ (.Y(_05122_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net362),
    .A1(\cpu.intr.r_timer_count[11] ));
 sg13g2_a22oi_1 _22541_ (.Y(_05123_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_reload[11] ),
    .A2(net396),
    .A1(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_buf_1 _22542_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05124_));
 sg13g2_a22oi_1 _22543_ (.Y(_05125_),
    .B1(net462),
    .B2(_10020_),
    .A2(net429),
    .A1(_05124_));
 sg13g2_nand3_1 _22544_ (.B(_05123_),
    .C(_05125_),
    .A(_05122_),
    .Y(_05126_));
 sg13g2_a22oi_1 _22545_ (.Y(_05127_),
    .B1(net372),
    .B2(\cpu.dcache.r_data[1][11] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][11] ));
 sg13g2_a22oi_1 _22546_ (.Y(_05128_),
    .B1(net532),
    .B2(\cpu.dcache.r_data[6][11] ),
    .A2(net414),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_mux2_1 _22547_ (.A0(\cpu.dcache.r_data[5][11] ),
    .A1(\cpu.dcache.r_data[7][11] ),
    .S(net552),
    .X(_05129_));
 sg13g2_a22oi_1 _22548_ (.Y(_05130_),
    .B1(_05129_),
    .B2(net620),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][11] ));
 sg13g2_nand2b_1 _22549_ (.Y(_05131_),
    .B(net537),
    .A_N(_05130_));
 sg13g2_and4_1 _22550_ (.A(net332),
    .B(_05127_),
    .C(_05128_),
    .D(_05131_),
    .X(_05132_));
 sg13g2_a21oi_2 _22551_ (.B1(_05132_),
    .Y(_05133_),
    .A2(net459),
    .A1(_00113_));
 sg13g2_a22oi_1 _22552_ (.Y(_05134_),
    .B1(_02899_),
    .B2(\cpu.dcache.r_data[5][27] ),
    .A2(net416),
    .A1(\cpu.dcache.r_data[1][27] ));
 sg13g2_a22oi_1 _22553_ (.Y(_05135_),
    .B1(_04799_),
    .B2(\cpu.dcache.r_data[3][27] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][27] ));
 sg13g2_mux2_1 _22554_ (.A0(\cpu.dcache.r_data[4][27] ),
    .A1(\cpu.dcache.r_data[6][27] ),
    .S(net514),
    .X(_05136_));
 sg13g2_a22oi_1 _22555_ (.Y(_05137_),
    .B1(_05136_),
    .B2(net713),
    .A2(_09815_),
    .A1(\cpu.dcache.r_data[7][27] ));
 sg13g2_nand2b_1 _22556_ (.Y(_05138_),
    .B(net603),
    .A_N(_05137_));
 sg13g2_and4_1 _22557_ (.A(_04808_),
    .B(_05134_),
    .C(_05135_),
    .D(_05138_),
    .X(_05139_));
 sg13g2_a21oi_1 _22558_ (.A1(_00112_),
    .A2(net463),
    .Y(_05140_),
    .B1(_05139_));
 sg13g2_mux2_1 _22559_ (.A0(_05133_),
    .A1(_05140_),
    .S(net580),
    .X(_05141_));
 sg13g2_a22oi_1 _22560_ (.Y(_05142_),
    .B1(_05141_),
    .B2(net460),
    .A2(_05126_),
    .A1(_05101_));
 sg13g2_a21oi_2 _22561_ (.B1(_11357_),
    .Y(_05143_),
    .A2(_05079_),
    .A1(net943));
 sg13g2_o21ai_1 _22562_ (.B1(_05143_),
    .Y(_05144_),
    .A1(net943),
    .A2(_05142_));
 sg13g2_o21ai_1 _22563_ (.B1(_05144_),
    .Y(_05145_),
    .A1(\cpu.ex.pc[11] ),
    .A2(_05118_));
 sg13g2_nor2_1 _22564_ (.A(_03448_),
    .B(_05145_),
    .Y(_05146_));
 sg13g2_a21oi_1 _22565_ (.A1(_02925_),
    .A2(_03448_),
    .Y(_05147_),
    .B1(_05146_));
 sg13g2_a21oi_1 _22566_ (.A1(_04989_),
    .A2(_05121_),
    .Y(_01033_),
    .B1(_05147_));
 sg13g2_a22oi_1 _22567_ (.Y(_05148_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net362),
    .A1(_09824_));
 sg13g2_a22oi_1 _22568_ (.Y(_05149_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_reload[12] ),
    .A2(net462),
    .A1(_10027_));
 sg13g2_buf_2 _22569_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05150_));
 sg13g2_a22oi_1 _22570_ (.Y(_05151_),
    .B1(net396),
    .B2(\cpu.intr.r_clock_cmp[28] ),
    .A2(net429),
    .A1(_05150_));
 sg13g2_nand3_1 _22571_ (.B(_05149_),
    .C(_05151_),
    .A(_05148_),
    .Y(_05152_));
 sg13g2_inv_1 _22572_ (.Y(_05153_),
    .A(_00124_));
 sg13g2_buf_1 _22573_ (.A(net403),
    .X(_05154_));
 sg13g2_buf_1 _22574_ (.A(_02892_),
    .X(_05155_));
 sg13g2_a22oi_1 _22575_ (.Y(_05156_),
    .B1(net364),
    .B2(\cpu.dcache.r_data[1][12] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][12] ));
 sg13g2_a22oi_1 _22576_ (.Y(_05157_),
    .B1(net532),
    .B2(\cpu.dcache.r_data[6][12] ),
    .A2(net477),
    .A1(\cpu.dcache.r_data[3][12] ));
 sg13g2_mux2_1 _22577_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(\cpu.dcache.r_data[7][12] ),
    .S(net514),
    .X(_05158_));
 sg13g2_a22oi_1 _22578_ (.Y(_05159_),
    .B1(_05158_),
    .B2(_09085_),
    .A2(net673),
    .A1(\cpu.dcache.r_data[4][12] ));
 sg13g2_nand2b_1 _22579_ (.Y(_05160_),
    .B(net603),
    .A_N(_05159_));
 sg13g2_nand4_1 _22580_ (.B(_05156_),
    .C(_05157_),
    .A(net365),
    .Y(_05161_),
    .D(_05160_));
 sg13g2_o21ai_1 _22581_ (.B1(_05161_),
    .Y(_05162_),
    .A1(_05153_),
    .A2(net360));
 sg13g2_a22oi_1 _22582_ (.Y(_05163_),
    .B1(_09346_),
    .B2(\cpu.dcache.r_data[5][28] ),
    .A2(_02887_),
    .A1(\cpu.dcache.r_data[1][28] ));
 sg13g2_a22oi_1 _22583_ (.Y(_05164_),
    .B1(_04799_),
    .B2(\cpu.dcache.r_data[3][28] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][28] ));
 sg13g2_mux2_1 _22584_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(\cpu.dcache.r_data[6][28] ),
    .S(net619),
    .X(_05165_));
 sg13g2_a22oi_1 _22585_ (.Y(_05166_),
    .B1(_05165_),
    .B2(net713),
    .A2(net669),
    .A1(\cpu.dcache.r_data[7][28] ));
 sg13g2_nand2b_1 _22586_ (.Y(_05167_),
    .B(_09814_),
    .A_N(_05166_));
 sg13g2_and4_1 _22587_ (.A(_04807_),
    .B(_05163_),
    .C(_05164_),
    .D(_05167_),
    .X(_05168_));
 sg13g2_a21oi_2 _22588_ (.B1(_05168_),
    .Y(_05169_),
    .A2(_04823_),
    .A1(_00123_));
 sg13g2_nand2_1 _22589_ (.Y(_05170_),
    .A(net668),
    .B(_05169_));
 sg13g2_o21ai_1 _22590_ (.B1(_05170_),
    .Y(_05171_),
    .A1(net580),
    .A2(_05162_));
 sg13g2_a22oi_1 _22591_ (.Y(_05172_),
    .B1(_05171_),
    .B2(net460),
    .A2(_05152_),
    .A1(_05101_));
 sg13g2_or2_1 _22592_ (.X(_05173_),
    .B(_05172_),
    .A(net943));
 sg13g2_nand3_1 _22593_ (.B(_05143_),
    .C(_05173_),
    .A(net32),
    .Y(_05174_));
 sg13g2_o21ai_1 _22594_ (.B1(_05174_),
    .Y(_05175_),
    .A1(net675),
    .A2(net31));
 sg13g2_buf_1 _22595_ (.A(_11348_),
    .X(_05176_));
 sg13g2_and2_1 _22596_ (.A(net710),
    .B(_04226_),
    .X(_05177_));
 sg13g2_a21oi_1 _22597_ (.A1(net635),
    .A2(_04268_),
    .Y(_05178_),
    .B1(_05177_));
 sg13g2_buf_1 _22598_ (.A(_04125_),
    .X(_05179_));
 sg13g2_nor3_1 _22599_ (.A(_08363_),
    .B(net231),
    .C(net153),
    .Y(_05180_));
 sg13g2_a221oi_1 _22600_ (.B2(_04989_),
    .C1(_05180_),
    .B1(_05178_),
    .A1(net128),
    .Y(_01034_),
    .A2(_05175_));
 sg13g2_a22oi_1 _22601_ (.Y(_05181_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net362),
    .A1(\cpu.intr.r_timer_count[13] ));
 sg13g2_a22oi_1 _22602_ (.Y(_05182_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_reload[13] ),
    .A2(net462),
    .A1(_10032_));
 sg13g2_buf_1 _22603_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05183_));
 sg13g2_a22oi_1 _22604_ (.Y(_05184_),
    .B1(net396),
    .B2(\cpu.intr.r_clock_cmp[29] ),
    .A2(net375),
    .A1(_05183_));
 sg13g2_nand3_1 _22605_ (.B(_05182_),
    .C(_05184_),
    .A(_05181_),
    .Y(_05185_));
 sg13g2_inv_1 _22606_ (.Y(_05186_),
    .A(_00131_));
 sg13g2_a22oi_1 _22607_ (.Y(_05187_),
    .B1(net364),
    .B2(\cpu.dcache.r_data[1][13] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][13] ));
 sg13g2_a22oi_1 _22608_ (.Y(_05188_),
    .B1(net532),
    .B2(\cpu.dcache.r_data[6][13] ),
    .A2(net477),
    .A1(\cpu.dcache.r_data[3][13] ));
 sg13g2_mux2_1 _22609_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(\cpu.dcache.r_data[7][13] ),
    .S(net552),
    .X(_05189_));
 sg13g2_a22oi_1 _22610_ (.Y(_05190_),
    .B1(_05189_),
    .B2(_09085_),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][13] ));
 sg13g2_nand2b_1 _22611_ (.Y(_05191_),
    .B(_11717_),
    .A_N(_05190_));
 sg13g2_nand4_1 _22612_ (.B(_05187_),
    .C(_05188_),
    .A(net365),
    .Y(_05192_),
    .D(_05191_));
 sg13g2_o21ai_1 _22613_ (.B1(_05192_),
    .Y(_05193_),
    .A1(_05186_),
    .A2(net360));
 sg13g2_inv_1 _22614_ (.Y(_05194_),
    .A(_00130_));
 sg13g2_a22oi_1 _22615_ (.Y(_05195_),
    .B1(_04824_),
    .B2(\cpu.dcache.r_data[1][29] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][29] ));
 sg13g2_a22oi_1 _22616_ (.Y(_05196_),
    .B1(_02902_),
    .B2(\cpu.dcache.r_data[6][29] ),
    .A2(net477),
    .A1(\cpu.dcache.r_data[3][29] ));
 sg13g2_mux2_1 _22617_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(\cpu.dcache.r_data[7][29] ),
    .S(_04802_),
    .X(_05197_));
 sg13g2_a22oi_1 _22618_ (.Y(_05198_),
    .B1(_05197_),
    .B2(net682),
    .A2(_11762_),
    .A1(\cpu.dcache.r_data[4][29] ));
 sg13g2_nand2b_1 _22619_ (.Y(_05199_),
    .B(_11717_),
    .A_N(_05198_));
 sg13g2_nand4_1 _22620_ (.B(_05195_),
    .C(_05196_),
    .A(_04808_),
    .Y(_05200_),
    .D(_05199_));
 sg13g2_o21ai_1 _22621_ (.B1(_05200_),
    .Y(_05201_),
    .A1(_05194_),
    .A2(net360));
 sg13g2_or2_1 _22622_ (.X(_05202_),
    .B(_05201_),
    .A(net759));
 sg13g2_o21ai_1 _22623_ (.B1(_05202_),
    .Y(_05203_),
    .A1(net580),
    .A2(_05193_));
 sg13g2_a22oi_1 _22624_ (.Y(_05204_),
    .B1(_05203_),
    .B2(net460),
    .A2(_05185_),
    .A1(_05101_));
 sg13g2_o21ai_1 _22625_ (.B1(_05143_),
    .Y(_05205_),
    .A1(net943),
    .A2(_05204_));
 sg13g2_mux2_1 _22626_ (.A0(_05205_),
    .A1(net611),
    .S(_03448_),
    .X(_05206_));
 sg13g2_o21ai_1 _22627_ (.B1(_05206_),
    .Y(_05207_),
    .A1(_08411_),
    .A2(_05118_));
 sg13g2_o21ai_1 _22628_ (.B1(net635),
    .Y(_05208_),
    .A1(net233),
    .A2(\cpu.ex.c_mult[13] ));
 sg13g2_and2_1 _22629_ (.A(_04984_),
    .B(_04322_),
    .X(_05209_));
 sg13g2_nor3_1 _22630_ (.A(_04988_),
    .B(_11360_),
    .C(_05209_),
    .Y(_05210_));
 sg13g2_o21ai_1 _22631_ (.B1(_05210_),
    .Y(_05211_),
    .A1(_04317_),
    .A2(_05208_));
 sg13g2_nor2b_1 _22632_ (.A(_05207_),
    .B_N(_05211_),
    .Y(_01035_));
 sg13g2_o21ai_1 _22633_ (.B1(_04125_),
    .Y(_05212_),
    .A1(_11348_),
    .A2(_04366_));
 sg13g2_o21ai_1 _22634_ (.B1(_05212_),
    .Y(_05213_),
    .A1(_08599_),
    .A2(_04125_));
 sg13g2_a22oi_1 _22635_ (.Y(_05214_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[14] ),
    .A2(_04951_),
    .A1(\cpu.intr.r_timer_count[14] ));
 sg13g2_a22oi_1 _22636_ (.Y(_05215_),
    .B1(_05104_),
    .B2(\cpu.intr.r_timer_reload[14] ),
    .A2(net462),
    .A1(_10038_));
 sg13g2_buf_1 _22637_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05216_));
 sg13g2_a22oi_1 _22638_ (.Y(_05217_),
    .B1(_05110_),
    .B2(\cpu.intr.r_clock_cmp[30] ),
    .A2(net375),
    .A1(_05216_));
 sg13g2_nand3_1 _22639_ (.B(_05215_),
    .C(_05217_),
    .A(_05214_),
    .Y(_05218_));
 sg13g2_a22oi_1 _22640_ (.Y(_05219_),
    .B1(_02888_),
    .B2(\cpu.dcache.r_data[1][14] ),
    .A2(_02893_),
    .A1(\cpu.dcache.r_data[2][14] ));
 sg13g2_a22oi_1 _22641_ (.Y(_05220_),
    .B1(_02902_),
    .B2(\cpu.dcache.r_data[6][14] ),
    .A2(_02896_),
    .A1(\cpu.dcache.r_data[3][14] ));
 sg13g2_mux2_1 _22642_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(\cpu.dcache.r_data[7][14] ),
    .S(_09093_),
    .X(_05221_));
 sg13g2_a22oi_1 _22643_ (.Y(_05222_),
    .B1(_05221_),
    .B2(_09086_),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][14] ));
 sg13g2_nand2b_1 _22644_ (.Y(_05223_),
    .B(net537),
    .A_N(_05222_));
 sg13g2_and4_1 _22645_ (.A(_05083_),
    .B(_05219_),
    .C(_05220_),
    .D(_05223_),
    .X(_05224_));
 sg13g2_a21oi_1 _22646_ (.A1(_00143_),
    .A2(net459),
    .Y(_05225_),
    .B1(_05224_));
 sg13g2_nand2_1 _22647_ (.Y(_05226_),
    .A(_09813_),
    .B(_05225_));
 sg13g2_a22oi_1 _22648_ (.Y(_05227_),
    .B1(_02888_),
    .B2(\cpu.dcache.r_data[1][30] ),
    .A2(_02893_),
    .A1(\cpu.dcache.r_data[2][30] ));
 sg13g2_a22oi_1 _22649_ (.Y(_05228_),
    .B1(_02903_),
    .B2(\cpu.dcache.r_data[6][30] ),
    .A2(_02896_),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_mux2_1 _22650_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(\cpu.dcache.r_data[7][30] ),
    .S(_09093_),
    .X(_05229_));
 sg13g2_a22oi_1 _22651_ (.Y(_05230_),
    .B1(_05229_),
    .B2(_09086_),
    .A2(_11762_),
    .A1(\cpu.dcache.r_data[4][30] ));
 sg13g2_nand2b_1 _22652_ (.Y(_05231_),
    .B(_11718_),
    .A_N(_05230_));
 sg13g2_and4_1 _22653_ (.A(net332),
    .B(_05227_),
    .C(_05228_),
    .D(_05231_),
    .X(_05232_));
 sg13g2_a21oi_1 _22654_ (.A1(_00142_),
    .A2(_05082_),
    .Y(_05233_),
    .B1(_05232_));
 sg13g2_nand2_1 _22655_ (.Y(_05234_),
    .A(net580),
    .B(_05233_));
 sg13g2_nand2_1 _22656_ (.Y(_05235_),
    .A(_05226_),
    .B(_05234_));
 sg13g2_a22oi_1 _22657_ (.Y(_05236_),
    .B1(_05235_),
    .B2(net460),
    .A2(_05218_),
    .A1(_05101_));
 sg13g2_o21ai_1 _22658_ (.B1(_05143_),
    .Y(_05237_),
    .A1(_05113_),
    .A2(_05236_));
 sg13g2_mux2_1 _22659_ (.A0(_05237_),
    .A1(net672),
    .S(_03448_),
    .X(_05238_));
 sg13g2_o21ai_1 _22660_ (.B1(_05238_),
    .Y(_05239_),
    .A1(_04983_),
    .A2(_05213_));
 sg13g2_a21oi_1 _22661_ (.A1(_04364_),
    .A2(_04794_),
    .Y(_01036_),
    .B1(_05239_));
 sg13g2_nand2_1 _22662_ (.Y(_05240_),
    .A(net635),
    .B(_04417_));
 sg13g2_a21oi_1 _22663_ (.A1(net711),
    .A2(_04420_),
    .Y(_05241_),
    .B1(_04793_));
 sg13g2_a22oi_1 _22664_ (.Y(_05242_),
    .B1(_05104_),
    .B2(\cpu.intr.r_timer_reload[15] ),
    .A2(_04951_),
    .A1(\cpu.intr.r_timer_count[15] ));
 sg13g2_a22oi_1 _22665_ (.Y(_05243_),
    .B1(_05110_),
    .B2(\cpu.intr.r_clock_cmp[31] ),
    .A2(net462),
    .A1(_10045_));
 sg13g2_buf_1 _22666_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05244_));
 sg13g2_a22oi_1 _22667_ (.Y(_05245_),
    .B1(_05107_),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net375),
    .A1(_05244_));
 sg13g2_nand3_1 _22668_ (.B(_05243_),
    .C(_05245_),
    .A(_05242_),
    .Y(_05246_));
 sg13g2_o21ai_1 _22669_ (.B1(_05042_),
    .Y(_05247_),
    .A1(net667),
    .A2(_05052_));
 sg13g2_a22oi_1 _22670_ (.Y(_05248_),
    .B1(_05247_),
    .B2(net460),
    .A2(_05246_),
    .A1(_05101_));
 sg13g2_o21ai_1 _22671_ (.B1(_05143_),
    .Y(_05249_),
    .A1(_05113_),
    .A2(_05248_));
 sg13g2_mux2_1 _22672_ (.A0(_05249_),
    .A1(net890),
    .S(_03448_),
    .X(_05250_));
 sg13g2_o21ai_1 _22673_ (.B1(_05250_),
    .Y(_05251_),
    .A1(_08379_),
    .A2(_05118_));
 sg13g2_a21oi_1 _22674_ (.A1(_05240_),
    .A2(_05241_),
    .Y(_01037_),
    .B1(_05251_));
 sg13g2_buf_1 _22675_ (.A(_11357_),
    .X(_05252_));
 sg13g2_mux2_1 _22676_ (.A0(_10206_),
    .A1(_04122_),
    .S(_11348_),
    .X(_05253_));
 sg13g2_nor2_1 _22677_ (.A(net913),
    .B(net231),
    .Y(_05254_));
 sg13g2_a21oi_1 _22678_ (.A1(_05179_),
    .A2(_05253_),
    .Y(_05255_),
    .B1(_05254_));
 sg13g2_nand2_1 _22679_ (.Y(_05256_),
    .A(\cpu.dcache.r_data[3][1] ),
    .B(net477));
 sg13g2_a22oi_1 _22680_ (.Y(_05257_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[7][1] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][1] ));
 sg13g2_nand3_1 _22681_ (.B(net1025),
    .C(\cpu.dcache.r_data[1][1] ),
    .A(net682),
    .Y(_05258_));
 sg13g2_o21ai_1 _22682_ (.B1(_05258_),
    .Y(_05259_),
    .A1(net682),
    .A2(_12360_));
 sg13g2_a22oi_1 _22683_ (.Y(_05260_),
    .B1(net773),
    .B2(\cpu.dcache.r_data[5][1] ),
    .A2(net894),
    .A1(\cpu.dcache.r_data[6][1] ));
 sg13g2_inv_1 _22684_ (.Y(_05261_),
    .A(_05260_));
 sg13g2_a22oi_1 _22685_ (.Y(_05262_),
    .B1(_05261_),
    .B2(net603),
    .A2(_05259_),
    .A1(net780));
 sg13g2_nand4_1 _22686_ (.B(_05256_),
    .C(_05257_),
    .A(net360),
    .Y(_05263_),
    .D(_05262_));
 sg13g2_o21ai_1 _22687_ (.B1(_05263_),
    .Y(_05264_),
    .A1(\cpu.dcache.r_data[0][1] ),
    .A2(net360));
 sg13g2_nand2_1 _22688_ (.Y(_05265_),
    .A(\cpu.dcache.r_data[3][17] ),
    .B(net464));
 sg13g2_a22oi_1 _22689_ (.Y(_05266_),
    .B1(_09394_),
    .B2(\cpu.dcache.r_data[4][17] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][17] ));
 sg13g2_a22oi_1 _22690_ (.Y(_05267_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[7][17] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[6][17] ));
 sg13g2_a22oi_1 _22691_ (.Y(_05268_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[5][17] ),
    .A2(net416),
    .A1(\cpu.dcache.r_data[1][17] ));
 sg13g2_nand4_1 _22692_ (.B(_05266_),
    .C(_05267_),
    .A(_05265_),
    .Y(_05269_),
    .D(_05268_));
 sg13g2_nand2_1 _22693_ (.Y(_05270_),
    .A(_00091_),
    .B(net550));
 sg13g2_o21ai_1 _22694_ (.B1(_05270_),
    .Y(_05271_),
    .A1(net463),
    .A2(_05269_));
 sg13g2_or2_1 _22695_ (.X(_05272_),
    .B(_05271_),
    .A(_09812_));
 sg13g2_o21ai_1 _22696_ (.B1(_05272_),
    .Y(_05273_),
    .A1(net580),
    .A2(_05264_));
 sg13g2_a22oi_1 _22697_ (.Y(_05274_),
    .B1(_02900_),
    .B2(\cpu.dcache.r_data[5][25] ),
    .A2(net364),
    .A1(\cpu.dcache.r_data[1][25] ));
 sg13g2_a22oi_1 _22698_ (.Y(_05275_),
    .B1(_02895_),
    .B2(\cpu.dcache.r_data[3][25] ),
    .A2(_05155_),
    .A1(\cpu.dcache.r_data[2][25] ));
 sg13g2_mux2_1 _22699_ (.A0(\cpu.dcache.r_data[4][25] ),
    .A1(\cpu.dcache.r_data[6][25] ),
    .S(net552),
    .X(_05276_));
 sg13g2_a22oi_1 _22700_ (.Y(_05277_),
    .B1(_05276_),
    .B2(net638),
    .A2(_09815_),
    .A1(\cpu.dcache.r_data[7][25] ));
 sg13g2_nand2b_1 _22701_ (.Y(_05278_),
    .B(_11718_),
    .A_N(_05277_));
 sg13g2_and4_1 _22702_ (.A(_05154_),
    .B(_05274_),
    .C(_05275_),
    .D(_05278_),
    .X(_05279_));
 sg13g2_a21oi_1 _22703_ (.A1(_00092_),
    .A2(_05082_),
    .Y(_05280_),
    .B1(_05279_));
 sg13g2_inv_1 _22704_ (.Y(_05281_),
    .A(_00093_));
 sg13g2_a22oi_1 _22705_ (.Y(_05282_),
    .B1(_02899_),
    .B2(\cpu.dcache.r_data[5][9] ),
    .A2(_04824_),
    .A1(\cpu.dcache.r_data[1][9] ));
 sg13g2_a22oi_1 _22706_ (.Y(_05283_),
    .B1(_02895_),
    .B2(\cpu.dcache.r_data[3][9] ),
    .A2(_05155_),
    .A1(\cpu.dcache.r_data[2][9] ));
 sg13g2_mux2_1 _22707_ (.A0(\cpu.dcache.r_data[4][9] ),
    .A1(\cpu.dcache.r_data[6][9] ),
    .S(net514),
    .X(_05284_));
 sg13g2_a22oi_1 _22708_ (.Y(_05285_),
    .B1(_05284_),
    .B2(_03698_),
    .A2(net669),
    .A1(\cpu.dcache.r_data[7][9] ));
 sg13g2_nand2b_1 _22709_ (.Y(_05286_),
    .B(net603),
    .A_N(_05285_));
 sg13g2_nand4_1 _22710_ (.B(_05282_),
    .C(_05283_),
    .A(net365),
    .Y(_05287_),
    .D(_05286_));
 sg13g2_o21ai_1 _22711_ (.B1(_05287_),
    .Y(_05288_),
    .A1(_05281_),
    .A2(_05154_));
 sg13g2_nor2_1 _22712_ (.A(_09118_),
    .B(_05288_),
    .Y(_05289_));
 sg13g2_a21oi_1 _22713_ (.A1(net991),
    .A2(_05280_),
    .Y(_05290_),
    .B1(_05289_));
 sg13g2_mux2_1 _22714_ (.A0(_05264_),
    .A1(_05272_),
    .S(net991),
    .X(_05291_));
 sg13g2_mux2_1 _22715_ (.A0(_05290_),
    .A1(_05291_),
    .S(net581),
    .X(_05292_));
 sg13g2_nor2_1 _22716_ (.A(net513),
    .B(_05292_),
    .Y(_05293_));
 sg13g2_a21oi_1 _22717_ (.A1(net513),
    .A2(_05273_),
    .Y(_05294_),
    .B1(_05293_));
 sg13g2_mux2_1 _22718_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(\cpu.intr.r_timer_reload[17] ),
    .S(net730),
    .X(_05295_));
 sg13g2_a22oi_1 _22719_ (.Y(_05296_),
    .B1(_05295_),
    .B2(net474),
    .A2(net402),
    .A1(_09036_));
 sg13g2_mux2_1 _22720_ (.A0(\cpu.intr.r_clock_cmp[1] ),
    .A1(\cpu.intr.r_clock_cmp[17] ),
    .S(net782),
    .X(_05297_));
 sg13g2_a22oi_1 _22721_ (.Y(_05298_),
    .B1(_05297_),
    .B2(net413),
    .A2(net401),
    .A1(_09037_));
 sg13g2_buf_1 _22722_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05299_));
 sg13g2_and2_1 _22723_ (.A(net898),
    .B(_09840_),
    .X(_05300_));
 sg13g2_a21oi_1 _22724_ (.A1(net885),
    .A2(_09826_),
    .Y(_05301_),
    .B1(_05300_));
 sg13g2_nor2_1 _22725_ (.A(net533),
    .B(_05301_),
    .Y(_05302_));
 sg13g2_a221oi_1 _22726_ (.B2(_09968_),
    .C1(_05302_),
    .B1(_04859_),
    .A1(_05299_),
    .Y(_05303_),
    .A2(net429));
 sg13g2_nand3_1 _22727_ (.B(_09037_),
    .C(net333),
    .A(_09036_),
    .Y(_05304_));
 sg13g2_nand4_1 _22728_ (.B(_05298_),
    .C(_05303_),
    .A(_05296_),
    .Y(_05305_),
    .D(_05304_));
 sg13g2_buf_1 _22729_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05306_));
 sg13g2_buf_1 _22730_ (.A(_05016_),
    .X(_05307_));
 sg13g2_mux2_1 _22731_ (.A0(_11705_),
    .A1(_11710_),
    .S(net995),
    .X(_05308_));
 sg13g2_a22oi_1 _22732_ (.Y(_05309_),
    .B1(_05308_),
    .B2(net400),
    .A2(_05014_),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_o21ai_1 _22733_ (.B1(_05309_),
    .Y(_05310_),
    .A1(_00095_),
    .A2(net310));
 sg13g2_a21oi_1 _22734_ (.A1(_05306_),
    .A2(_04971_),
    .Y(_05311_),
    .B1(_05310_));
 sg13g2_nor2_1 _22735_ (.A(_00094_),
    .B(_04968_),
    .Y(_05312_));
 sg13g2_a21oi_1 _22736_ (.A1(_11706_),
    .A2(_04918_),
    .Y(_05313_),
    .B1(_05312_));
 sg13g2_nand2_1 _22737_ (.Y(_05314_),
    .A(_09162_),
    .B(_04963_));
 sg13g2_nand3_1 _22738_ (.B(_05313_),
    .C(_05314_),
    .A(_05311_),
    .Y(_05315_));
 sg13g2_a22oi_1 _22739_ (.Y(_05316_),
    .B1(net400),
    .B2(\cpu.uart.r_div_value[1] ),
    .A2(net461),
    .A1(\cpu.uart.r_r_invert ));
 sg13g2_a22oi_1 _22740_ (.Y(_05317_),
    .B1(net399),
    .B2(\cpu.uart.r_div_value[9] ),
    .A2(net401),
    .A1(_09034_));
 sg13g2_nand2_1 _22741_ (.Y(_05318_),
    .A(_05316_),
    .B(_05317_));
 sg13g2_a21oi_1 _22742_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04883_),
    .Y(_05319_),
    .B1(_05318_));
 sg13g2_o21ai_1 _22743_ (.B1(net1031),
    .Y(_05320_),
    .A1(net512),
    .A2(_05319_));
 sg13g2_a221oi_1 _22744_ (.B2(_04978_),
    .C1(_05320_),
    .B1(_05315_),
    .A1(_04847_),
    .Y(_05321_),
    .A2(_05305_));
 sg13g2_and3_1 _22745_ (.X(_05322_),
    .A(_09042_),
    .B(_09043_),
    .C(_04914_));
 sg13g2_buf_2 _22746_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05323_));
 sg13g2_inv_1 _22747_ (.Y(_05324_),
    .A(_00097_));
 sg13g2_a22oi_1 _22748_ (.Y(_05325_),
    .B1(_04940_),
    .B2(_05324_),
    .A2(net398),
    .A1(_05323_));
 sg13g2_nor2b_1 _22749_ (.A(_00099_),
    .B_N(_04918_),
    .Y(_05326_));
 sg13g2_nand2_1 _22750_ (.Y(_05327_),
    .A(_04932_),
    .B(_04935_));
 sg13g2_nor2_1 _22751_ (.A(_00100_),
    .B(_05327_),
    .Y(_05328_));
 sg13g2_nand2_1 _22752_ (.Y(_05329_),
    .A(_04907_),
    .B(_04869_));
 sg13g2_nand2b_1 _22753_ (.Y(_05330_),
    .B(net397),
    .A_N(_00096_));
 sg13g2_o21ai_1 _22754_ (.B1(_05330_),
    .Y(_05331_),
    .A1(_00098_),
    .A2(_05329_));
 sg13g2_nor3_1 _22755_ (.A(_05326_),
    .B(_05328_),
    .C(_05331_),
    .Y(_05332_));
 sg13g2_a22oi_1 _22756_ (.Y(_05333_),
    .B1(_04930_),
    .B2(_09043_),
    .A2(_04923_),
    .A1(_09042_));
 sg13g2_nand3_1 _22757_ (.B(_05332_),
    .C(_05333_),
    .A(_05325_),
    .Y(_05334_));
 sg13g2_o21ai_1 _22758_ (.B1(_04901_),
    .Y(_05335_),
    .A1(_05322_),
    .A2(_05334_));
 sg13g2_a22oi_1 _22759_ (.Y(_05336_),
    .B1(_05321_),
    .B2(_05335_),
    .A2(_05294_),
    .A1(net886));
 sg13g2_nand2_1 _22760_ (.Y(_05337_),
    .A(net32),
    .B(_05336_));
 sg13g2_o21ai_1 _22761_ (.B1(_05337_),
    .Y(_05338_),
    .A1(_09975_),
    .A2(net31));
 sg13g2_nor2_1 _22762_ (.A(net152),
    .B(_05338_),
    .Y(_05339_));
 sg13g2_a21oi_1 _22763_ (.A1(net152),
    .A2(_05255_),
    .Y(_01038_),
    .B1(_05339_));
 sg13g2_buf_1 _22764_ (.A(net153),
    .X(_05340_));
 sg13g2_nand2_1 _22765_ (.Y(_05341_),
    .A(\cpu.dcache.r_data[3][2] ),
    .B(net414));
 sg13g2_a22oi_1 _22766_ (.Y(_05342_),
    .B1(net474),
    .B2(\cpu.dcache.r_data[7][2] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][2] ));
 sg13g2_nor2_1 _22767_ (.A(net712),
    .B(net780),
    .Y(_05343_));
 sg13g2_a22oi_1 _22768_ (.Y(_05344_),
    .B1(_05343_),
    .B2(\cpu.dcache.r_data[6][2] ),
    .A2(\cpu.dcache.r_data[4][2] ),
    .A1(net780));
 sg13g2_nor2_1 _22769_ (.A(net620),
    .B(_05344_),
    .Y(_05345_));
 sg13g2_a221oi_1 _22770_ (.B2(\cpu.dcache.r_data[5][2] ),
    .C1(_05345_),
    .B1(net413),
    .A1(\cpu.dcache.r_data[1][2] ),
    .Y(_05346_),
    .A2(net364));
 sg13g2_nand4_1 _22771_ (.B(_05341_),
    .C(_05342_),
    .A(net360),
    .Y(_05347_),
    .D(_05346_));
 sg13g2_o21ai_1 _22772_ (.B1(_05347_),
    .Y(_05348_),
    .A1(\cpu.dcache.r_data[0][2] ),
    .A2(net332));
 sg13g2_inv_1 _22773_ (.Y(_05349_),
    .A(_05348_));
 sg13g2_a22oi_1 _22774_ (.Y(_05350_),
    .B1(net476),
    .B2(\cpu.dcache.r_data[5][18] ),
    .A2(net364),
    .A1(\cpu.dcache.r_data[1][18] ));
 sg13g2_a22oi_1 _22775_ (.Y(_05351_),
    .B1(net477),
    .B2(\cpu.dcache.r_data[3][18] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][18] ));
 sg13g2_mux2_1 _22776_ (.A0(\cpu.dcache.r_data[4][18] ),
    .A1(\cpu.dcache.r_data[6][18] ),
    .S(net552),
    .X(_05352_));
 sg13g2_a22oi_1 _22777_ (.Y(_05353_),
    .B1(_05352_),
    .B2(net713),
    .A2(net669),
    .A1(\cpu.dcache.r_data[7][18] ));
 sg13g2_nand2b_1 _22778_ (.Y(_05354_),
    .B(net603),
    .A_N(_05353_));
 sg13g2_and4_1 _22779_ (.A(net360),
    .B(_05350_),
    .C(_05351_),
    .D(_05354_),
    .X(_05355_));
 sg13g2_a21oi_1 _22780_ (.A1(_00101_),
    .A2(net459),
    .Y(_05356_),
    .B1(_05355_));
 sg13g2_nand2_1 _22781_ (.Y(_05357_),
    .A(net668),
    .B(_05356_));
 sg13g2_nor2_1 _22782_ (.A(net945),
    .B(_05357_),
    .Y(_05358_));
 sg13g2_a21oi_1 _22783_ (.A1(net945),
    .A2(_05349_),
    .Y(_05359_),
    .B1(_05358_));
 sg13g2_a221oi_1 _22784_ (.B2(net991),
    .C1(net581),
    .B1(_05097_),
    .A1(net667),
    .Y(_05360_),
    .A2(_05090_));
 sg13g2_a21oi_1 _22785_ (.A1(net581),
    .A2(_05359_),
    .Y(_05361_),
    .B1(_05360_));
 sg13g2_o21ai_1 _22786_ (.B1(_05357_),
    .Y(_05362_),
    .A1(net609),
    .A2(_05348_));
 sg13g2_mux2_1 _22787_ (.A0(_05361_),
    .A1(_05362_),
    .S(net460),
    .X(_05363_));
 sg13g2_buf_1 _22788_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05364_));
 sg13g2_nand2_1 _22789_ (.Y(_05365_),
    .A(net864),
    .B(_11691_));
 sg13g2_o21ai_1 _22790_ (.B1(_05365_),
    .Y(_05366_),
    .A1(net864),
    .A2(_00282_));
 sg13g2_a22oi_1 _22791_ (.Y(_05367_),
    .B1(_05366_),
    .B2(net400),
    .A2(_05014_),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _22792_ (.B1(_05367_),
    .Y(_05368_),
    .A1(_00105_),
    .A2(net310));
 sg13g2_a21oi_1 _22793_ (.A1(_05364_),
    .A2(_04971_),
    .Y(_05369_),
    .B1(_05368_));
 sg13g2_nor2_1 _22794_ (.A(_00104_),
    .B(_04968_),
    .Y(_05370_));
 sg13g2_a21oi_1 _22795_ (.A1(_11716_),
    .A2(_04918_),
    .Y(_05371_),
    .B1(_05370_));
 sg13g2_nand2_1 _22796_ (.Y(_05372_),
    .A(_09166_),
    .B(_04963_));
 sg13g2_nand3_1 _22797_ (.B(_05371_),
    .C(_05372_),
    .A(_05369_),
    .Y(_05373_));
 sg13g2_and2_1 _22798_ (.A(\cpu.uart.r_in[2] ),
    .B(_04883_),
    .X(_05374_));
 sg13g2_a221oi_1 _22799_ (.B2(_09802_),
    .C1(_05374_),
    .B1(net399),
    .A1(\cpu.uart.r_div_value[2] ),
    .Y(_05375_),
    .A2(net363));
 sg13g2_o21ai_1 _22800_ (.B1(net854),
    .Y(_05376_),
    .A1(net512),
    .A2(_05375_));
 sg13g2_a21oi_1 _22801_ (.A1(_04978_),
    .A2(_05373_),
    .Y(_05377_),
    .B1(_05376_));
 sg13g2_a22oi_1 _22802_ (.Y(_05378_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_reload[2] ),
    .A2(net362),
    .A1(\cpu.intr.r_timer_count[2] ));
 sg13g2_nand2_1 _22803_ (.Y(_05379_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(net396));
 sg13g2_buf_1 _22804_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05380_));
 sg13g2_a22oi_1 _22805_ (.Y(_05381_),
    .B1(net402),
    .B2(_09030_),
    .A2(net375),
    .A1(_05380_));
 sg13g2_a21o_1 _22806_ (.A2(net333),
    .A1(_09030_),
    .B1(net401),
    .X(_05382_));
 sg13g2_a22oi_1 _22807_ (.Y(_05383_),
    .B1(net474),
    .B2(\cpu.intr.r_timer_reload[18] ),
    .A2(net475),
    .A1(_09842_));
 sg13g2_a221oi_1 _22808_ (.B2(\cpu.intr.r_clock_cmp[2] ),
    .C1(net730),
    .B1(net413),
    .A1(_09972_),
    .Y(_05384_),
    .A2(net598));
 sg13g2_a21oi_1 _22809_ (.A1(net668),
    .A2(_05383_),
    .Y(_05385_),
    .B1(_05384_));
 sg13g2_a21oi_1 _22810_ (.A1(\cpu.intr.r_enable[2] ),
    .A2(_05382_),
    .Y(_05386_),
    .B1(_05385_));
 sg13g2_nand4_1 _22811_ (.B(_05379_),
    .C(_05381_),
    .A(_05378_),
    .Y(_05387_),
    .D(_05386_));
 sg13g2_nand3_1 _22812_ (.B(_09045_),
    .C(_04914_),
    .A(_09044_),
    .Y(_05388_));
 sg13g2_buf_1 _22813_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05389_));
 sg13g2_inv_1 _22814_ (.Y(_05390_),
    .A(_00108_));
 sg13g2_a22oi_1 _22815_ (.Y(_05391_),
    .B1(_04942_),
    .B2(_05390_),
    .A2(net398),
    .A1(_05389_));
 sg13g2_inv_1 _22816_ (.Y(_05392_),
    .A(_00106_));
 sg13g2_a22oi_1 _22817_ (.Y(_05393_),
    .B1(_04930_),
    .B2(_09045_),
    .A2(net397),
    .A1(_05392_));
 sg13g2_inv_1 _22818_ (.Y(_05394_),
    .A(_00109_));
 sg13g2_inv_1 _22819_ (.Y(_05395_),
    .A(_00107_));
 sg13g2_a22oi_1 _22820_ (.Y(_05396_),
    .B1(_04940_),
    .B2(_05395_),
    .A2(_04923_),
    .A1(_09044_));
 sg13g2_o21ai_1 _22821_ (.B1(_05396_),
    .Y(_05397_),
    .A1(_00110_),
    .A2(_05327_));
 sg13g2_a21oi_1 _22822_ (.A1(_05394_),
    .A2(_04918_),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_nand4_1 _22823_ (.B(_05391_),
    .C(_05393_),
    .A(_05388_),
    .Y(_05399_),
    .D(_05398_));
 sg13g2_a22oi_1 _22824_ (.Y(_05400_),
    .B1(_05399_),
    .B2(_04901_),
    .A2(_05387_),
    .A1(_04847_));
 sg13g2_nand2_1 _22825_ (.Y(_05401_),
    .A(_05377_),
    .B(_05400_));
 sg13g2_o21ai_1 _22826_ (.B1(_05401_),
    .Y(_05402_),
    .A1(net854),
    .A2(_05363_));
 sg13g2_mux2_1 _22827_ (.A0(net638),
    .A1(_05402_),
    .S(net31),
    .X(_05403_));
 sg13g2_o21ai_1 _22828_ (.B1(_04125_),
    .Y(_05404_),
    .A1(net919),
    .A2(net635));
 sg13g2_nand3_1 _22829_ (.B(net919),
    .C(net710),
    .A(net796),
    .Y(_05405_));
 sg13g2_o21ai_1 _22830_ (.B1(_05405_),
    .Y(_05406_),
    .A1(net711),
    .A2(_04453_));
 sg13g2_a221oi_1 _22831_ (.B2(net231),
    .C1(net153),
    .B1(_05406_),
    .A1(net798),
    .Y(_05407_),
    .A2(_05404_));
 sg13g2_a21oi_1 _22832_ (.A1(net127),
    .A2(_05403_),
    .Y(_01039_),
    .B1(_05407_));
 sg13g2_nand2_1 _22833_ (.Y(_05408_),
    .A(net710),
    .B(_04495_));
 sg13g2_o21ai_1 _22834_ (.B1(_05408_),
    .Y(_05409_),
    .A1(net711),
    .A2(_04493_));
 sg13g2_nand2_1 _22835_ (.Y(_05410_),
    .A(_04984_),
    .B(_04213_));
 sg13g2_a21oi_1 _22836_ (.A1(net231),
    .A2(_05410_),
    .Y(_05411_),
    .B1(net918));
 sg13g2_a21oi_1 _22837_ (.A1(_05179_),
    .A2(_05409_),
    .Y(_05412_),
    .B1(_05411_));
 sg13g2_buf_1 _22838_ (.A(_11360_),
    .X(_05413_));
 sg13g2_and2_1 _22839_ (.A(_09160_),
    .B(_04963_),
    .X(_05414_));
 sg13g2_buf_1 _22840_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05415_));
 sg13g2_nor2_1 _22841_ (.A(_00115_),
    .B(net310),
    .Y(_05416_));
 sg13g2_a221oi_1 _22842_ (.B2(\cpu.spi.r_timeout[3] ),
    .C1(_05416_),
    .B1(_05014_),
    .A1(_05415_),
    .Y(_05417_),
    .A2(_04971_));
 sg13g2_o21ai_1 _22843_ (.B1(_05417_),
    .Y(_05418_),
    .A1(_00114_),
    .A2(_04968_));
 sg13g2_o21ai_1 _22844_ (.B1(_04978_),
    .Y(_05419_),
    .A1(_05414_),
    .A2(_05418_));
 sg13g2_nand3_1 _22845_ (.B(_09055_),
    .C(_04914_),
    .A(_09054_),
    .Y(_05420_));
 sg13g2_nand2_2 _22846_ (.Y(_05421_),
    .A(net898),
    .B(net413));
 sg13g2_nand2_1 _22847_ (.Y(_05422_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(_04859_));
 sg13g2_o21ai_1 _22848_ (.B1(_05422_),
    .Y(_05423_),
    .A1(_00119_),
    .A2(_05421_));
 sg13g2_nand2_1 _22849_ (.Y(_05424_),
    .A(net837),
    .B(_05423_));
 sg13g2_buf_1 _22850_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05425_));
 sg13g2_nand2_1 _22851_ (.Y(_05426_),
    .A(_05425_),
    .B(net398));
 sg13g2_o21ai_1 _22852_ (.B1(_05426_),
    .Y(_05427_),
    .A1(_00117_),
    .A2(_04939_));
 sg13g2_a221oi_1 _22853_ (.B2(_09055_),
    .C1(_05427_),
    .B1(_04930_),
    .A1(_09054_),
    .Y(_05428_),
    .A2(_04923_));
 sg13g2_inv_1 _22854_ (.Y(_05429_),
    .A(_00116_));
 sg13g2_inv_1 _22855_ (.Y(_05430_),
    .A(_00118_));
 sg13g2_a22oi_1 _22856_ (.Y(_05431_),
    .B1(_04942_),
    .B2(_05430_),
    .A2(_04928_),
    .A1(_05429_));
 sg13g2_nand4_1 _22857_ (.B(_05424_),
    .C(_05428_),
    .A(_05420_),
    .Y(_05432_),
    .D(_05431_));
 sg13g2_a22oi_1 _22858_ (.Y(_05433_),
    .B1(net474),
    .B2(\cpu.intr.r_timer_reload[19] ),
    .A2(net475),
    .A1(\cpu.intr.r_timer_count[19] ));
 sg13g2_a221oi_1 _22859_ (.B2(\cpu.intr.r_clock_cmp[3] ),
    .C1(net730),
    .B1(net413),
    .A1(_09978_),
    .Y(_05434_),
    .A2(net598));
 sg13g2_a21o_1 _22860_ (.A2(_05433_),
    .A1(net668),
    .B1(_05434_),
    .X(_05435_));
 sg13g2_buf_2 _22861_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05436_));
 sg13g2_and2_1 _22862_ (.A(_09031_),
    .B(net402),
    .X(_05437_));
 sg13g2_a221oi_1 _22863_ (.B2(\cpu.intr.r_timer_reload[3] ),
    .C1(_05437_),
    .B1(_05103_),
    .A1(_05436_),
    .Y(_05438_),
    .A2(net429));
 sg13g2_a22oi_1 _22864_ (.Y(_05439_),
    .B1(net396),
    .B2(\cpu.intr.r_clock_cmp[19] ),
    .A2(_04950_),
    .A1(\cpu.intr.r_timer_count[3] ));
 sg13g2_a21oi_1 _22865_ (.A1(_09031_),
    .A2(net333),
    .Y(_05440_),
    .B1(net401));
 sg13g2_nand2b_1 _22866_ (.Y(_05441_),
    .B(\cpu.intr.r_enable[3] ),
    .A_N(_05440_));
 sg13g2_nand4_1 _22867_ (.B(_05438_),
    .C(_05439_),
    .A(_05435_),
    .Y(_05442_),
    .D(_05441_));
 sg13g2_and2_1 _22868_ (.A(\cpu.uart.r_in[3] ),
    .B(_04883_),
    .X(_05443_));
 sg13g2_a221oi_1 _22869_ (.B2(\cpu.uart.r_div_value[11] ),
    .C1(_05443_),
    .B1(net399),
    .A1(\cpu.uart.r_div_value[3] ),
    .Y(_05444_),
    .A2(net363));
 sg13g2_o21ai_1 _22870_ (.B1(net1031),
    .Y(_05445_),
    .A1(net512),
    .A2(_05444_));
 sg13g2_a221oi_1 _22871_ (.B2(_04847_),
    .C1(_05445_),
    .B1(_05442_),
    .A1(_04901_),
    .Y(_05446_),
    .A2(_05432_));
 sg13g2_a22oi_1 _22872_ (.Y(_05447_),
    .B1(net414),
    .B2(\cpu.dcache.r_data[3][3] ),
    .A2(net372),
    .A1(\cpu.dcache.r_data[1][3] ));
 sg13g2_a22oi_1 _22873_ (.Y(_05448_),
    .B1(net532),
    .B2(\cpu.dcache.r_data[6][3] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][3] ));
 sg13g2_mux2_1 _22874_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(\cpu.dcache.r_data[7][3] ),
    .S(net552),
    .X(_05449_));
 sg13g2_a22oi_1 _22875_ (.Y(_05450_),
    .B1(_05449_),
    .B2(net620),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][3] ));
 sg13g2_nand2b_1 _22876_ (.Y(_05451_),
    .B(net537),
    .A_N(_05450_));
 sg13g2_nand3_1 _22877_ (.B(_05448_),
    .C(_05451_),
    .A(_05447_),
    .Y(_05452_));
 sg13g2_mux2_1 _22878_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(_05452_),
    .S(net332),
    .X(_05453_));
 sg13g2_nand2_1 _22879_ (.Y(_05454_),
    .A(\cpu.dcache.r_data[3][19] ),
    .B(net464));
 sg13g2_a22oi_1 _22880_ (.Y(_05455_),
    .B1(_09394_),
    .B2(\cpu.dcache.r_data[4][19] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][19] ));
 sg13g2_a22oi_1 _22881_ (.Y(_05456_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[7][19] ),
    .A2(net612),
    .A1(\cpu.dcache.r_data[6][19] ));
 sg13g2_a22oi_1 _22882_ (.Y(_05457_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net416),
    .A1(\cpu.dcache.r_data[1][19] ));
 sg13g2_nand4_1 _22883_ (.B(_05455_),
    .C(_05456_),
    .A(_05454_),
    .Y(_05458_),
    .D(_05457_));
 sg13g2_nor2_1 _22884_ (.A(net463),
    .B(_05458_),
    .Y(_05459_));
 sg13g2_a21oi_1 _22885_ (.A1(_00111_),
    .A2(net463),
    .Y(_05460_),
    .B1(_05459_));
 sg13g2_nand2_1 _22886_ (.Y(_05461_),
    .A(_11850_),
    .B(_05460_));
 sg13g2_nor2_1 _22887_ (.A(_11790_),
    .B(_05461_),
    .Y(_05462_));
 sg13g2_a21oi_1 _22888_ (.A1(net945),
    .A2(_05453_),
    .Y(_05463_),
    .B1(_05462_));
 sg13g2_a221oi_1 _22889_ (.B2(net991),
    .C1(net581),
    .B1(_05140_),
    .A1(_09813_),
    .Y(_05464_),
    .A2(_05133_));
 sg13g2_a21oi_1 _22890_ (.A1(net581),
    .A2(_05463_),
    .Y(_05465_),
    .B1(_05464_));
 sg13g2_nand2_1 _22891_ (.Y(_05466_),
    .A(net667),
    .B(_05453_));
 sg13g2_nand3_1 _22892_ (.B(_05461_),
    .C(_05466_),
    .A(net513),
    .Y(_05467_));
 sg13g2_o21ai_1 _22893_ (.B1(_05467_),
    .Y(_05468_),
    .A1(net460),
    .A2(_05465_));
 sg13g2_a22oi_1 _22894_ (.Y(_05469_),
    .B1(_05468_),
    .B2(net886),
    .A2(_05446_),
    .A1(_05419_));
 sg13g2_nand2_1 _22895_ (.Y(_05470_),
    .A(_03446_),
    .B(_05469_));
 sg13g2_o21ai_1 _22896_ (.B1(_05470_),
    .Y(_05471_),
    .A1(net780),
    .A2(net31));
 sg13g2_nand2_1 _22897_ (.Y(_05472_),
    .A(net151),
    .B(_05471_));
 sg13g2_o21ai_1 _22898_ (.B1(_05472_),
    .Y(_01040_),
    .A1(net127),
    .A2(_05412_));
 sg13g2_and2_1 _22899_ (.A(net710),
    .B(_04503_),
    .X(_05473_));
 sg13g2_a21oi_1 _22900_ (.A1(net635),
    .A2(_04539_),
    .Y(_05474_),
    .B1(_05473_));
 sg13g2_nor2_1 _22901_ (.A(_11348_),
    .B(_04214_),
    .Y(_05475_));
 sg13g2_o21ai_1 _22902_ (.B1(net1116),
    .Y(_05476_),
    .A1(net232),
    .A2(_05475_));
 sg13g2_o21ai_1 _22903_ (.B1(_05476_),
    .Y(_05477_),
    .A1(net232),
    .A2(_05474_));
 sg13g2_a22oi_1 _22904_ (.Y(_05478_),
    .B1(_05103_),
    .B2(\cpu.intr.r_timer_reload[4] ),
    .A2(_04859_),
    .A1(_09983_));
 sg13g2_a22oi_1 _22905_ (.Y(_05479_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[4] ),
    .A2(_04950_),
    .A1(\cpu.intr.r_timer_count[4] ));
 sg13g2_nand2_1 _22906_ (.Y(_05480_),
    .A(_05478_),
    .B(_05479_));
 sg13g2_nand2_1 _22907_ (.Y(_05481_),
    .A(net782),
    .B(net537));
 sg13g2_mux2_1 _22908_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(net496),
    .X(_05482_));
 sg13g2_a22oi_1 _22909_ (.Y(_05483_),
    .B1(_05482_),
    .B2(net551),
    .A2(net894),
    .A1(_09846_));
 sg13g2_buf_2 _22910_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05484_));
 sg13g2_a221oi_1 _22911_ (.B2(_09071_),
    .C1(_04875_),
    .B1(_04869_),
    .A1(_05484_),
    .Y(_05485_),
    .A2(_09961_));
 sg13g2_o21ai_1 _22912_ (.B1(_05485_),
    .Y(_05486_),
    .A1(_05481_),
    .A2(_05483_));
 sg13g2_nor2_1 _22913_ (.A(_05480_),
    .B(_05486_),
    .Y(_05487_));
 sg13g2_nand3_1 _22914_ (.B(net713),
    .C(_04851_),
    .A(net1036),
    .Y(_05488_));
 sg13g2_buf_2 _22915_ (.A(_05488_),
    .X(_05489_));
 sg13g2_a221oi_1 _22916_ (.B2(_05489_),
    .C1(_09821_),
    .B1(_05487_),
    .A1(_10185_),
    .Y(_05490_),
    .A2(net333));
 sg13g2_nor2_1 _22917_ (.A(_09060_),
    .B(_09070_),
    .Y(_05491_));
 sg13g2_o21ai_1 _22918_ (.B1(_05491_),
    .Y(_05492_),
    .A1(net333),
    .A2(_05487_));
 sg13g2_buf_2 _22919_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05493_));
 sg13g2_nand3_1 _22920_ (.B(_05493_),
    .C(net402),
    .A(net864),
    .Y(_05494_));
 sg13g2_nand3_1 _22921_ (.B(_10431_),
    .C(net363),
    .A(\cpu.gpio.r_enable_in[4] ),
    .Y(_05495_));
 sg13g2_buf_2 _22922_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05496_));
 sg13g2_nor3_1 _22923_ (.A(net898),
    .B(_04907_),
    .C(net597),
    .Y(_05497_));
 sg13g2_buf_2 _22924_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05498_));
 sg13g2_a22oi_1 _22925_ (.Y(_05499_),
    .B1(_05498_),
    .B2(net864),
    .A2(net837),
    .A1(_09052_));
 sg13g2_nor2b_1 _22926_ (.A(_05499_),
    .B_N(net461),
    .Y(_05500_));
 sg13g2_a221oi_1 _22927_ (.B2(net7),
    .C1(_05500_),
    .B1(_05497_),
    .A1(_05496_),
    .Y(_05501_),
    .A2(net397));
 sg13g2_nor2_1 _22928_ (.A(_09066_),
    .B(_04913_),
    .Y(_05502_));
 sg13g2_buf_2 _22929_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05503_));
 sg13g2_a22oi_1 _22930_ (.Y(_05504_),
    .B1(_04935_),
    .B2(_05503_),
    .A2(_04859_),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_nor2_1 _22931_ (.A(_04907_),
    .B(_05504_),
    .Y(_05505_));
 sg13g2_and3_1 _22932_ (.X(_05506_),
    .A(_09052_),
    .B(net944),
    .C(net402));
 sg13g2_o21ai_1 _22933_ (.B1(\cpu.gpio.r_enable_io[4] ),
    .Y(_05507_),
    .A1(_04961_),
    .A2(_05506_));
 sg13g2_nand3_1 _22934_ (.B(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .C(net429),
    .A(net837),
    .Y(_05508_));
 sg13g2_buf_2 _22935_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05509_));
 sg13g2_nand2_1 _22936_ (.Y(_05510_),
    .A(_05509_),
    .B(net398));
 sg13g2_buf_2 _22937_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05511_));
 sg13g2_a22oi_1 _22938_ (.Y(_05512_),
    .B1(_04942_),
    .B2(_05511_),
    .A2(_04930_),
    .A1(_09065_));
 sg13g2_nand4_1 _22939_ (.B(_05508_),
    .C(_05510_),
    .A(_05507_),
    .Y(_05513_),
    .D(_05512_));
 sg13g2_nor3_1 _22940_ (.A(_05502_),
    .B(_05505_),
    .C(_05513_),
    .Y(_05514_));
 sg13g2_nand4_1 _22941_ (.B(_05495_),
    .C(_05501_),
    .A(_05494_),
    .Y(_05515_),
    .D(_05514_));
 sg13g2_buf_1 _22942_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05516_));
 sg13g2_nor2_1 _22943_ (.A(_00126_),
    .B(_05016_),
    .Y(_05517_));
 sg13g2_a221oi_1 _22944_ (.B2(\cpu.spi.r_timeout[4] ),
    .C1(_05517_),
    .B1(_05014_),
    .A1(_05516_),
    .Y(_05518_),
    .A2(_04971_));
 sg13g2_o21ai_1 _22945_ (.B1(_05518_),
    .Y(_05519_),
    .A1(_00125_),
    .A2(_04968_));
 sg13g2_a21oi_1 _22946_ (.A1(_09168_),
    .A2(_04963_),
    .Y(_05520_),
    .B1(_05519_));
 sg13g2_nor2_1 _22947_ (.A(_09017_),
    .B(_05520_),
    .Y(_05521_));
 sg13g2_a221oi_1 _22948_ (.B2(_04901_),
    .C1(_05521_),
    .B1(_05515_),
    .A1(_05490_),
    .Y(_05522_),
    .A2(_05492_));
 sg13g2_a221oi_1 _22949_ (.B2(\cpu.uart.r_in[4] ),
    .C1(net512),
    .B1(_04883_),
    .A1(\cpu.uart.r_div_value[4] ),
    .Y(_05523_),
    .A2(net363));
 sg13g2_a21oi_1 _22950_ (.A1(net512),
    .A2(_05522_),
    .Y(_05524_),
    .B1(_05523_));
 sg13g2_nor3_1 _22951_ (.A(net580),
    .B(_04822_),
    .C(_05162_),
    .Y(_05525_));
 sg13g2_inv_1 _22952_ (.Y(_05526_),
    .A(_00121_));
 sg13g2_a22oi_1 _22953_ (.Y(_05527_),
    .B1(net372),
    .B2(\cpu.dcache.r_data[1][4] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][4] ));
 sg13g2_a22oi_1 _22954_ (.Y(_05528_),
    .B1(net475),
    .B2(\cpu.dcache.r_data[6][4] ),
    .A2(net414),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_mux2_1 _22955_ (.A0(\cpu.dcache.r_data[5][4] ),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(net552),
    .X(_05529_));
 sg13g2_a22oi_1 _22956_ (.Y(_05530_),
    .B1(_05529_),
    .B2(net620),
    .A2(net601),
    .A1(\cpu.dcache.r_data[4][4] ));
 sg13g2_nand2b_1 _22957_ (.Y(_05531_),
    .B(net537),
    .A_N(_05530_));
 sg13g2_nand4_1 _22958_ (.B(_05527_),
    .C(_05528_),
    .A(net332),
    .Y(_05532_),
    .D(_05531_));
 sg13g2_o21ai_1 _22959_ (.B1(_05532_),
    .Y(_05533_),
    .A1(_05526_),
    .A2(net332));
 sg13g2_nor2_1 _22960_ (.A(_05064_),
    .B(_05533_),
    .Y(_05534_));
 sg13g2_nand2_1 _22961_ (.Y(_05535_),
    .A(_05054_),
    .B(_05169_));
 sg13g2_a22oi_1 _22962_ (.Y(_05536_),
    .B1(net476),
    .B2(\cpu.dcache.r_data[5][20] ),
    .A2(net416),
    .A1(\cpu.dcache.r_data[1][20] ));
 sg13g2_a22oi_1 _22963_ (.Y(_05537_),
    .B1(net464),
    .B2(\cpu.dcache.r_data[3][20] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[2][20] ));
 sg13g2_mux2_1 _22964_ (.A0(\cpu.dcache.r_data[4][20] ),
    .A1(\cpu.dcache.r_data[6][20] ),
    .S(net514),
    .X(_05538_));
 sg13g2_a22oi_1 _22965_ (.Y(_05539_),
    .B1(_05538_),
    .B2(net713),
    .A2(net669),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_nand2b_1 _22966_ (.Y(_05540_),
    .B(net670),
    .A_N(_05539_));
 sg13g2_and4_1 _22967_ (.A(net403),
    .B(_05536_),
    .C(_05537_),
    .D(_05540_),
    .X(_05541_));
 sg13g2_a21oi_1 _22968_ (.A1(_00122_),
    .A2(net463),
    .Y(_05542_),
    .B1(_05541_));
 sg13g2_and2_1 _22969_ (.A(net668),
    .B(_05542_),
    .X(_05543_));
 sg13g2_nand2_1 _22970_ (.Y(_05544_),
    .A(net581),
    .B(_05543_));
 sg13g2_a21oi_1 _22971_ (.A1(_05535_),
    .A2(_05544_),
    .Y(_05545_),
    .B1(net945));
 sg13g2_nor4_1 _22972_ (.A(_04842_),
    .B(_05525_),
    .C(_05534_),
    .D(_05545_),
    .Y(_05546_));
 sg13g2_nor2_1 _22973_ (.A(net580),
    .B(_05533_),
    .Y(_05547_));
 sg13g2_nor4_1 _22974_ (.A(_08771_),
    .B(_04822_),
    .C(_05543_),
    .D(_05547_),
    .Y(_05548_));
 sg13g2_nor3_1 _22975_ (.A(net854),
    .B(_05546_),
    .C(_05548_),
    .Y(_05549_));
 sg13g2_a21oi_1 _22976_ (.A1(net854),
    .A2(_05524_),
    .Y(_05550_),
    .B1(_05549_));
 sg13g2_nor2_1 _22977_ (.A(net366),
    .B(net32),
    .Y(_05551_));
 sg13g2_a21oi_1 _22978_ (.A1(net31),
    .A2(_05550_),
    .Y(_05552_),
    .B1(_05551_));
 sg13g2_mux2_1 _22979_ (.A0(_05477_),
    .A1(_05552_),
    .S(net151),
    .X(_01041_));
 sg13g2_and2_1 _22980_ (.A(net710),
    .B(_04571_),
    .X(_05553_));
 sg13g2_a21oi_1 _22981_ (.A1(_05176_),
    .A2(_04568_),
    .Y(_05554_),
    .B1(_05553_));
 sg13g2_nand2_1 _22982_ (.Y(_05555_),
    .A(net947),
    .B(net232));
 sg13g2_o21ai_1 _22983_ (.B1(_05555_),
    .Y(_05556_),
    .A1(net232),
    .A2(_05554_));
 sg13g2_buf_1 _22984_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05557_));
 sg13g2_nor2_1 _22985_ (.A(_00133_),
    .B(net310),
    .Y(_05558_));
 sg13g2_a221oi_1 _22986_ (.B2(\cpu.spi.r_timeout[5] ),
    .C1(_05558_),
    .B1(_05014_),
    .A1(_05557_),
    .Y(_05559_),
    .A2(_04971_));
 sg13g2_o21ai_1 _22987_ (.B1(_05559_),
    .Y(_05560_),
    .A1(_00132_),
    .A2(_04968_));
 sg13g2_a21o_1 _22988_ (.A2(_04963_),
    .A1(_09167_),
    .B1(_05560_),
    .X(_05561_));
 sg13g2_and3_1 _22989_ (.X(_05562_),
    .A(_09056_),
    .B(_09057_),
    .C(_04854_));
 sg13g2_a221oi_1 _22990_ (.B2(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .C1(_05562_),
    .B1(_04859_),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .Y(_05563_),
    .A2(_09962_));
 sg13g2_o21ai_1 _22991_ (.B1(_05563_),
    .Y(_05564_),
    .A1(_00138_),
    .A2(_05421_));
 sg13g2_nand2b_1 _22992_ (.Y(_05565_),
    .B(net461),
    .A_N(_00135_));
 sg13g2_o21ai_1 _22993_ (.B1(_05565_),
    .Y(_05566_),
    .A1(_00137_),
    .A2(_05489_));
 sg13g2_a22oi_1 _22994_ (.Y(_05567_),
    .B1(_05566_),
    .B2(_11725_),
    .A2(_05497_),
    .A1(net8));
 sg13g2_inv_1 _22995_ (.Y(_05568_),
    .A(_00134_));
 sg13g2_a22oi_1 _22996_ (.Y(_05569_),
    .B1(_04930_),
    .B2(_09061_),
    .A2(net397),
    .A1(_05568_));
 sg13g2_nor2_1 _22997_ (.A(_00136_),
    .B(_05329_),
    .Y(_05570_));
 sg13g2_a221oi_1 _22998_ (.B2(_09056_),
    .C1(_05570_),
    .B1(_04961_),
    .A1(\cpu.gpio.r_enable_in[5] ),
    .Y(_05571_),
    .A2(_04923_));
 sg13g2_buf_2 _22999_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05572_));
 sg13g2_and2_1 _23000_ (.A(_09057_),
    .B(_04926_),
    .X(_05573_));
 sg13g2_a22oi_1 _23001_ (.Y(_05574_),
    .B1(_05573_),
    .B2(net461),
    .A2(net398),
    .A1(_05572_));
 sg13g2_nand4_1 _23002_ (.B(_05569_),
    .C(_05571_),
    .A(_05567_),
    .Y(_05575_),
    .D(_05574_));
 sg13g2_a21oi_1 _23003_ (.A1(net837),
    .A2(_05564_),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_o21ai_1 _23004_ (.B1(_05576_),
    .Y(_05577_),
    .A1(_09062_),
    .A2(_04913_));
 sg13g2_a22oi_1 _23005_ (.Y(_05578_),
    .B1(_04883_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net363),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_a22oi_1 _23006_ (.Y(_05579_),
    .B1(net474),
    .B2(\cpu.intr.r_timer_reload[21] ),
    .A2(net475),
    .A1(_09847_));
 sg13g2_a221oi_1 _23007_ (.B2(\cpu.intr.r_clock_cmp[5] ),
    .C1(net782),
    .B1(net413),
    .A1(_09987_),
    .Y(_05580_),
    .A2(net598));
 sg13g2_a21o_1 _23008_ (.A2(_05579_),
    .A1(net730),
    .B1(_05580_),
    .X(_05581_));
 sg13g2_nand2_1 _23009_ (.Y(_05582_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(_05103_));
 sg13g2_buf_1 _23010_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05583_));
 sg13g2_a22oi_1 _23011_ (.Y(_05584_),
    .B1(net402),
    .B2(_09038_),
    .A2(net429),
    .A1(_05583_));
 sg13g2_a22oi_1 _23012_ (.Y(_05585_),
    .B1(net396),
    .B2(\cpu.intr.r_clock_cmp[21] ),
    .A2(_04950_),
    .A1(\cpu.intr.r_timer_count[5] ));
 sg13g2_nand4_1 _23013_ (.B(_05582_),
    .C(_05584_),
    .A(_05581_),
    .Y(_05586_),
    .D(_05585_));
 sg13g2_a21oi_1 _23014_ (.A1(_09038_),
    .A2(net333),
    .Y(_05587_),
    .B1(net401));
 sg13g2_nor2b_1 _23015_ (.A(_05587_),
    .B_N(\cpu.intr.r_enable[5] ),
    .Y(_05588_));
 sg13g2_o21ai_1 _23016_ (.B1(_04847_),
    .Y(_05589_),
    .A1(_05586_),
    .A2(_05588_));
 sg13g2_o21ai_1 _23017_ (.B1(_05589_),
    .Y(_05590_),
    .A1(net512),
    .A2(_05578_));
 sg13g2_a221oi_1 _23018_ (.B2(_04901_),
    .C1(_05590_),
    .B1(_05577_),
    .A1(_04978_),
    .Y(_05591_),
    .A2(_05561_));
 sg13g2_nand2_1 _23019_ (.Y(_05592_),
    .A(\cpu.dcache.r_data[1][5] ),
    .B(net372));
 sg13g2_a22oi_1 _23020_ (.Y(_05593_),
    .B1(net598),
    .B2(\cpu.dcache.r_data[4][5] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_a22oi_1 _23021_ (.Y(_05594_),
    .B1(net474),
    .B2(\cpu.dcache.r_data[7][5] ),
    .A2(net532),
    .A1(\cpu.dcache.r_data[6][5] ));
 sg13g2_a22oi_1 _23022_ (.Y(_05595_),
    .B1(net476),
    .B2(\cpu.dcache.r_data[5][5] ),
    .A2(net477),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_nand4_1 _23023_ (.B(_05593_),
    .C(_05594_),
    .A(_05592_),
    .Y(_05596_),
    .D(_05595_));
 sg13g2_nand2_1 _23024_ (.Y(_05597_),
    .A(_00128_),
    .B(net463));
 sg13g2_o21ai_1 _23025_ (.B1(_05597_),
    .Y(_05598_),
    .A1(net459),
    .A2(_05596_));
 sg13g2_inv_1 _23026_ (.Y(_05599_),
    .A(_05598_));
 sg13g2_inv_1 _23027_ (.Y(_05600_),
    .A(_00129_));
 sg13g2_a22oi_1 _23028_ (.Y(_05601_),
    .B1(net364),
    .B2(\cpu.dcache.r_data[1][21] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][21] ));
 sg13g2_a22oi_1 _23029_ (.Y(_05602_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[7][21] ),
    .A2(net464),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_mux2_1 _23030_ (.A0(\cpu.dcache.r_data[4][21] ),
    .A1(\cpu.dcache.r_data[6][21] ),
    .S(net514),
    .X(_05603_));
 sg13g2_a22oi_1 _23031_ (.Y(_05604_),
    .B1(_05603_),
    .B2(net713),
    .A2(net773),
    .A1(\cpu.dcache.r_data[5][21] ));
 sg13g2_nand2b_1 _23032_ (.Y(_05605_),
    .B(net603),
    .A_N(_05604_));
 sg13g2_nand4_1 _23033_ (.B(_05601_),
    .C(_05602_),
    .A(net365),
    .Y(_05606_),
    .D(_05605_));
 sg13g2_o21ai_1 _23034_ (.B1(_05606_),
    .Y(_05607_),
    .A1(_05600_),
    .A2(net360));
 sg13g2_nor2_1 _23035_ (.A(_09812_),
    .B(_05607_),
    .Y(_05608_));
 sg13g2_a21oi_1 _23036_ (.A1(net667),
    .A2(_05599_),
    .Y(_05609_),
    .B1(_05608_));
 sg13g2_nor2_1 _23037_ (.A(net636),
    .B(_05201_),
    .Y(_05610_));
 sg13g2_a21oi_1 _23038_ (.A1(net636),
    .A2(_05608_),
    .Y(_05611_),
    .B1(_05610_));
 sg13g2_nor3_1 _23039_ (.A(_11850_),
    .B(net636),
    .C(_05193_),
    .Y(_05612_));
 sg13g2_a21oi_1 _23040_ (.A1(_05065_),
    .A2(_05599_),
    .Y(_05613_),
    .B1(_05612_));
 sg13g2_o21ai_1 _23041_ (.B1(_05613_),
    .Y(_05614_),
    .A1(net945),
    .A2(_05611_));
 sg13g2_nor2_1 _23042_ (.A(net513),
    .B(_05614_),
    .Y(_05615_));
 sg13g2_a21oi_1 _23043_ (.A1(net513),
    .A2(_05609_),
    .Y(_05616_),
    .B1(_05615_));
 sg13g2_nor2_1 _23044_ (.A(net854),
    .B(_05616_),
    .Y(_05617_));
 sg13g2_a21oi_1 _23045_ (.A1(net854),
    .A2(_05591_),
    .Y(_05618_),
    .B1(_05617_));
 sg13g2_nand2_1 _23046_ (.Y(_05619_),
    .A(net32),
    .B(_05618_));
 sg13g2_o21ai_1 _23047_ (.B1(_05619_),
    .Y(_05620_),
    .A1(net865),
    .A2(net31));
 sg13g2_mux2_1 _23048_ (.A0(_05556_),
    .A1(_05620_),
    .S(net151),
    .X(_01042_));
 sg13g2_and2_1 _23049_ (.A(net710),
    .B(_04604_),
    .X(_05621_));
 sg13g2_nor3_1 _23050_ (.A(net711),
    .B(_04574_),
    .C(_04601_),
    .Y(_05622_));
 sg13g2_nor3_1 _23051_ (.A(net232),
    .B(_05621_),
    .C(_05622_),
    .Y(_05623_));
 sg13g2_o21ai_1 _23052_ (.B1(_11357_),
    .Y(_05624_),
    .A1(_08669_),
    .A2(net231));
 sg13g2_nand2_1 _23053_ (.Y(_05625_),
    .A(\cpu.dcache.r_data[3][6] ),
    .B(net477));
 sg13g2_a22oi_1 _23054_ (.Y(_05626_),
    .B1(net598),
    .B2(\cpu.dcache.r_data[4][6] ),
    .A2(net395),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_a22oi_1 _23055_ (.Y(_05627_),
    .B1(net531),
    .B2(\cpu.dcache.r_data[7][6] ),
    .A2(net532),
    .A1(\cpu.dcache.r_data[6][6] ));
 sg13g2_a22oi_1 _23056_ (.Y(_05628_),
    .B1(net476),
    .B2(\cpu.dcache.r_data[5][6] ),
    .A2(net364),
    .A1(\cpu.dcache.r_data[1][6] ));
 sg13g2_nand4_1 _23057_ (.B(_05626_),
    .C(_05627_),
    .A(_05625_),
    .Y(_05629_),
    .D(_05628_));
 sg13g2_nand2_1 _23058_ (.Y(_05630_),
    .A(_00140_),
    .B(net463));
 sg13g2_o21ai_1 _23059_ (.B1(_05630_),
    .Y(_05631_),
    .A1(net459),
    .A2(_05629_));
 sg13g2_buf_1 _23060_ (.A(_05631_),
    .X(_05632_));
 sg13g2_a22oi_1 _23061_ (.Y(_05633_),
    .B1(_05632_),
    .B2(net581),
    .A2(_05226_),
    .A1(_05044_));
 sg13g2_nor2b_1 _23062_ (.A(_05233_),
    .B_N(_05044_),
    .Y(_05634_));
 sg13g2_a22oi_1 _23063_ (.Y(_05635_),
    .B1(net372),
    .B2(\cpu.dcache.r_data[1][22] ),
    .A2(net415),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_a22oi_1 _23064_ (.Y(_05636_),
    .B1(_02906_),
    .B2(\cpu.dcache.r_data[7][22] ),
    .A2(net414),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_mux2_1 _23065_ (.A0(\cpu.dcache.r_data[4][22] ),
    .A1(\cpu.dcache.r_data[6][22] ),
    .S(net552),
    .X(_05637_));
 sg13g2_a22oi_1 _23066_ (.Y(_05638_),
    .B1(_05637_),
    .B2(net638),
    .A2(net773),
    .A1(\cpu.dcache.r_data[5][22] ));
 sg13g2_nand2b_1 _23067_ (.Y(_05639_),
    .B(net537),
    .A_N(_05638_));
 sg13g2_and4_1 _23068_ (.A(net332),
    .B(_05635_),
    .C(_05636_),
    .D(_05639_),
    .X(_05640_));
 sg13g2_a21oi_1 _23069_ (.A1(_00141_),
    .A2(net459),
    .Y(_05641_),
    .B1(_05640_));
 sg13g2_o21ai_1 _23070_ (.B1(_05043_),
    .Y(_05642_),
    .A1(_09942_),
    .A2(_05632_));
 sg13g2_nor2_1 _23071_ (.A(_05064_),
    .B(_05632_),
    .Y(_05643_));
 sg13g2_a221oi_1 _23072_ (.B2(_05054_),
    .C1(_05643_),
    .B1(_05642_),
    .A1(_09942_),
    .Y(_05644_),
    .A2(_05641_));
 sg13g2_a21oi_1 _23073_ (.A1(_05226_),
    .A2(_05634_),
    .Y(_05645_),
    .B1(_05644_));
 sg13g2_o21ai_1 _23074_ (.B1(_05645_),
    .Y(_05646_),
    .A1(net991),
    .A2(_05633_));
 sg13g2_buf_1 _23075_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05647_));
 sg13g2_nor2_1 _23076_ (.A(_00145_),
    .B(_05016_),
    .Y(_05648_));
 sg13g2_a221oi_1 _23077_ (.B2(\cpu.spi.r_timeout[6] ),
    .C1(_05648_),
    .B1(_05014_),
    .A1(_05647_),
    .Y(_05649_),
    .A2(_04971_));
 sg13g2_o21ai_1 _23078_ (.B1(_05649_),
    .Y(_05650_),
    .A1(_00144_),
    .A2(_04968_));
 sg13g2_a21o_1 _23079_ (.A2(_04963_),
    .A1(_09161_),
    .B1(_05650_),
    .X(_05651_));
 sg13g2_a22oi_1 _23080_ (.Y(_05652_),
    .B1(net461),
    .B2(_09047_),
    .A2(_09961_),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_o21ai_1 _23081_ (.B1(_05652_),
    .Y(_05653_),
    .A1(_00150_),
    .A2(_05421_));
 sg13g2_a21o_1 _23082_ (.A2(_04859_),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B1(_05653_),
    .X(_05654_));
 sg13g2_and3_1 _23083_ (.X(_05655_),
    .A(_09047_),
    .B(_04926_),
    .C(_04854_));
 sg13g2_o21ai_1 _23084_ (.B1(\cpu.gpio.r_enable_io[6] ),
    .Y(_05656_),
    .A1(_04961_),
    .A2(_05655_));
 sg13g2_nand2b_1 _23085_ (.Y(_05657_),
    .B(_04887_),
    .A_N(_00147_));
 sg13g2_o21ai_1 _23086_ (.B1(_05657_),
    .Y(_05658_),
    .A1(_00149_),
    .A2(_05489_));
 sg13g2_nor2b_1 _23087_ (.A(net995),
    .B_N(\cpu.gpio.r_enable_in[6] ),
    .Y(_05659_));
 sg13g2_a22oi_1 _23088_ (.Y(_05660_),
    .B1(_05659_),
    .B2(net400),
    .A2(_05658_),
    .A1(net864));
 sg13g2_buf_1 _23089_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05661_));
 sg13g2_nand2b_1 _23090_ (.Y(_05662_),
    .B(net397),
    .A_N(_00146_));
 sg13g2_o21ai_1 _23091_ (.B1(_05662_),
    .Y(_05663_),
    .A1(_00148_),
    .A2(_05329_));
 sg13g2_a221oi_1 _23092_ (.B2(_09067_),
    .C1(_05663_),
    .B1(_04930_),
    .A1(_05661_),
    .Y(_05664_),
    .A2(net398));
 sg13g2_nand2_1 _23093_ (.Y(_05665_),
    .A(net9),
    .B(_05497_));
 sg13g2_nand4_1 _23094_ (.B(_05660_),
    .C(_05664_),
    .A(_05656_),
    .Y(_05666_),
    .D(_05665_));
 sg13g2_a21oi_1 _23095_ (.A1(net837),
    .A2(_05654_),
    .Y(_05667_),
    .B1(_05666_));
 sg13g2_o21ai_1 _23096_ (.B1(_05667_),
    .Y(_05668_),
    .A1(_09068_),
    .A2(_04913_));
 sg13g2_a22oi_1 _23097_ (.Y(_05669_),
    .B1(_04883_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net363),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_a22oi_1 _23098_ (.Y(_05670_),
    .B1(net474),
    .B2(\cpu.intr.r_timer_reload[22] ),
    .A2(net475),
    .A1(_09848_));
 sg13g2_a221oi_1 _23099_ (.B2(\cpu.intr.r_clock_cmp[6] ),
    .C1(net782),
    .B1(net413),
    .A1(_09991_),
    .Y(_05671_),
    .A2(net598));
 sg13g2_a21oi_1 _23100_ (.A1(net730),
    .A2(_05670_),
    .Y(_05672_),
    .B1(_05671_));
 sg13g2_buf_2 _23101_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05673_));
 sg13g2_a22oi_1 _23102_ (.Y(_05674_),
    .B1(_04950_),
    .B2(\cpu.intr.r_timer_count[6] ),
    .A2(net429),
    .A1(_05673_));
 sg13g2_a22oi_1 _23103_ (.Y(_05675_),
    .B1(_05103_),
    .B2(\cpu.intr.r_timer_reload[6] ),
    .A2(_04935_),
    .A1(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_nand2_1 _23104_ (.Y(_05676_),
    .A(_05674_),
    .B(_05675_));
 sg13g2_o21ai_1 _23105_ (.B1(_05021_),
    .Y(_05677_),
    .A1(_05672_),
    .A2(_05676_));
 sg13g2_o21ai_1 _23106_ (.B1(_05677_),
    .Y(_05678_),
    .A1(net512),
    .A2(_05669_));
 sg13g2_a221oi_1 _23107_ (.B2(_04901_),
    .C1(_05678_),
    .B1(_05668_),
    .A1(_04978_),
    .Y(_05679_),
    .A2(_05651_));
 sg13g2_nand2b_1 _23108_ (.Y(_05680_),
    .B(net854),
    .A_N(_05679_));
 sg13g2_o21ai_1 _23109_ (.B1(_05680_),
    .Y(_05681_),
    .A1(_02878_),
    .A2(_05646_));
 sg13g2_mux2_1 _23110_ (.A0(_02914_),
    .A1(_05681_),
    .S(_04797_),
    .X(_05682_));
 sg13g2_nand2_1 _23111_ (.Y(_05683_),
    .A(_05413_),
    .B(_05682_));
 sg13g2_o21ai_1 _23112_ (.B1(_05683_),
    .Y(_01043_),
    .A1(_05623_),
    .A2(_05624_));
 sg13g2_nand2_1 _23113_ (.Y(_05684_),
    .A(net32),
    .B(_05078_));
 sg13g2_o21ai_1 _23114_ (.B1(_05684_),
    .Y(_05685_),
    .A1(net1037),
    .A2(net31));
 sg13g2_nand2_1 _23115_ (.Y(_05686_),
    .A(net635),
    .B(_04629_));
 sg13g2_o21ai_1 _23116_ (.B1(_05686_),
    .Y(_05687_),
    .A1(net635),
    .A2(_04630_));
 sg13g2_nor3_1 _23117_ (.A(\cpu.ex.pc[7] ),
    .B(net231),
    .C(net153),
    .Y(_05688_));
 sg13g2_a221oi_1 _23118_ (.B2(_04989_),
    .C1(_05688_),
    .B1(_05687_),
    .A1(net128),
    .Y(_01044_),
    .A2(_05685_));
 sg13g2_mux2_1 _23119_ (.A0(_04831_),
    .A1(_04838_),
    .S(_05098_),
    .X(_05689_));
 sg13g2_a22oi_1 _23120_ (.Y(_05690_),
    .B1(net458),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(net361),
    .A1(\cpu.intr.r_timer_reload[8] ));
 sg13g2_a22oi_1 _23121_ (.Y(_05691_),
    .B1(net362),
    .B2(\cpu.intr.r_timer_count[8] ),
    .A2(net462),
    .A1(_10003_));
 sg13g2_buf_2 _23122_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05692_));
 sg13g2_a22oi_1 _23123_ (.Y(_05693_),
    .B1(net396),
    .B2(\cpu.intr.r_clock_cmp[24] ),
    .A2(net375),
    .A1(_05692_));
 sg13g2_nand3_1 _23124_ (.B(_05691_),
    .C(_05693_),
    .A(_05690_),
    .Y(_05694_));
 sg13g2_a221oi_1 _23125_ (.B2(_05101_),
    .C1(net943),
    .B1(_05694_),
    .A1(_05081_),
    .Y(_05695_),
    .A2(_05689_));
 sg13g2_nor2_1 _23126_ (.A(_05080_),
    .B(_05695_),
    .Y(_05696_));
 sg13g2_mux2_1 _23127_ (.A0(_09012_),
    .A1(_05696_),
    .S(net32),
    .X(_05697_));
 sg13g2_nand2_1 _23128_ (.Y(_05698_),
    .A(_05176_),
    .B(_04658_));
 sg13g2_a21oi_1 _23129_ (.A1(net710),
    .A2(_04660_),
    .Y(_05699_),
    .B1(_04988_));
 sg13g2_a221oi_1 _23130_ (.B2(_05699_),
    .C1(net153),
    .B1(_05698_),
    .A1(net948),
    .Y(_05700_),
    .A2(net232));
 sg13g2_a21o_1 _23131_ (.A2(_05697_),
    .A1(_05117_),
    .B1(_05700_),
    .X(_01045_));
 sg13g2_a22oi_1 _23132_ (.Y(_05701_),
    .B1(net361),
    .B2(\cpu.intr.r_timer_reload[9] ),
    .A2(net362),
    .A1(\cpu.intr.r_timer_count[9] ));
 sg13g2_buf_2 _23133_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05702_));
 sg13g2_mux2_1 _23134_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(\cpu.intr.r_clock_cmp[25] ),
    .S(net668),
    .X(_05703_));
 sg13g2_a22oi_1 _23135_ (.Y(_05704_),
    .B1(_05703_),
    .B2(net413),
    .A2(_09963_),
    .A1(_05702_));
 sg13g2_nand2_1 _23136_ (.Y(_05705_),
    .A(_10010_),
    .B(_04860_));
 sg13g2_nand3_1 _23137_ (.B(_05704_),
    .C(_05705_),
    .A(_05701_),
    .Y(_05706_));
 sg13g2_a21o_1 _23138_ (.A2(_05280_),
    .A1(net609),
    .B1(_05289_),
    .X(_05707_));
 sg13g2_a221oi_1 _23139_ (.B2(_05081_),
    .C1(net943),
    .B1(_05707_),
    .A1(_05101_),
    .Y(_05708_),
    .A2(_05706_));
 sg13g2_o21ai_1 _23140_ (.B1(_04797_),
    .Y(_05709_),
    .A1(_05080_),
    .A2(_05708_));
 sg13g2_o21ai_1 _23141_ (.B1(_05709_),
    .Y(_05710_),
    .A1(_10627_),
    .A2(_04992_));
 sg13g2_nand2_1 _23142_ (.Y(_05711_),
    .A(net635),
    .B(_04692_));
 sg13g2_a21oi_1 _23143_ (.A1(net711),
    .A2(_04662_),
    .Y(_05712_),
    .B1(_04793_));
 sg13g2_nor3_1 _23144_ (.A(_08719_),
    .B(net231),
    .C(_04983_),
    .Y(_05713_));
 sg13g2_a221oi_1 _23145_ (.B2(_05712_),
    .C1(_05713_),
    .B1(_05711_),
    .A1(net151),
    .Y(_01046_),
    .A2(_05710_));
 sg13g2_nand2b_1 _23146_ (.Y(_05714_),
    .B(\cpu.dec.r_rd[0] ),
    .A_N(_03337_));
 sg13g2_a21oi_1 _23147_ (.A1(net231),
    .A2(_05714_),
    .Y(_05715_),
    .B1(net153));
 sg13g2_a21o_1 _23148_ (.A2(_05117_),
    .A1(net1010),
    .B1(_05715_),
    .X(_01047_));
 sg13g2_nor2b_1 _23149_ (.A(_03337_),
    .B_N(\cpu.dec.r_rd[1] ),
    .Y(_05716_));
 sg13g2_o21ai_1 _23150_ (.B1(net152),
    .Y(_05717_),
    .A1(net232),
    .A2(_05716_));
 sg13g2_o21ai_1 _23151_ (.B1(_05717_),
    .Y(_01048_),
    .A1(_03410_),
    .A2(net152));
 sg13g2_nor3_1 _23152_ (.A(_03337_),
    .B(_09181_),
    .C(_10183_),
    .Y(_05718_));
 sg13g2_nand3_1 _23153_ (.B(net152),
    .C(_05718_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05719_));
 sg13g2_o21ai_1 _23154_ (.B1(_05719_),
    .Y(_01049_),
    .A1(_10058_),
    .A2(_05252_));
 sg13g2_inv_1 _23155_ (.Y(_05720_),
    .A(_10056_));
 sg13g2_nand3_1 _23156_ (.B(_11357_),
    .C(_05718_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05721_));
 sg13g2_o21ai_1 _23157_ (.B1(_05721_),
    .Y(_01050_),
    .A1(_05720_),
    .A2(_05252_));
 sg13g2_mux2_1 _23158_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_05413_),
    .X(_01051_));
 sg13g2_nor2_1 _23159_ (.A(_10937_),
    .B(_10942_),
    .Y(_05722_));
 sg13g2_nand2_1 _23160_ (.Y(_05723_),
    .A(net718),
    .B(net425));
 sg13g2_o21ai_1 _23161_ (.B1(_05723_),
    .Y(_05724_),
    .A1(_10815_),
    .A2(_05722_));
 sg13g2_mux2_1 _23162_ (.A0(net884),
    .A1(_05724_),
    .S(net152),
    .X(_01052_));
 sg13g2_a22oi_1 _23163_ (.Y(_05725_),
    .B1(net490),
    .B2(_11114_),
    .A2(net425),
    .A1(net1089));
 sg13g2_nand2_1 _23164_ (.Y(_05726_),
    .A(net551),
    .B(net425));
 sg13g2_o21ai_1 _23165_ (.B1(_05726_),
    .Y(_05727_),
    .A1(_10815_),
    .A2(_10844_));
 sg13g2_nor2_1 _23166_ (.A(net1033),
    .B(_05727_),
    .Y(_05728_));
 sg13g2_a21o_1 _23167_ (.A2(_05725_),
    .A1(net1033),
    .B1(_05728_),
    .X(_05729_));
 sg13g2_nand2_1 _23168_ (.Y(_05730_),
    .A(_10018_),
    .B(net151));
 sg13g2_o21ai_1 _23169_ (.B1(_05730_),
    .Y(_01053_),
    .A1(net127),
    .A2(_05729_));
 sg13g2_buf_1 _23170_ (.A(net943),
    .X(_05731_));
 sg13g2_nand2_1 _23171_ (.Y(_05732_),
    .A(_10869_),
    .B(_10878_));
 sg13g2_a22oi_1 _23172_ (.Y(_05733_),
    .B1(net490),
    .B2(_05732_),
    .A2(net425),
    .A1(_09094_));
 sg13g2_a221oi_1 _23173_ (.B2(_10156_),
    .C1(net836),
    .B1(net490),
    .A1(net1094),
    .Y(_05734_),
    .A2(net425));
 sg13g2_a21oi_1 _23174_ (.A1(net836),
    .A2(_05733_),
    .Y(_05735_),
    .B1(_05734_));
 sg13g2_mux2_1 _23175_ (.A0(_10025_),
    .A1(_05735_),
    .S(net152),
    .X(_01054_));
 sg13g2_a22oi_1 _23176_ (.Y(_05736_),
    .B1(_11049_),
    .B2(_10802_),
    .A2(_11182_),
    .A1(net366));
 sg13g2_nor3_1 _23177_ (.A(net836),
    .B(_11167_),
    .C(_11168_),
    .Y(_05737_));
 sg13g2_a21o_1 _23178_ (.A2(_05736_),
    .A1(_05731_),
    .B1(_05737_),
    .X(_05738_));
 sg13g2_nand2_1 _23179_ (.Y(_05739_),
    .A(_10030_),
    .B(net151));
 sg13g2_o21ai_1 _23180_ (.B1(_05739_),
    .Y(_01055_),
    .A1(net127),
    .A2(_05738_));
 sg13g2_mux2_1 _23181_ (.A0(_11259_),
    .A1(_10758_),
    .S(net836),
    .X(_05740_));
 sg13g2_nand2_1 _23182_ (.Y(_05741_),
    .A(_10036_),
    .B(net151));
 sg13g2_o21ai_1 _23183_ (.B1(_05741_),
    .Y(_01056_),
    .A1(_05340_),
    .A2(_05740_));
 sg13g2_mux2_1 _23184_ (.A0(_11234_),
    .A1(_10995_),
    .S(net836),
    .X(_05742_));
 sg13g2_nand2_1 _23185_ (.Y(_05743_),
    .A(_10043_),
    .B(net151));
 sg13g2_o21ai_1 _23186_ (.B1(_05743_),
    .Y(_01057_),
    .A1(_05340_),
    .A2(_05742_));
 sg13g2_mux2_1 _23187_ (.A0(_11200_),
    .A1(_10971_),
    .S(net836),
    .X(_05744_));
 sg13g2_nand2_1 _23188_ (.Y(_05745_),
    .A(_10048_),
    .B(_04796_));
 sg13g2_o21ai_1 _23189_ (.B1(_05745_),
    .Y(_01058_),
    .A1(net128),
    .A2(_05744_));
 sg13g2_nand2_1 _23190_ (.Y(_05746_),
    .A(_10895_),
    .B(_10913_));
 sg13g2_a22oi_1 _23191_ (.Y(_05747_),
    .B1(net490),
    .B2(_05746_),
    .A2(net425),
    .A1(_09943_));
 sg13g2_nand2_1 _23192_ (.Y(_05748_),
    .A(_02808_),
    .B(net154));
 sg13g2_o21ai_1 _23193_ (.B1(_05748_),
    .Y(_01059_),
    .A1(net128),
    .A2(_05747_));
 sg13g2_mux2_1 _23194_ (.A0(net862),
    .A1(_05727_),
    .S(net152),
    .X(_01060_));
 sg13g2_nand2_1 _23195_ (.Y(_05749_),
    .A(net964),
    .B(net154));
 sg13g2_o21ai_1 _23196_ (.B1(_05749_),
    .Y(_01061_),
    .A1(net128),
    .A2(_05733_));
 sg13g2_nand2_1 _23197_ (.Y(_05750_),
    .A(net1016),
    .B(net154));
 sg13g2_o21ai_1 _23198_ (.B1(_05750_),
    .Y(_01062_),
    .A1(_05736_),
    .A2(net127));
 sg13g2_nand2_1 _23199_ (.Y(_05751_),
    .A(net1015),
    .B(net154));
 sg13g2_o21ai_1 _23200_ (.B1(_05751_),
    .Y(_01063_),
    .A1(_10758_),
    .A2(net127));
 sg13g2_nand2_1 _23201_ (.Y(_05752_),
    .A(_09934_),
    .B(net154));
 sg13g2_o21ai_1 _23202_ (.B1(_05752_),
    .Y(_01064_),
    .A1(_10995_),
    .A2(net127));
 sg13g2_nand2_1 _23203_ (.Y(_05753_),
    .A(net1012),
    .B(net154));
 sg13g2_o21ai_1 _23204_ (.B1(_05753_),
    .Y(_01065_),
    .A1(_10971_),
    .A2(net127));
 sg13g2_a22oi_1 _23205_ (.Y(_05754_),
    .B1(net490),
    .B2(_11089_),
    .A2(net425),
    .A1(net1038));
 sg13g2_nor2_1 _23206_ (.A(_05731_),
    .B(_05754_),
    .Y(_05755_));
 sg13g2_a21oi_1 _23207_ (.A1(net836),
    .A2(_05724_),
    .Y(_05756_),
    .B1(_05755_));
 sg13g2_nand2_1 _23208_ (.Y(_05757_),
    .A(_10008_),
    .B(net154));
 sg13g2_o21ai_1 _23209_ (.B1(_05757_),
    .Y(_01066_),
    .A1(net128),
    .A2(_05756_));
 sg13g2_mux2_1 _23210_ (.A0(_11070_),
    .A1(_05747_),
    .S(net836),
    .X(_05758_));
 sg13g2_nand2_1 _23211_ (.Y(_05759_),
    .A(_10013_),
    .B(net154));
 sg13g2_o21ai_1 _23212_ (.B1(_05759_),
    .Y(_01067_),
    .A1(net128),
    .A2(_05758_));
 sg13g2_nand2_1 _23213_ (.Y(_05760_),
    .A(_08363_),
    .B(net497));
 sg13g2_o21ai_1 _23214_ (.B1(_05760_),
    .Y(_05761_),
    .A1(_08822_),
    .A2(net497));
 sg13g2_or3_1 _23215_ (.A(_10921_),
    .B(_10811_),
    .C(_10852_),
    .X(_05762_));
 sg13g2_o21ai_1 _23216_ (.B1(_03219_),
    .Y(_05763_),
    .A1(_10888_),
    .A2(_05762_));
 sg13g2_buf_1 _23217_ (.A(_05763_),
    .X(_05764_));
 sg13g2_nor4_1 _23218_ (.A(_08737_),
    .B(_04724_),
    .C(_03752_),
    .D(_03411_),
    .Y(_05765_));
 sg13g2_buf_1 _23219_ (.A(_05765_),
    .X(_05766_));
 sg13g2_buf_1 _23220_ (.A(_00288_),
    .X(_05767_));
 sg13g2_nand2b_1 _23221_ (.Y(_05768_),
    .B(net841),
    .A_N(net1068));
 sg13g2_o21ai_1 _23222_ (.B1(_05768_),
    .Y(_05769_),
    .A1(net841),
    .A2(net675));
 sg13g2_nand4_1 _23223_ (.B(_05764_),
    .C(net579),
    .A(net347),
    .Y(_05770_),
    .D(_05769_));
 sg13g2_o21ai_1 _23224_ (.B1(_05770_),
    .Y(_05771_),
    .A1(net347),
    .A2(_05761_));
 sg13g2_buf_1 _23225_ (.A(_10525_),
    .X(_05772_));
 sg13g2_buf_1 _23226_ (.A(_05772_),
    .X(_05773_));
 sg13g2_nand2_1 _23227_ (.Y(_05774_),
    .A(_05764_),
    .B(net579));
 sg13g2_a21oi_2 _23228_ (.B1(_09182_),
    .Y(_05775_),
    .A2(_05774_),
    .A1(net347));
 sg13g2_nor2_1 _23229_ (.A(_05773_),
    .B(_05775_),
    .Y(_05776_));
 sg13g2_a21oi_1 _23230_ (.A1(_09129_),
    .A2(_05771_),
    .Y(_01070_),
    .B1(_05776_));
 sg13g2_buf_1 _23231_ (.A(_10594_),
    .X(_05777_));
 sg13g2_nand2b_1 _23232_ (.Y(_05778_),
    .B(net941),
    .A_N(net942));
 sg13g2_buf_1 _23233_ (.A(_05778_),
    .X(_05779_));
 sg13g2_nand2b_1 _23234_ (.Y(_05780_),
    .B(net942),
    .A_N(_10594_));
 sg13g2_buf_1 _23235_ (.A(_05780_),
    .X(_05781_));
 sg13g2_nand3_1 _23236_ (.B(net709),
    .C(_05781_),
    .A(net841),
    .Y(_05782_));
 sg13g2_o21ai_1 _23237_ (.B1(_05782_),
    .Y(_05783_),
    .A1(net841),
    .A2(net611));
 sg13g2_nand3_1 _23238_ (.B(net579),
    .C(_05783_),
    .A(_05764_),
    .Y(_05784_));
 sg13g2_nor2_1 _23239_ (.A(net611),
    .B(net497),
    .Y(_05785_));
 sg13g2_a21oi_1 _23240_ (.A1(_08423_),
    .A2(net497),
    .Y(_05786_),
    .B1(_05785_));
 sg13g2_mux2_1 _23241_ (.A0(_05784_),
    .A1(_05786_),
    .S(net311),
    .X(_05787_));
 sg13g2_nor2_1 _23242_ (.A(net679),
    .B(_05787_),
    .Y(_05788_));
 sg13g2_nor2_1 _23243_ (.A(net941),
    .B(_05775_),
    .Y(_05789_));
 sg13g2_nor2_1 _23244_ (.A(_05788_),
    .B(_05789_),
    .Y(_01071_));
 sg13g2_nand2_1 _23245_ (.Y(_05790_),
    .A(_10525_),
    .B(_10594_));
 sg13g2_buf_2 _23246_ (.A(_05790_),
    .X(_05791_));
 sg13g2_inv_2 _23247_ (.Y(_05792_),
    .A(_10566_));
 sg13g2_nand2b_1 _23248_ (.Y(_05793_),
    .B(_05792_),
    .A_N(_05791_));
 sg13g2_buf_1 _23249_ (.A(_10566_),
    .X(_05794_));
 sg13g2_nand2_1 _23250_ (.Y(_05795_),
    .A(net940),
    .B(_05791_));
 sg13g2_nand3_1 _23251_ (.B(_05793_),
    .C(_05795_),
    .A(net841),
    .Y(_05796_));
 sg13g2_o21ai_1 _23252_ (.B1(_05796_),
    .Y(_05797_),
    .A1(_03377_),
    .A2(net672));
 sg13g2_nand3_1 _23253_ (.B(net579),
    .C(_05797_),
    .A(_05764_),
    .Y(_05798_));
 sg13g2_nor2_1 _23254_ (.A(net672),
    .B(net497),
    .Y(_05799_));
 sg13g2_a21oi_1 _23255_ (.A1(_08599_),
    .A2(net497),
    .Y(_05800_),
    .B1(_05799_));
 sg13g2_mux2_1 _23256_ (.A0(_05798_),
    .A1(_05800_),
    .S(net311),
    .X(_05801_));
 sg13g2_nor2_1 _23257_ (.A(net679),
    .B(_05801_),
    .Y(_05802_));
 sg13g2_nor2_1 _23258_ (.A(net940),
    .B(_05775_),
    .Y(_05803_));
 sg13g2_nor2_1 _23259_ (.A(_05802_),
    .B(_05803_),
    .Y(_01072_));
 sg13g2_nor2_1 _23260_ (.A(net890),
    .B(net497),
    .Y(_05804_));
 sg13g2_a21oi_1 _23261_ (.A1(_08382_),
    .A2(net497),
    .Y(_05805_),
    .B1(_05804_));
 sg13g2_buf_1 _23262_ (.A(_10614_),
    .X(_05806_));
 sg13g2_buf_1 _23263_ (.A(net939),
    .X(_05807_));
 sg13g2_nor2_2 _23264_ (.A(_05792_),
    .B(_05791_),
    .Y(_05808_));
 sg13g2_xnor2_1 _23265_ (.Y(_05809_),
    .A(net834),
    .B(_05808_));
 sg13g2_nand2_1 _23266_ (.Y(_05810_),
    .A(net841),
    .B(_05809_));
 sg13g2_o21ai_1 _23267_ (.B1(_05810_),
    .Y(_05811_),
    .A1(net841),
    .A2(net890));
 sg13g2_nand4_1 _23268_ (.B(_05764_),
    .C(net579),
    .A(net347),
    .Y(_05812_),
    .D(_05811_));
 sg13g2_o21ai_1 _23269_ (.B1(_05812_),
    .Y(_05813_),
    .A1(net347),
    .A2(_05805_));
 sg13g2_nor2_1 _23270_ (.A(_05807_),
    .B(_05775_),
    .Y(_05814_));
 sg13g2_a21oi_1 _23271_ (.A1(_09129_),
    .A2(_05813_),
    .Y(_01073_),
    .B1(_05814_));
 sg13g2_buf_2 _23272_ (.A(_00188_),
    .X(_05815_));
 sg13g2_buf_1 _23273_ (.A(net1090),
    .X(_05816_));
 sg13g2_nor2_2 _23274_ (.A(net938),
    .B(net834),
    .Y(_05817_));
 sg13g2_nand2_1 _23275_ (.Y(_05818_),
    .A(_05815_),
    .B(_05817_));
 sg13g2_nand3b_1 _23276_ (.B(net579),
    .C(_09098_),
    .Y(_05819_),
    .A_N(_10242_));
 sg13g2_buf_1 _23277_ (.A(_05819_),
    .X(_05820_));
 sg13g2_or3_1 _23278_ (.A(net835),
    .B(_05777_),
    .C(_05820_),
    .X(_05821_));
 sg13g2_buf_1 _23279_ (.A(_05821_),
    .X(_05822_));
 sg13g2_nor2_1 _23280_ (.A(_05818_),
    .B(_05822_),
    .Y(_05823_));
 sg13g2_buf_1 _23281_ (.A(_05823_),
    .X(_05824_));
 sg13g2_buf_1 _23282_ (.A(_05824_),
    .X(_05825_));
 sg13g2_mux2_1 _23283_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(_03399_),
    .S(net230),
    .X(_01141_));
 sg13g2_mux2_1 _23284_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net524),
    .S(net230),
    .X(_01142_));
 sg13g2_mux2_1 _23285_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(net641),
    .S(net230),
    .X(_01143_));
 sg13g2_mux2_1 _23286_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net591),
    .S(net230),
    .X(_01144_));
 sg13g2_mux2_1 _23287_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(net840),
    .S(net230),
    .X(_01145_));
 sg13g2_mux2_1 _23288_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net716),
    .S(net230),
    .X(_01146_));
 sg13g2_mux2_1 _23289_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net715),
    .S(_05825_),
    .X(_01147_));
 sg13g2_mux2_1 _23290_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net839),
    .S(net230),
    .X(_01148_));
 sg13g2_mux2_1 _23291_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net838),
    .S(_05825_),
    .X(_01149_));
 sg13g2_mux2_1 _23292_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net949),
    .S(net230),
    .X(_01150_));
 sg13g2_mux2_1 _23293_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(_03387_),
    .S(_05824_),
    .X(_01151_));
 sg13g2_mux2_1 _23294_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net468),
    .S(_05824_),
    .X(_01152_));
 sg13g2_buf_1 _23295_ (.A(_05820_),
    .X(_05826_));
 sg13g2_nand3_1 _23296_ (.B(_05792_),
    .C(_05806_),
    .A(_10594_),
    .Y(_05827_));
 sg13g2_buf_1 _23297_ (.A(_05827_),
    .X(_05828_));
 sg13g2_nor3_2 _23298_ (.A(net938),
    .B(net835),
    .C(_05828_),
    .Y(_05829_));
 sg13g2_nor2b_1 _23299_ (.A(net394),
    .B_N(_05829_),
    .Y(_05830_));
 sg13g2_buf_1 _23300_ (.A(_05830_),
    .X(_05831_));
 sg13g2_buf_1 _23301_ (.A(_05831_),
    .X(_05832_));
 sg13g2_mux2_1 _23302_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(_03399_),
    .S(net309),
    .X(_01153_));
 sg13g2_mux2_1 _23303_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net524),
    .S(net309),
    .X(_01154_));
 sg13g2_mux2_1 _23304_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(net641),
    .S(net309),
    .X(_01155_));
 sg13g2_mux2_1 _23305_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net591),
    .S(_05832_),
    .X(_01156_));
 sg13g2_mux2_1 _23306_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net840),
    .S(net309),
    .X(_01157_));
 sg13g2_mux2_1 _23307_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net716),
    .S(net309),
    .X(_01158_));
 sg13g2_mux2_1 _23308_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net715),
    .S(net309),
    .X(_01159_));
 sg13g2_mux2_1 _23309_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(net839),
    .S(net309),
    .X(_01160_));
 sg13g2_mux2_1 _23310_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net838),
    .S(net309),
    .X(_01161_));
 sg13g2_mux2_1 _23311_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net949),
    .S(_05832_),
    .X(_01162_));
 sg13g2_buf_1 _23312_ (.A(net595),
    .X(_05833_));
 sg13g2_mux2_1 _23313_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net511),
    .S(_05831_),
    .X(_01163_));
 sg13g2_mux2_1 _23314_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net468),
    .S(_05831_),
    .X(_01164_));
 sg13g2_buf_1 _23315_ (.A(_03397_),
    .X(_05834_));
 sg13g2_inv_2 _23316_ (.Y(_05835_),
    .A(net1090));
 sg13g2_nand2_1 _23317_ (.Y(_05836_),
    .A(_05835_),
    .B(_05772_));
 sg13g2_nor2_1 _23318_ (.A(_05828_),
    .B(_05836_),
    .Y(_05837_));
 sg13g2_buf_2 _23319_ (.A(_05837_),
    .X(_05838_));
 sg13g2_nor2b_1 _23320_ (.A(_05826_),
    .B_N(_05838_),
    .Y(_05839_));
 sg13g2_buf_1 _23321_ (.A(_05839_),
    .X(_05840_));
 sg13g2_buf_1 _23322_ (.A(_05840_),
    .X(_05841_));
 sg13g2_mux2_1 _23323_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(_05834_),
    .S(net308),
    .X(_01165_));
 sg13g2_mux2_1 _23324_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net524),
    .S(net308),
    .X(_01166_));
 sg13g2_mux2_1 _23325_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(_03417_),
    .S(net308),
    .X(_01167_));
 sg13g2_mux2_1 _23326_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net591),
    .S(_05841_),
    .X(_01168_));
 sg13g2_mux2_1 _23327_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(net840),
    .S(net308),
    .X(_01169_));
 sg13g2_mux2_1 _23328_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net716),
    .S(net308),
    .X(_01170_));
 sg13g2_mux2_1 _23329_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net715),
    .S(net308),
    .X(_01171_));
 sg13g2_mux2_1 _23330_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(net839),
    .S(net308),
    .X(_01172_));
 sg13g2_mux2_1 _23331_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net838),
    .S(net308),
    .X(_01173_));
 sg13g2_mux2_1 _23332_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net949),
    .S(_05841_),
    .X(_01174_));
 sg13g2_mux2_1 _23333_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net511),
    .S(_05840_),
    .X(_01175_));
 sg13g2_mux2_1 _23334_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(_03415_),
    .S(_05840_),
    .X(_01176_));
 sg13g2_nor2b_1 _23335_ (.A(net1090),
    .B_N(_10614_),
    .Y(_05842_));
 sg13g2_buf_1 _23336_ (.A(_05842_),
    .X(_05843_));
 sg13g2_nand2b_1 _23337_ (.Y(_05844_),
    .B(_05843_),
    .A_N(_05815_));
 sg13g2_buf_1 _23338_ (.A(_05844_),
    .X(_05845_));
 sg13g2_nor2_1 _23339_ (.A(_05822_),
    .B(_05845_),
    .Y(_05846_));
 sg13g2_buf_1 _23340_ (.A(_05846_),
    .X(_05847_));
 sg13g2_buf_1 _23341_ (.A(_05847_),
    .X(_05848_));
 sg13g2_mux2_1 _23342_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net331),
    .S(net229),
    .X(_01177_));
 sg13g2_mux2_1 _23343_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(_03416_),
    .S(net229),
    .X(_01178_));
 sg13g2_mux2_1 _23344_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(_03417_),
    .S(net229),
    .X(_01179_));
 sg13g2_mux2_1 _23345_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(net591),
    .S(net229),
    .X(_01180_));
 sg13g2_mux2_1 _23346_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(net840),
    .S(net229),
    .X(_01181_));
 sg13g2_mux2_1 _23347_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(net716),
    .S(net229),
    .X(_01182_));
 sg13g2_mux2_1 _23348_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(net715),
    .S(_05848_),
    .X(_01183_));
 sg13g2_mux2_1 _23349_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(net839),
    .S(net229),
    .X(_01184_));
 sg13g2_mux2_1 _23350_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(net838),
    .S(_05848_),
    .X(_01185_));
 sg13g2_mux2_1 _23351_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net949),
    .S(net229),
    .X(_01186_));
 sg13g2_mux2_1 _23352_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net511),
    .S(_05847_),
    .X(_01187_));
 sg13g2_mux2_1 _23353_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(_03415_),
    .S(_05847_),
    .X(_01188_));
 sg13g2_or2_1 _23354_ (.X(_05849_),
    .B(_05820_),
    .A(_05781_));
 sg13g2_buf_1 _23355_ (.A(_05849_),
    .X(_05850_));
 sg13g2_nor2_1 _23356_ (.A(_05845_),
    .B(_05850_),
    .Y(_05851_));
 sg13g2_buf_1 _23357_ (.A(_05851_),
    .X(_05852_));
 sg13g2_buf_1 _23358_ (.A(_05852_),
    .X(_05853_));
 sg13g2_mux2_1 _23359_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net331),
    .S(net228),
    .X(_01189_));
 sg13g2_mux2_1 _23360_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(_03416_),
    .S(net228),
    .X(_01190_));
 sg13g2_buf_1 _23361_ (.A(net890),
    .X(_05854_));
 sg13g2_mux2_1 _23362_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net708),
    .S(net228),
    .X(_01191_));
 sg13g2_mux2_1 _23363_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(net591),
    .S(net228),
    .X(_01192_));
 sg13g2_mux2_1 _23364_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(_03426_),
    .S(net228),
    .X(_01193_));
 sg13g2_mux2_1 _23365_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(_03427_),
    .S(net228),
    .X(_01194_));
 sg13g2_mux2_1 _23366_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(_03428_),
    .S(net228),
    .X(_01195_));
 sg13g2_mux2_1 _23367_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net839),
    .S(net228),
    .X(_01196_));
 sg13g2_mux2_1 _23368_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(net838),
    .S(_05853_),
    .X(_01197_));
 sg13g2_mux2_1 _23369_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net949),
    .S(_05853_),
    .X(_01198_));
 sg13g2_mux2_1 _23370_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net511),
    .S(_05852_),
    .X(_01199_));
 sg13g2_buf_1 _23371_ (.A(_09313_),
    .X(_05855_));
 sg13g2_mux2_1 _23372_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net510),
    .S(_05852_),
    .X(_01200_));
 sg13g2_buf_1 _23373_ (.A(_05820_),
    .X(_05856_));
 sg13g2_nor3_1 _23374_ (.A(net709),
    .B(_05856_),
    .C(_05845_),
    .Y(_05857_));
 sg13g2_buf_1 _23375_ (.A(_05857_),
    .X(_05858_));
 sg13g2_buf_1 _23376_ (.A(_05858_),
    .X(_05859_));
 sg13g2_mux2_1 _23377_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(net331),
    .S(net307),
    .X(_01201_));
 sg13g2_buf_1 _23378_ (.A(_09478_),
    .X(_05860_));
 sg13g2_mux2_1 _23379_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(_05860_),
    .S(net307),
    .X(_01202_));
 sg13g2_mux2_1 _23380_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(net708),
    .S(net307),
    .X(_01203_));
 sg13g2_mux2_1 _23381_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(_03425_),
    .S(net307),
    .X(_01204_));
 sg13g2_mux2_1 _23382_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(_03426_),
    .S(net307),
    .X(_01205_));
 sg13g2_mux2_1 _23383_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(_03427_),
    .S(net307),
    .X(_01206_));
 sg13g2_mux2_1 _23384_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(_03428_),
    .S(net307),
    .X(_01207_));
 sg13g2_mux2_1 _23385_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(_03429_),
    .S(net307),
    .X(_01208_));
 sg13g2_mux2_1 _23386_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(_03433_),
    .S(_05859_),
    .X(_01209_));
 sg13g2_mux2_1 _23387_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(_03424_),
    .S(_05859_),
    .X(_01210_));
 sg13g2_mux2_1 _23388_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(net511),
    .S(_05858_),
    .X(_01211_));
 sg13g2_mux2_1 _23389_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(net510),
    .S(_05858_),
    .X(_01212_));
 sg13g2_nor3_1 _23390_ (.A(_05791_),
    .B(_05856_),
    .C(_05845_),
    .Y(_05861_));
 sg13g2_buf_1 _23391_ (.A(_05861_),
    .X(_05862_));
 sg13g2_buf_1 _23392_ (.A(_05862_),
    .X(_05863_));
 sg13g2_mux2_1 _23393_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(_05834_),
    .S(net306),
    .X(_01213_));
 sg13g2_mux2_1 _23394_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(net578),
    .S(net306),
    .X(_01214_));
 sg13g2_mux2_1 _23395_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(_05854_),
    .S(net306),
    .X(_01215_));
 sg13g2_mux2_1 _23396_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(_03425_),
    .S(net306),
    .X(_01216_));
 sg13g2_buf_1 _23397_ (.A(_02914_),
    .X(_05864_));
 sg13g2_mux2_1 _23398_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(net833),
    .S(net306),
    .X(_01217_));
 sg13g2_buf_1 _23399_ (.A(_09014_),
    .X(_05865_));
 sg13g2_mux2_1 _23400_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(_05865_),
    .S(net306),
    .X(_01218_));
 sg13g2_buf_1 _23401_ (.A(_09012_),
    .X(_05866_));
 sg13g2_mux2_1 _23402_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(_05866_),
    .S(net306),
    .X(_01219_));
 sg13g2_mux2_1 _23403_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(_03429_),
    .S(net306),
    .X(_01220_));
 sg13g2_mux2_1 _23404_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(_03433_),
    .S(_05863_),
    .X(_01221_));
 sg13g2_mux2_1 _23405_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(_03424_),
    .S(_05863_),
    .X(_01222_));
 sg13g2_mux2_1 _23406_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(_05833_),
    .S(_05862_),
    .X(_01223_));
 sg13g2_mux2_1 _23407_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_05855_),
    .S(_05862_),
    .X(_01224_));
 sg13g2_nand2b_1 _23408_ (.Y(_05867_),
    .B(net938),
    .A_N(net939));
 sg13g2_nor2_2 _23409_ (.A(_10594_),
    .B(_10566_),
    .Y(_05868_));
 sg13g2_nand2b_1 _23410_ (.Y(_05869_),
    .B(_05868_),
    .A_N(net942));
 sg13g2_buf_1 _23411_ (.A(_05869_),
    .X(_05870_));
 sg13g2_nor3_1 _23412_ (.A(net393),
    .B(_05867_),
    .C(_05870_),
    .Y(_05871_));
 sg13g2_buf_1 _23413_ (.A(_05871_),
    .X(_05872_));
 sg13g2_buf_1 _23414_ (.A(_05872_),
    .X(_05873_));
 sg13g2_mux2_1 _23415_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net331),
    .S(net305),
    .X(_01225_));
 sg13g2_mux2_1 _23416_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net578),
    .S(net305),
    .X(_01226_));
 sg13g2_mux2_1 _23417_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net708),
    .S(net305),
    .X(_01227_));
 sg13g2_buf_1 _23418_ (.A(net643),
    .X(_05874_));
 sg13g2_mux2_1 _23419_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net577),
    .S(net305),
    .X(_01228_));
 sg13g2_mux2_1 _23420_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net833),
    .S(net305),
    .X(_01229_));
 sg13g2_mux2_1 _23421_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net832),
    .S(_05873_),
    .X(_01230_));
 sg13g2_mux2_1 _23422_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net831),
    .S(_05873_),
    .X(_01231_));
 sg13g2_buf_1 _23423_ (.A(_10627_),
    .X(_05875_));
 sg13g2_mux2_1 _23424_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net937),
    .S(net305),
    .X(_01232_));
 sg13g2_buf_1 _23425_ (.A(net1089),
    .X(_05876_));
 sg13g2_mux2_1 _23426_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net936),
    .S(net305),
    .X(_01233_));
 sg13g2_buf_1 _23427_ (.A(net1094),
    .X(_05877_));
 sg13g2_mux2_1 _23428_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net935),
    .S(net305),
    .X(_01234_));
 sg13g2_mux2_1 _23429_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(net511),
    .S(_05872_),
    .X(_01235_));
 sg13g2_mux2_1 _23430_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net510),
    .S(_05872_),
    .X(_01236_));
 sg13g2_nor2_1 _23431_ (.A(_05835_),
    .B(net834),
    .Y(_05878_));
 sg13g2_nor2_1 _23432_ (.A(_05794_),
    .B(_05850_),
    .Y(_05879_));
 sg13g2_nand2_1 _23433_ (.Y(_05880_),
    .A(_05878_),
    .B(_05879_));
 sg13g2_buf_2 _23434_ (.A(_05880_),
    .X(_05881_));
 sg13g2_buf_1 _23435_ (.A(_05881_),
    .X(_05882_));
 sg13g2_nand2_1 _23436_ (.Y(_05883_),
    .A(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .B(_05881_));
 sg13g2_o21ai_1 _23437_ (.B1(_05883_),
    .Y(_01237_),
    .A1(_03704_),
    .A2(net197));
 sg13g2_mux2_1 _23438_ (.A0(_03696_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .S(net197),
    .X(_01238_));
 sg13g2_mux2_1 _23439_ (.A0(_03697_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .S(net197),
    .X(_01239_));
 sg13g2_nand2_1 _23440_ (.Y(_05884_),
    .A(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .B(_05881_));
 sg13g2_o21ai_1 _23441_ (.B1(_05884_),
    .Y(_01240_),
    .A1(_02908_),
    .A2(net197));
 sg13g2_mux2_1 _23442_ (.A0(_02916_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .S(net197),
    .X(_01241_));
 sg13g2_mux2_1 _23443_ (.A0(_02918_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .S(net197),
    .X(_01242_));
 sg13g2_mux2_1 _23444_ (.A0(_02920_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .S(_05882_),
    .X(_01243_));
 sg13g2_mux2_1 _23445_ (.A0(_02922_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .S(_05882_),
    .X(_01244_));
 sg13g2_mux2_1 _23446_ (.A0(_02924_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .S(_05881_),
    .X(_01245_));
 sg13g2_mux2_1 _23447_ (.A0(_02926_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .S(_05881_),
    .X(_01246_));
 sg13g2_nand2_1 _23448_ (.Y(_05885_),
    .A(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .B(_05881_));
 sg13g2_o21ai_1 _23449_ (.B1(_05885_),
    .Y(_01247_),
    .A1(_03693_),
    .A2(net197));
 sg13g2_mux2_1 _23450_ (.A0(_03695_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .S(_05881_),
    .X(_01248_));
 sg13g2_nand2_1 _23451_ (.Y(_05886_),
    .A(net941),
    .B(_05792_));
 sg13g2_nand2b_1 _23452_ (.Y(_05887_),
    .B(net938),
    .A_N(net835));
 sg13g2_nor3_2 _23453_ (.A(net834),
    .B(_05886_),
    .C(_05887_),
    .Y(_05888_));
 sg13g2_nor2b_1 _23454_ (.A(net394),
    .B_N(_05888_),
    .Y(_05889_));
 sg13g2_buf_1 _23455_ (.A(_05889_),
    .X(_05890_));
 sg13g2_buf_1 _23456_ (.A(_05890_),
    .X(_05891_));
 sg13g2_mux2_1 _23457_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net331),
    .S(net304),
    .X(_01249_));
 sg13g2_mux2_1 _23458_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(net578),
    .S(net304),
    .X(_01250_));
 sg13g2_mux2_1 _23459_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net708),
    .S(net304),
    .X(_01251_));
 sg13g2_mux2_1 _23460_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net577),
    .S(net304),
    .X(_01252_));
 sg13g2_mux2_1 _23461_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net833),
    .S(net304),
    .X(_01253_));
 sg13g2_mux2_1 _23462_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(net832),
    .S(_05891_),
    .X(_01254_));
 sg13g2_mux2_1 _23463_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(net831),
    .S(_05891_),
    .X(_01255_));
 sg13g2_mux2_1 _23464_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(net937),
    .S(net304),
    .X(_01256_));
 sg13g2_mux2_1 _23465_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net936),
    .S(net304),
    .X(_01257_));
 sg13g2_mux2_1 _23466_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net935),
    .S(net304),
    .X(_01258_));
 sg13g2_mux2_1 _23467_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net511),
    .S(_05890_),
    .X(_01259_));
 sg13g2_mux2_1 _23468_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net510),
    .S(_05890_),
    .X(_01260_));
 sg13g2_nand2_1 _23469_ (.Y(_05892_),
    .A(net1090),
    .B(net835));
 sg13g2_nor3_1 _23470_ (.A(net834),
    .B(_05886_),
    .C(_05892_),
    .Y(_05893_));
 sg13g2_buf_2 _23471_ (.A(_05893_),
    .X(_05894_));
 sg13g2_nor2b_1 _23472_ (.A(net394),
    .B_N(_05894_),
    .Y(_05895_));
 sg13g2_buf_1 _23473_ (.A(_05895_),
    .X(_05896_));
 sg13g2_buf_1 _23474_ (.A(_05896_),
    .X(_05897_));
 sg13g2_mux2_1 _23475_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(net331),
    .S(net303),
    .X(_01261_));
 sg13g2_mux2_1 _23476_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(net578),
    .S(net303),
    .X(_01262_));
 sg13g2_mux2_1 _23477_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(net708),
    .S(net303),
    .X(_01263_));
 sg13g2_mux2_1 _23478_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net577),
    .S(net303),
    .X(_01264_));
 sg13g2_mux2_1 _23479_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(_05864_),
    .S(net303),
    .X(_01265_));
 sg13g2_mux2_1 _23480_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(net832),
    .S(_05897_),
    .X(_01266_));
 sg13g2_mux2_1 _23481_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(net831),
    .S(_05897_),
    .X(_01267_));
 sg13g2_mux2_1 _23482_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net937),
    .S(net303),
    .X(_01268_));
 sg13g2_mux2_1 _23483_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(net936),
    .S(net303),
    .X(_01269_));
 sg13g2_mux2_1 _23484_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(net935),
    .S(net303),
    .X(_01270_));
 sg13g2_mux2_1 _23485_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net511),
    .S(_05896_),
    .X(_01271_));
 sg13g2_mux2_1 _23486_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net510),
    .S(_05896_),
    .X(_01272_));
 sg13g2_nor2_1 _23487_ (.A(_05818_),
    .B(_05850_),
    .Y(_05898_));
 sg13g2_buf_1 _23488_ (.A(_05898_),
    .X(_05899_));
 sg13g2_buf_1 _23489_ (.A(_05899_),
    .X(_05900_));
 sg13g2_mux2_1 _23490_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(net331),
    .S(net227),
    .X(_01273_));
 sg13g2_mux2_1 _23491_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(_05860_),
    .S(net227),
    .X(_01274_));
 sg13g2_mux2_1 _23492_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(_05854_),
    .S(net227),
    .X(_01275_));
 sg13g2_mux2_1 _23493_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05874_),
    .S(net227),
    .X(_01276_));
 sg13g2_mux2_1 _23494_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(_05864_),
    .S(net227),
    .X(_01277_));
 sg13g2_mux2_1 _23495_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(_05865_),
    .S(net227),
    .X(_01278_));
 sg13g2_mux2_1 _23496_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(_05866_),
    .S(_05900_),
    .X(_01279_));
 sg13g2_mux2_1 _23497_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(net937),
    .S(net227),
    .X(_01280_));
 sg13g2_mux2_1 _23498_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(_05876_),
    .S(net227),
    .X(_01281_));
 sg13g2_mux2_1 _23499_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(_05877_),
    .S(_05900_),
    .X(_01282_));
 sg13g2_mux2_1 _23500_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(_05833_),
    .S(_05899_),
    .X(_01283_));
 sg13g2_mux2_1 _23501_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05855_),
    .S(_05899_),
    .X(_01284_));
 sg13g2_or2_1 _23502_ (.X(_05901_),
    .B(_05867_),
    .A(_05815_));
 sg13g2_buf_1 _23503_ (.A(_05901_),
    .X(_05902_));
 sg13g2_nor2_1 _23504_ (.A(_05822_),
    .B(_05902_),
    .Y(_05903_));
 sg13g2_buf_1 _23505_ (.A(_05903_),
    .X(_05904_));
 sg13g2_buf_1 _23506_ (.A(_05904_),
    .X(_05905_));
 sg13g2_mux2_1 _23507_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net331),
    .S(net226),
    .X(_01285_));
 sg13g2_mux2_1 _23508_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net578),
    .S(net226),
    .X(_01286_));
 sg13g2_mux2_1 _23509_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net708),
    .S(net226),
    .X(_01287_));
 sg13g2_mux2_1 _23510_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net577),
    .S(net226),
    .X(_01288_));
 sg13g2_mux2_1 _23511_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net833),
    .S(net226),
    .X(_01289_));
 sg13g2_mux2_1 _23512_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net832),
    .S(_05905_),
    .X(_01290_));
 sg13g2_mux2_1 _23513_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net831),
    .S(_05905_),
    .X(_01291_));
 sg13g2_mux2_1 _23514_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net937),
    .S(net226),
    .X(_01292_));
 sg13g2_mux2_1 _23515_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net936),
    .S(net226),
    .X(_01293_));
 sg13g2_mux2_1 _23516_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net935),
    .S(net226),
    .X(_01294_));
 sg13g2_buf_1 _23517_ (.A(_09231_),
    .X(_05906_));
 sg13g2_mux2_1 _23518_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net576),
    .S(_05904_),
    .X(_01295_));
 sg13g2_mux2_1 _23519_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net510),
    .S(_05904_),
    .X(_01296_));
 sg13g2_buf_1 _23520_ (.A(_03397_),
    .X(_05907_));
 sg13g2_nor2_1 _23521_ (.A(_05850_),
    .B(_05902_),
    .Y(_05908_));
 sg13g2_buf_1 _23522_ (.A(_05908_),
    .X(_05909_));
 sg13g2_buf_1 _23523_ (.A(_05909_),
    .X(_05910_));
 sg13g2_mux2_1 _23524_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net330),
    .S(net225),
    .X(_01297_));
 sg13g2_mux2_1 _23525_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net578),
    .S(net225),
    .X(_01298_));
 sg13g2_mux2_1 _23526_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net708),
    .S(net225),
    .X(_01299_));
 sg13g2_mux2_1 _23527_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net577),
    .S(net225),
    .X(_01300_));
 sg13g2_mux2_1 _23528_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net833),
    .S(net225),
    .X(_01301_));
 sg13g2_mux2_1 _23529_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net832),
    .S(_05910_),
    .X(_01302_));
 sg13g2_mux2_1 _23530_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net831),
    .S(_05910_),
    .X(_01303_));
 sg13g2_mux2_1 _23531_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net937),
    .S(net225),
    .X(_01304_));
 sg13g2_mux2_1 _23532_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net936),
    .S(net225),
    .X(_01305_));
 sg13g2_mux2_1 _23533_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net935),
    .S(net225),
    .X(_01306_));
 sg13g2_mux2_1 _23534_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net576),
    .S(_05909_),
    .X(_01307_));
 sg13g2_mux2_1 _23535_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net510),
    .S(_05909_),
    .X(_01308_));
 sg13g2_nor3_1 _23536_ (.A(net709),
    .B(net393),
    .C(_05902_),
    .Y(_05911_));
 sg13g2_buf_1 _23537_ (.A(_05911_),
    .X(_05912_));
 sg13g2_buf_1 _23538_ (.A(_05912_),
    .X(_05913_));
 sg13g2_mux2_1 _23539_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net330),
    .S(net302),
    .X(_01309_));
 sg13g2_mux2_1 _23540_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net578),
    .S(net302),
    .X(_01310_));
 sg13g2_mux2_1 _23541_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net708),
    .S(net302),
    .X(_01311_));
 sg13g2_mux2_1 _23542_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net577),
    .S(net302),
    .X(_01312_));
 sg13g2_mux2_1 _23543_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net833),
    .S(net302),
    .X(_01313_));
 sg13g2_mux2_1 _23544_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net832),
    .S(_05913_),
    .X(_01314_));
 sg13g2_mux2_1 _23545_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net831),
    .S(_05913_),
    .X(_01315_));
 sg13g2_mux2_1 _23546_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net937),
    .S(net302),
    .X(_01316_));
 sg13g2_mux2_1 _23547_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net936),
    .S(net302),
    .X(_01317_));
 sg13g2_mux2_1 _23548_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net935),
    .S(net302),
    .X(_01318_));
 sg13g2_mux2_1 _23549_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net576),
    .S(_05912_),
    .X(_01319_));
 sg13g2_mux2_1 _23550_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net510),
    .S(_05912_),
    .X(_01320_));
 sg13g2_nor3_1 _23551_ (.A(_05791_),
    .B(net393),
    .C(_05902_),
    .Y(_05914_));
 sg13g2_buf_1 _23552_ (.A(_05914_),
    .X(_05915_));
 sg13g2_buf_1 _23553_ (.A(_05915_),
    .X(_05916_));
 sg13g2_mux2_1 _23554_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net330),
    .S(net301),
    .X(_01321_));
 sg13g2_mux2_1 _23555_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net578),
    .S(net301),
    .X(_01322_));
 sg13g2_buf_1 _23556_ (.A(_09428_),
    .X(_05917_));
 sg13g2_mux2_1 _23557_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net707),
    .S(net301),
    .X(_01323_));
 sg13g2_mux2_1 _23558_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net577),
    .S(net301),
    .X(_01324_));
 sg13g2_mux2_1 _23559_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net833),
    .S(net301),
    .X(_01325_));
 sg13g2_mux2_1 _23560_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(net832),
    .S(_05916_),
    .X(_01326_));
 sg13g2_mux2_1 _23561_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net831),
    .S(_05916_),
    .X(_01327_));
 sg13g2_mux2_1 _23562_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net937),
    .S(net301),
    .X(_01328_));
 sg13g2_mux2_1 _23563_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net936),
    .S(net301),
    .X(_01329_));
 sg13g2_mux2_1 _23564_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net935),
    .S(net301),
    .X(_01330_));
 sg13g2_mux2_1 _23565_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net576),
    .S(_05915_),
    .X(_01331_));
 sg13g2_buf_1 _23566_ (.A(_09313_),
    .X(_05918_));
 sg13g2_mux2_1 _23567_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net509),
    .S(_05915_),
    .X(_01332_));
 sg13g2_nand2_1 _23568_ (.Y(_05919_),
    .A(net1090),
    .B(net834));
 sg13g2_nor3_1 _23569_ (.A(net393),
    .B(_05870_),
    .C(_05919_),
    .Y(_05920_));
 sg13g2_buf_1 _23570_ (.A(_05920_),
    .X(_05921_));
 sg13g2_buf_1 _23571_ (.A(_05921_),
    .X(_05922_));
 sg13g2_mux2_1 _23572_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net330),
    .S(net300),
    .X(_01333_));
 sg13g2_buf_1 _23573_ (.A(net672),
    .X(_05923_));
 sg13g2_mux2_1 _23574_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net575),
    .S(net300),
    .X(_01334_));
 sg13g2_mux2_1 _23575_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net707),
    .S(net300),
    .X(_01335_));
 sg13g2_mux2_1 _23576_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net577),
    .S(net300),
    .X(_01336_));
 sg13g2_mux2_1 _23577_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net833),
    .S(net300),
    .X(_01337_));
 sg13g2_mux2_1 _23578_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net832),
    .S(_05922_),
    .X(_01338_));
 sg13g2_mux2_1 _23579_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net831),
    .S(_05922_),
    .X(_01339_));
 sg13g2_mux2_1 _23580_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(_05875_),
    .S(net300),
    .X(_01340_));
 sg13g2_mux2_1 _23581_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(_05876_),
    .S(net300),
    .X(_01341_));
 sg13g2_mux2_1 _23582_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net935),
    .S(net300),
    .X(_01342_));
 sg13g2_mux2_1 _23583_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net576),
    .S(_05921_),
    .X(_01343_));
 sg13g2_mux2_1 _23584_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net509),
    .S(_05921_),
    .X(_01344_));
 sg13g2_nand3_1 _23585_ (.B(_05807_),
    .C(_05879_),
    .A(_05816_),
    .Y(_05924_));
 sg13g2_buf_2 _23586_ (.A(_05924_),
    .X(_05925_));
 sg13g2_buf_1 _23587_ (.A(_05925_),
    .X(_05926_));
 sg13g2_nand2_1 _23588_ (.Y(_05927_),
    .A(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .B(_05925_));
 sg13g2_o21ai_1 _23589_ (.B1(_05927_),
    .Y(_01345_),
    .A1(_03704_),
    .A2(net196));
 sg13g2_mux2_1 _23590_ (.A0(_03696_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .S(net196),
    .X(_01346_));
 sg13g2_mux2_1 _23591_ (.A0(_03697_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .S(net196),
    .X(_01347_));
 sg13g2_nand2_1 _23592_ (.Y(_05928_),
    .A(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .B(_05925_));
 sg13g2_o21ai_1 _23593_ (.B1(_05928_),
    .Y(_01348_),
    .A1(_02908_),
    .A2(net196));
 sg13g2_mux2_1 _23594_ (.A0(_02916_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .S(net196),
    .X(_01349_));
 sg13g2_mux2_1 _23595_ (.A0(_02918_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .S(_05926_),
    .X(_01350_));
 sg13g2_mux2_1 _23596_ (.A0(_02920_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .S(_05926_),
    .X(_01351_));
 sg13g2_mux2_1 _23597_ (.A0(_02922_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .S(net196),
    .X(_01352_));
 sg13g2_mux2_1 _23598_ (.A0(_02924_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .S(_05925_),
    .X(_01353_));
 sg13g2_mux2_1 _23599_ (.A0(_02926_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .S(_05925_),
    .X(_01354_));
 sg13g2_nand2_1 _23600_ (.Y(_05929_),
    .A(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .B(_05925_));
 sg13g2_o21ai_1 _23601_ (.B1(_05929_),
    .Y(_01355_),
    .A1(_03693_),
    .A2(net196));
 sg13g2_mux2_1 _23602_ (.A0(_03695_),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .S(_05925_),
    .X(_01356_));
 sg13g2_nor2_2 _23603_ (.A(_05828_),
    .B(_05887_),
    .Y(_05930_));
 sg13g2_nor2b_1 _23604_ (.A(net394),
    .B_N(_05930_),
    .Y(_05931_));
 sg13g2_buf_1 _23605_ (.A(_05931_),
    .X(_05932_));
 sg13g2_buf_1 _23606_ (.A(_05932_),
    .X(_05933_));
 sg13g2_mux2_1 _23607_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(_05907_),
    .S(net299),
    .X(_01357_));
 sg13g2_mux2_1 _23608_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net575),
    .S(net299),
    .X(_01358_));
 sg13g2_mux2_1 _23609_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net707),
    .S(net299),
    .X(_01359_));
 sg13g2_mux2_1 _23610_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(_05874_),
    .S(net299),
    .X(_01360_));
 sg13g2_buf_1 _23611_ (.A(net953),
    .X(_05934_));
 sg13g2_mux2_1 _23612_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(_05934_),
    .S(net299),
    .X(_01361_));
 sg13g2_buf_1 _23613_ (.A(_09014_),
    .X(_05935_));
 sg13g2_mux2_1 _23614_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net829),
    .S(_05933_),
    .X(_01362_));
 sg13g2_buf_1 _23615_ (.A(net1038),
    .X(_05936_));
 sg13g2_mux2_1 _23616_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net828),
    .S(_05933_),
    .X(_01363_));
 sg13g2_mux2_1 _23617_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(_05875_),
    .S(net299),
    .X(_01364_));
 sg13g2_mux2_1 _23618_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net936),
    .S(net299),
    .X(_01365_));
 sg13g2_mux2_1 _23619_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(_05877_),
    .S(net299),
    .X(_01366_));
 sg13g2_mux2_1 _23620_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(_05906_),
    .S(_05932_),
    .X(_01367_));
 sg13g2_mux2_1 _23621_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net509),
    .S(_05932_),
    .X(_01368_));
 sg13g2_nor2_1 _23622_ (.A(_05828_),
    .B(_05892_),
    .Y(_05937_));
 sg13g2_buf_1 _23623_ (.A(_05937_),
    .X(_05938_));
 sg13g2_nor2b_1 _23624_ (.A(net394),
    .B_N(_05938_),
    .Y(_05939_));
 sg13g2_buf_1 _23625_ (.A(_05939_),
    .X(_05940_));
 sg13g2_buf_1 _23626_ (.A(_05940_),
    .X(_05941_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(_05907_),
    .S(net298),
    .X(_01369_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net575),
    .S(net298),
    .X(_01370_));
 sg13g2_mux2_1 _23629_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net707),
    .S(net298),
    .X(_01371_));
 sg13g2_buf_1 _23630_ (.A(net643),
    .X(_05942_));
 sg13g2_mux2_1 _23631_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net574),
    .S(net298),
    .X(_01372_));
 sg13g2_mux2_1 _23632_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(_05934_),
    .S(net298),
    .X(_01373_));
 sg13g2_mux2_1 _23633_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net829),
    .S(net298),
    .X(_01374_));
 sg13g2_mux2_1 _23634_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net828),
    .S(_05941_),
    .X(_01375_));
 sg13g2_buf_1 _23635_ (.A(_10627_),
    .X(_05943_));
 sg13g2_mux2_1 _23636_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net934),
    .S(net298),
    .X(_01376_));
 sg13g2_buf_1 _23637_ (.A(net1089),
    .X(_05944_));
 sg13g2_mux2_1 _23638_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net933),
    .S(net298),
    .X(_01377_));
 sg13g2_buf_1 _23639_ (.A(net1094),
    .X(_05945_));
 sg13g2_mux2_1 _23640_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net932),
    .S(_05941_),
    .X(_01378_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net576),
    .S(_05940_),
    .X(_01379_));
 sg13g2_mux2_1 _23642_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net509),
    .S(_05940_),
    .X(_01380_));
 sg13g2_or2_1 _23643_ (.X(_05946_),
    .B(_05919_),
    .A(_05815_));
 sg13g2_buf_1 _23644_ (.A(_05946_),
    .X(_05947_));
 sg13g2_nor2_1 _23645_ (.A(_05822_),
    .B(_05947_),
    .Y(_05948_));
 sg13g2_buf_1 _23646_ (.A(_05948_),
    .X(_05949_));
 sg13g2_buf_1 _23647_ (.A(_05949_),
    .X(_05950_));
 sg13g2_mux2_1 _23648_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net330),
    .S(net224),
    .X(_01381_));
 sg13g2_mux2_1 _23649_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net575),
    .S(net224),
    .X(_01382_));
 sg13g2_mux2_1 _23650_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net707),
    .S(net224),
    .X(_01383_));
 sg13g2_mux2_1 _23651_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net574),
    .S(net224),
    .X(_01384_));
 sg13g2_mux2_1 _23652_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net830),
    .S(net224),
    .X(_01385_));
 sg13g2_mux2_1 _23653_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net829),
    .S(net224),
    .X(_01386_));
 sg13g2_mux2_1 _23654_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net828),
    .S(_05950_),
    .X(_01387_));
 sg13g2_mux2_1 _23655_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net934),
    .S(net224),
    .X(_01388_));
 sg13g2_mux2_1 _23656_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net933),
    .S(net224),
    .X(_01389_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net932),
    .S(_05950_),
    .X(_01390_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(_05906_),
    .S(_05949_),
    .X(_01391_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net509),
    .S(_05949_),
    .X(_01392_));
 sg13g2_nor2_1 _23660_ (.A(_05850_),
    .B(_05947_),
    .Y(_05951_));
 sg13g2_buf_1 _23661_ (.A(_05951_),
    .X(_05952_));
 sg13g2_buf_1 _23662_ (.A(_05952_),
    .X(_05953_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net330),
    .S(net223),
    .X(_01393_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net575),
    .S(net223),
    .X(_01394_));
 sg13g2_mux2_1 _23665_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net707),
    .S(net223),
    .X(_01395_));
 sg13g2_mux2_1 _23666_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net574),
    .S(net223),
    .X(_01396_));
 sg13g2_mux2_1 _23667_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net830),
    .S(net223),
    .X(_01397_));
 sg13g2_mux2_1 _23668_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net829),
    .S(net223),
    .X(_01398_));
 sg13g2_mux2_1 _23669_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net828),
    .S(_05953_),
    .X(_01399_));
 sg13g2_mux2_1 _23670_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net934),
    .S(net223),
    .X(_01400_));
 sg13g2_mux2_1 _23671_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net933),
    .S(net223),
    .X(_01401_));
 sg13g2_mux2_1 _23672_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net932),
    .S(_05953_),
    .X(_01402_));
 sg13g2_mux2_1 _23673_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net576),
    .S(_05952_),
    .X(_01403_));
 sg13g2_mux2_1 _23674_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net509),
    .S(_05952_),
    .X(_01404_));
 sg13g2_nor3_1 _23675_ (.A(_05779_),
    .B(_05818_),
    .C(_05826_),
    .Y(_05954_));
 sg13g2_buf_1 _23676_ (.A(_05954_),
    .X(_05955_));
 sg13g2_buf_1 _23677_ (.A(_05955_),
    .X(_05956_));
 sg13g2_mux2_1 _23678_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net330),
    .S(net297),
    .X(_01405_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(_05923_),
    .S(net297),
    .X(_01406_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(_05917_),
    .S(net297),
    .X(_01407_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(net574),
    .S(net297),
    .X(_01408_));
 sg13g2_mux2_1 _23682_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(net830),
    .S(net297),
    .X(_01409_));
 sg13g2_mux2_1 _23683_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net829),
    .S(net297),
    .X(_01410_));
 sg13g2_mux2_1 _23684_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net828),
    .S(_05956_),
    .X(_01411_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(_05943_),
    .S(net297),
    .X(_01412_));
 sg13g2_mux2_1 _23686_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(_05944_),
    .S(net297),
    .X(_01413_));
 sg13g2_mux2_1 _23687_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(_05945_),
    .S(_05956_),
    .X(_01414_));
 sg13g2_mux2_1 _23688_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(net576),
    .S(_05955_),
    .X(_01415_));
 sg13g2_mux2_1 _23689_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(net509),
    .S(_05955_),
    .X(_01416_));
 sg13g2_nor3_1 _23690_ (.A(_05779_),
    .B(net393),
    .C(_05947_),
    .Y(_05957_));
 sg13g2_buf_1 _23691_ (.A(_05957_),
    .X(_05958_));
 sg13g2_buf_1 _23692_ (.A(_05958_),
    .X(_05959_));
 sg13g2_mux2_1 _23693_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net330),
    .S(net296),
    .X(_01417_));
 sg13g2_mux2_1 _23694_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net575),
    .S(net296),
    .X(_01418_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net707),
    .S(net296),
    .X(_01419_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(net574),
    .S(net296),
    .X(_01420_));
 sg13g2_mux2_1 _23697_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net830),
    .S(net296),
    .X(_01421_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net829),
    .S(net296),
    .X(_01422_));
 sg13g2_mux2_1 _23699_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net828),
    .S(_05959_),
    .X(_01423_));
 sg13g2_mux2_1 _23700_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net934),
    .S(net296),
    .X(_01424_));
 sg13g2_mux2_1 _23701_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(net933),
    .S(net296),
    .X(_01425_));
 sg13g2_mux2_1 _23702_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net932),
    .S(_05959_),
    .X(_01426_));
 sg13g2_mux2_1 _23703_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net595),
    .S(_05958_),
    .X(_01427_));
 sg13g2_mux2_1 _23704_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(_05918_),
    .S(_05958_),
    .X(_01428_));
 sg13g2_nor3_1 _23705_ (.A(_05791_),
    .B(net393),
    .C(_05947_),
    .Y(_05960_));
 sg13g2_buf_1 _23706_ (.A(_05960_),
    .X(_05961_));
 sg13g2_buf_1 _23707_ (.A(_05961_),
    .X(_05962_));
 sg13g2_mux2_1 _23708_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net335),
    .S(net295),
    .X(_01429_));
 sg13g2_mux2_1 _23709_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net575),
    .S(net295),
    .X(_01430_));
 sg13g2_mux2_1 _23710_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net707),
    .S(net295),
    .X(_01431_));
 sg13g2_mux2_1 _23711_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(net574),
    .S(net295),
    .X(_01432_));
 sg13g2_mux2_1 _23712_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net830),
    .S(net295),
    .X(_01433_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net829),
    .S(net295),
    .X(_01434_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(net828),
    .S(_05962_),
    .X(_01435_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(net934),
    .S(net295),
    .X(_01436_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net933),
    .S(net295),
    .X(_01437_));
 sg13g2_mux2_1 _23717_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net932),
    .S(_05962_),
    .X(_01438_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net595),
    .S(_05961_),
    .X(_01439_));
 sg13g2_mux2_1 _23719_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(_05918_),
    .S(_05961_),
    .X(_01440_));
 sg13g2_nor3_1 _23720_ (.A(_05791_),
    .B(_05818_),
    .C(net393),
    .Y(_05963_));
 sg13g2_buf_1 _23721_ (.A(_05963_),
    .X(_05964_));
 sg13g2_buf_1 _23722_ (.A(_05964_),
    .X(_05965_));
 sg13g2_mux2_1 _23723_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net335),
    .S(net294),
    .X(_01441_));
 sg13g2_mux2_1 _23724_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(_05923_),
    .S(net294),
    .X(_01442_));
 sg13g2_mux2_1 _23725_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(_05917_),
    .S(net294),
    .X(_01443_));
 sg13g2_mux2_1 _23726_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net574),
    .S(net294),
    .X(_01444_));
 sg13g2_mux2_1 _23727_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(net830),
    .S(net294),
    .X(_01445_));
 sg13g2_mux2_1 _23728_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(_05935_),
    .S(net294),
    .X(_01446_));
 sg13g2_mux2_1 _23729_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net828),
    .S(_05965_),
    .X(_01447_));
 sg13g2_mux2_1 _23730_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net934),
    .S(net294),
    .X(_01448_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(_05944_),
    .S(net294),
    .X(_01449_));
 sg13g2_mux2_1 _23732_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(net932),
    .S(_05965_),
    .X(_01450_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(net595),
    .S(_05964_),
    .X(_01451_));
 sg13g2_mux2_1 _23734_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(net509),
    .S(_05964_),
    .X(_01452_));
 sg13g2_nand2b_1 _23735_ (.Y(_05966_),
    .B(_10566_),
    .A_N(_05806_));
 sg13g2_nor3_1 _23736_ (.A(_05816_),
    .B(_05822_),
    .C(_05966_),
    .Y(_05967_));
 sg13g2_buf_1 _23737_ (.A(_05967_),
    .X(_05968_));
 sg13g2_buf_1 _23738_ (.A(_05968_),
    .X(_05969_));
 sg13g2_mux2_1 _23739_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net335),
    .S(net222),
    .X(_01453_));
 sg13g2_mux2_1 _23740_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net575),
    .S(net222),
    .X(_01454_));
 sg13g2_mux2_1 _23741_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net717),
    .S(_05969_),
    .X(_01455_));
 sg13g2_mux2_1 _23742_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net574),
    .S(net222),
    .X(_01456_));
 sg13g2_mux2_1 _23743_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net830),
    .S(net222),
    .X(_01457_));
 sg13g2_mux2_1 _23744_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net829),
    .S(net222),
    .X(_01458_));
 sg13g2_mux2_1 _23745_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(_05936_),
    .S(net222),
    .X(_01459_));
 sg13g2_mux2_1 _23746_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net934),
    .S(net222),
    .X(_01460_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net933),
    .S(net222),
    .X(_01461_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net932),
    .S(_05969_),
    .X(_01462_));
 sg13g2_mux2_1 _23749_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(_03386_),
    .S(_05968_),
    .X(_01463_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(net528),
    .S(_05968_),
    .X(_01464_));
 sg13g2_nor3_1 _23751_ (.A(_05777_),
    .B(_05836_),
    .C(_05966_),
    .Y(_05970_));
 sg13g2_buf_1 _23752_ (.A(_05970_),
    .X(_05971_));
 sg13g2_nor2b_1 _23753_ (.A(net394),
    .B_N(_05971_),
    .Y(_05972_));
 sg13g2_buf_1 _23754_ (.A(_05972_),
    .X(_05973_));
 sg13g2_buf_1 _23755_ (.A(_05973_),
    .X(_05974_));
 sg13g2_mux2_1 _23756_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net335),
    .S(net293),
    .X(_01465_));
 sg13g2_mux2_1 _23757_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(net594),
    .S(net293),
    .X(_01466_));
 sg13g2_mux2_1 _23758_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net717),
    .S(_05974_),
    .X(_01467_));
 sg13g2_mux2_1 _23759_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(_05942_),
    .S(net293),
    .X(_01468_));
 sg13g2_mux2_1 _23760_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net830),
    .S(net293),
    .X(_01469_));
 sg13g2_mux2_1 _23761_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(_05935_),
    .S(net293),
    .X(_01470_));
 sg13g2_mux2_1 _23762_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(_05936_),
    .S(net293),
    .X(_01471_));
 sg13g2_mux2_1 _23763_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net934),
    .S(net293),
    .X(_01472_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net933),
    .S(net293),
    .X(_01473_));
 sg13g2_mux2_1 _23765_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net932),
    .S(_05974_),
    .X(_01474_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net595),
    .S(_05973_),
    .X(_01475_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net528),
    .S(_05973_),
    .X(_01476_));
 sg13g2_nor2_1 _23768_ (.A(_05792_),
    .B(net939),
    .Y(_05975_));
 sg13g2_nand2_2 _23769_ (.Y(_05976_),
    .A(net941),
    .B(_05975_));
 sg13g2_nor3_2 _23770_ (.A(net938),
    .B(_05773_),
    .C(_05976_),
    .Y(_05977_));
 sg13g2_nor2b_1 _23771_ (.A(net394),
    .B_N(_05977_),
    .Y(_05978_));
 sg13g2_buf_1 _23772_ (.A(_05978_),
    .X(_05979_));
 sg13g2_buf_1 _23773_ (.A(_05979_),
    .X(_05980_));
 sg13g2_mux2_1 _23774_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(net335),
    .S(net292),
    .X(_01477_));
 sg13g2_mux2_1 _23775_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(net594),
    .S(net292),
    .X(_01478_));
 sg13g2_mux2_1 _23776_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net717),
    .S(net292),
    .X(_01479_));
 sg13g2_mux2_1 _23777_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(_05942_),
    .S(net292),
    .X(_01480_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(net853),
    .S(net292),
    .X(_01481_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(net852),
    .S(_05980_),
    .X(_01482_));
 sg13g2_mux2_1 _23780_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(net851),
    .S(_05980_),
    .X(_01483_));
 sg13g2_mux2_1 _23781_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(_05943_),
    .S(net292),
    .X(_01484_));
 sg13g2_mux2_1 _23782_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(net933),
    .S(net292),
    .X(_01485_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(_05945_),
    .S(net292),
    .X(_01486_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(_03386_),
    .S(_05979_),
    .X(_01487_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net528),
    .S(_05979_),
    .X(_01488_));
 sg13g2_nor2_1 _23786_ (.A(_05836_),
    .B(_05976_),
    .Y(_05981_));
 sg13g2_buf_1 _23787_ (.A(_05981_),
    .X(_05982_));
 sg13g2_nor2b_1 _23788_ (.A(net394),
    .B_N(_05982_),
    .Y(_05983_));
 sg13g2_buf_1 _23789_ (.A(_05983_),
    .X(_05984_));
 sg13g2_buf_1 _23790_ (.A(_05984_),
    .X(_05985_));
 sg13g2_mux2_1 _23791_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_03398_),
    .S(net291),
    .X(_01489_));
 sg13g2_mux2_1 _23792_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(_03390_),
    .S(net291),
    .X(_01490_));
 sg13g2_mux2_1 _23793_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(_03392_),
    .S(_05985_),
    .X(_01491_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(_02927_),
    .S(net291),
    .X(_01492_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net853),
    .S(net291),
    .X(_01493_));
 sg13g2_mux2_1 _23796_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net852),
    .S(net291),
    .X(_01494_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net851),
    .S(net291),
    .X(_01495_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(net952),
    .S(net291),
    .X(_01496_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net951),
    .S(net291),
    .X(_01497_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net950),
    .S(_05985_),
    .X(_01498_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net595),
    .S(_05984_),
    .X(_01499_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(_03388_),
    .S(_05984_),
    .X(_01500_));
 sg13g2_inv_1 _23803_ (.Y(_05986_),
    .A(_05843_));
 sg13g2_nor3_1 _23804_ (.A(net393),
    .B(_05986_),
    .C(_05870_),
    .Y(_05987_));
 sg13g2_buf_1 _23805_ (.A(_05987_),
    .X(_05988_));
 sg13g2_buf_1 _23806_ (.A(_05988_),
    .X(_05989_));
 sg13g2_mux2_1 _23807_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_03398_),
    .S(net290),
    .X(_01501_));
 sg13g2_mux2_1 _23808_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(net594),
    .S(net290),
    .X(_01502_));
 sg13g2_mux2_1 _23809_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_03392_),
    .S(net290),
    .X(_01503_));
 sg13g2_mux2_1 _23810_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_02927_),
    .S(_05989_),
    .X(_01504_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(_02915_),
    .S(net290),
    .X(_01505_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(_02917_),
    .S(net290),
    .X(_01506_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(_02919_),
    .S(net290),
    .X(_01507_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(_02921_),
    .S(net290),
    .X(_01508_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(_02923_),
    .S(_05989_),
    .X(_01509_));
 sg13g2_mux2_1 _23816_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net950),
    .S(net290),
    .X(_01510_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(net595),
    .S(_05988_),
    .X(_01511_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_03388_),
    .S(_05988_),
    .X(_01512_));
 sg13g2_nand2_1 _23819_ (.Y(_05990_),
    .A(_05843_),
    .B(_05879_));
 sg13g2_buf_2 _23820_ (.A(_05990_),
    .X(_05991_));
 sg13g2_buf_1 _23821_ (.A(_05991_),
    .X(_05992_));
 sg13g2_nand2_1 _23822_ (.Y(_05993_),
    .A(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .B(_05991_));
 sg13g2_o21ai_1 _23823_ (.B1(_05993_),
    .Y(_01513_),
    .A1(net586),
    .A2(net195));
 sg13g2_mux2_1 _23824_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .S(net195),
    .X(_01514_));
 sg13g2_mux2_1 _23825_ (.A0(net639),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .S(net195),
    .X(_01515_));
 sg13g2_nand2_1 _23826_ (.Y(_05994_),
    .A(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .B(_05991_));
 sg13g2_o21ai_1 _23827_ (.B1(_05994_),
    .Y(_01516_),
    .A1(net729),
    .A2(_05992_));
 sg13g2_mux2_1 _23828_ (.A0(net728),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .S(net195),
    .X(_01517_));
 sg13g2_mux2_1 _23829_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .S(net195),
    .X(_01518_));
 sg13g2_mux2_1 _23830_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .S(_05992_),
    .X(_01519_));
 sg13g2_mux2_1 _23831_ (.A0(net850),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .S(net195),
    .X(_01520_));
 sg13g2_mux2_1 _23832_ (.A0(net849),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .S(_05991_),
    .X(_01521_));
 sg13g2_mux2_1 _23833_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .S(_05991_),
    .X(_01522_));
 sg13g2_nand2_1 _23834_ (.Y(_05995_),
    .A(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .B(_05991_));
 sg13g2_o21ai_1 _23835_ (.B1(_05995_),
    .Y(_01523_),
    .A1(net640),
    .A2(net195));
 sg13g2_mux2_1 _23836_ (.A0(net467),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .S(_05991_),
    .X(_01524_));
 sg13g2_and2_1 _23837_ (.A(_05815_),
    .B(_05817_),
    .X(_05996_));
 sg13g2_buf_1 _23838_ (.A(_05996_),
    .X(_05997_));
 sg13g2_nand3_1 _23839_ (.B(_10242_),
    .C(net579),
    .A(net1032),
    .Y(_05998_));
 sg13g2_buf_1 _23840_ (.A(_05998_),
    .X(_05999_));
 sg13g2_nor3_2 _23841_ (.A(net835),
    .B(net941),
    .C(_05999_),
    .Y(_06000_));
 sg13g2_nand2_1 _23842_ (.Y(_06001_),
    .A(_05997_),
    .B(_06000_));
 sg13g2_buf_2 _23843_ (.A(_06001_),
    .X(_06002_));
 sg13g2_buf_1 _23844_ (.A(_06002_),
    .X(_06003_));
 sg13g2_nand2_1 _23845_ (.Y(_06004_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(_06002_));
 sg13g2_o21ai_1 _23846_ (.B1(_06004_),
    .Y(_01525_),
    .A1(net586),
    .A2(net289));
 sg13g2_mux2_1 _23847_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(_06003_),
    .X(_01526_));
 sg13g2_mux2_1 _23848_ (.A0(net639),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .S(_06003_),
    .X(_01527_));
 sg13g2_nand2_1 _23849_ (.Y(_06005_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(_06002_));
 sg13g2_o21ai_1 _23850_ (.B1(_06005_),
    .Y(_01528_),
    .A1(net729),
    .A2(net289));
 sg13g2_mux2_1 _23851_ (.A0(net728),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .S(net289),
    .X(_01529_));
 sg13g2_mux2_1 _23852_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .S(net289),
    .X(_01530_));
 sg13g2_mux2_1 _23853_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .S(net289),
    .X(_01531_));
 sg13g2_mux2_1 _23854_ (.A0(net850),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .S(net289),
    .X(_01532_));
 sg13g2_mux2_1 _23855_ (.A0(net849),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(net289),
    .X(_01533_));
 sg13g2_mux2_1 _23856_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(_06002_),
    .X(_01534_));
 sg13g2_nand2_1 _23857_ (.Y(_06006_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .B(_06002_));
 sg13g2_o21ai_1 _23858_ (.B1(_06006_),
    .Y(_01535_),
    .A1(net640),
    .A2(net289));
 sg13g2_mux2_1 _23859_ (.A0(net467),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(_06002_),
    .X(_01536_));
 sg13g2_and3_1 _23860_ (.X(_06007_),
    .A(net1032),
    .B(_10242_),
    .C(net579));
 sg13g2_buf_1 _23861_ (.A(_06007_),
    .X(_06008_));
 sg13g2_buf_1 _23862_ (.A(_06008_),
    .X(_06009_));
 sg13g2_nand2_1 _23863_ (.Y(_06010_),
    .A(_05829_),
    .B(net392));
 sg13g2_buf_2 _23864_ (.A(_06010_),
    .X(_06011_));
 sg13g2_buf_1 _23865_ (.A(_06011_),
    .X(_06012_));
 sg13g2_nand2_1 _23866_ (.Y(_06013_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(_06011_));
 sg13g2_o21ai_1 _23867_ (.B1(_06013_),
    .Y(_01537_),
    .A1(net586),
    .A2(net288));
 sg13g2_mux2_1 _23868_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(_06012_),
    .X(_01538_));
 sg13g2_mux2_1 _23869_ (.A0(net639),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .S(net288),
    .X(_01539_));
 sg13g2_nand2_1 _23870_ (.Y(_06014_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(_06011_));
 sg13g2_o21ai_1 _23871_ (.B1(_06014_),
    .Y(_01540_),
    .A1(net729),
    .A2(net288));
 sg13g2_mux2_1 _23872_ (.A0(net728),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .S(net288),
    .X(_01541_));
 sg13g2_mux2_1 _23873_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .S(net288),
    .X(_01542_));
 sg13g2_mux2_1 _23874_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .S(net288),
    .X(_01543_));
 sg13g2_mux2_1 _23875_ (.A0(net850),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .S(net288),
    .X(_01544_));
 sg13g2_mux2_1 _23876_ (.A0(net849),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(net288),
    .X(_01545_));
 sg13g2_mux2_1 _23877_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(_06011_),
    .X(_01546_));
 sg13g2_nand2_1 _23878_ (.Y(_06015_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .B(_06011_));
 sg13g2_o21ai_1 _23879_ (.B1(_06015_),
    .Y(_01547_),
    .A1(net640),
    .A2(_06012_));
 sg13g2_mux2_1 _23880_ (.A0(net467),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(_06011_),
    .X(_01548_));
 sg13g2_nand2_1 _23881_ (.Y(_06016_),
    .A(_05838_),
    .B(_06009_));
 sg13g2_buf_2 _23882_ (.A(_06016_),
    .X(_06017_));
 sg13g2_buf_1 _23883_ (.A(_06017_),
    .X(_06018_));
 sg13g2_nand2_1 _23884_ (.Y(_06019_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(_06017_));
 sg13g2_o21ai_1 _23885_ (.B1(_06019_),
    .Y(_01549_),
    .A1(net586),
    .A2(net287));
 sg13g2_mux2_1 _23886_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(_06018_),
    .X(_01550_));
 sg13g2_mux2_1 _23887_ (.A0(net639),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S(net287),
    .X(_01551_));
 sg13g2_nand2_1 _23888_ (.Y(_06020_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(_06017_));
 sg13g2_o21ai_1 _23889_ (.B1(_06020_),
    .Y(_01552_),
    .A1(net729),
    .A2(net287));
 sg13g2_mux2_1 _23890_ (.A0(net728),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S(net287),
    .X(_01553_));
 sg13g2_mux2_1 _23891_ (.A0(net727),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S(net287),
    .X(_01554_));
 sg13g2_mux2_1 _23892_ (.A0(net726),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S(net287),
    .X(_01555_));
 sg13g2_mux2_1 _23893_ (.A0(net850),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S(net287),
    .X(_01556_));
 sg13g2_mux2_1 _23894_ (.A0(net849),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(net287),
    .X(_01557_));
 sg13g2_mux2_1 _23895_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(_06017_),
    .X(_01558_));
 sg13g2_nand2_1 _23896_ (.Y(_06021_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .B(_06017_));
 sg13g2_o21ai_1 _23897_ (.B1(_06021_),
    .Y(_01559_),
    .A1(net640),
    .A2(_06018_));
 sg13g2_mux2_1 _23898_ (.A0(net467),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(_06017_),
    .X(_01560_));
 sg13g2_nor2_1 _23899_ (.A(_05815_),
    .B(_05986_),
    .Y(_06022_));
 sg13g2_nand2_1 _23900_ (.Y(_06023_),
    .A(_06022_),
    .B(_06000_));
 sg13g2_buf_2 _23901_ (.A(_06023_),
    .X(_06024_));
 sg13g2_buf_1 _23902_ (.A(_06024_),
    .X(_06025_));
 sg13g2_nand2_1 _23903_ (.Y(_06026_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(_06024_));
 sg13g2_o21ai_1 _23904_ (.B1(_06026_),
    .Y(_01561_),
    .A1(net586),
    .A2(net286));
 sg13g2_mux2_1 _23905_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(net286),
    .X(_01562_));
 sg13g2_mux2_1 _23906_ (.A0(net639),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .S(_06025_),
    .X(_01563_));
 sg13g2_buf_1 _23907_ (.A(_11715_),
    .X(_06027_));
 sg13g2_nand2_1 _23908_ (.Y(_06028_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(_06024_));
 sg13g2_o21ai_1 _23909_ (.B1(_06028_),
    .Y(_01564_),
    .A1(net706),
    .A2(net286));
 sg13g2_buf_1 _23910_ (.A(net853),
    .X(_06029_));
 sg13g2_mux2_1 _23911_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .S(net286),
    .X(_01565_));
 sg13g2_buf_1 _23912_ (.A(net852),
    .X(_06030_));
 sg13g2_mux2_1 _23913_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .S(net286),
    .X(_01566_));
 sg13g2_buf_1 _23914_ (.A(net851),
    .X(_06031_));
 sg13g2_mux2_1 _23915_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .S(net286),
    .X(_01567_));
 sg13g2_buf_1 _23916_ (.A(net952),
    .X(_06032_));
 sg13g2_mux2_1 _23917_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .S(net286),
    .X(_01568_));
 sg13g2_buf_1 _23918_ (.A(net951),
    .X(_06033_));
 sg13g2_mux2_1 _23919_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(net286),
    .X(_01569_));
 sg13g2_buf_1 _23920_ (.A(net950),
    .X(_06034_));
 sg13g2_mux2_1 _23921_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(_06024_),
    .X(_01570_));
 sg13g2_nand2_1 _23922_ (.Y(_06035_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .B(_06024_));
 sg13g2_o21ai_1 _23923_ (.B1(_06035_),
    .Y(_01571_),
    .A1(net640),
    .A2(_06025_));
 sg13g2_mux2_1 _23924_ (.A0(net467),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(_06024_),
    .X(_01572_));
 sg13g2_nor2_1 _23925_ (.A(_05781_),
    .B(_05999_),
    .Y(_06036_));
 sg13g2_nand2_1 _23926_ (.Y(_06037_),
    .A(_06022_),
    .B(_06036_));
 sg13g2_buf_2 _23927_ (.A(_06037_),
    .X(_06038_));
 sg13g2_buf_1 _23928_ (.A(_06038_),
    .X(_06039_));
 sg13g2_nand2_1 _23929_ (.Y(_06040_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(_06038_));
 sg13g2_o21ai_1 _23930_ (.B1(_06040_),
    .Y(_01573_),
    .A1(net586),
    .A2(net285));
 sg13g2_mux2_1 _23931_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(net285),
    .X(_01574_));
 sg13g2_mux2_1 _23932_ (.A0(net639),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .S(_06039_),
    .X(_01575_));
 sg13g2_nand2_1 _23933_ (.Y(_06041_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(_06038_));
 sg13g2_o21ai_1 _23934_ (.B1(_06041_),
    .Y(_01576_),
    .A1(net706),
    .A2(net285));
 sg13g2_mux2_1 _23935_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .S(net285),
    .X(_01577_));
 sg13g2_mux2_1 _23936_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .S(net285),
    .X(_01578_));
 sg13g2_mux2_1 _23937_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .S(net285),
    .X(_01579_));
 sg13g2_mux2_1 _23938_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .S(net285),
    .X(_01580_));
 sg13g2_mux2_1 _23939_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(net285),
    .X(_01581_));
 sg13g2_mux2_1 _23940_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(_06038_),
    .X(_01582_));
 sg13g2_nand2_1 _23941_ (.Y(_06042_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .B(_06038_));
 sg13g2_o21ai_1 _23942_ (.B1(_06042_),
    .Y(_01583_),
    .A1(net640),
    .A2(_06039_));
 sg13g2_mux2_1 _23943_ (.A0(net467),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(_06038_),
    .X(_01584_));
 sg13g2_buf_1 _23944_ (.A(net637),
    .X(_06043_));
 sg13g2_nor2_1 _23945_ (.A(net709),
    .B(_05999_),
    .Y(_06044_));
 sg13g2_nand2_1 _23946_ (.Y(_06045_),
    .A(_06022_),
    .B(_06044_));
 sg13g2_buf_2 _23947_ (.A(_06045_),
    .X(_06046_));
 sg13g2_buf_1 _23948_ (.A(_06046_),
    .X(_06047_));
 sg13g2_nand2_1 _23949_ (.Y(_06048_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(_06046_));
 sg13g2_o21ai_1 _23950_ (.B1(_06048_),
    .Y(_01585_),
    .A1(net573),
    .A2(net284));
 sg13g2_buf_1 _23951_ (.A(net594),
    .X(_06049_));
 sg13g2_mux2_1 _23952_ (.A0(_06049_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net284),
    .X(_01586_));
 sg13g2_buf_1 _23953_ (.A(net717),
    .X(_06050_));
 sg13g2_mux2_1 _23954_ (.A0(_06050_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .S(net284),
    .X(_01587_));
 sg13g2_nand2_1 _23955_ (.Y(_06051_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(_06046_));
 sg13g2_o21ai_1 _23956_ (.B1(_06051_),
    .Y(_01588_),
    .A1(_06027_),
    .A2(_06047_));
 sg13g2_mux2_1 _23957_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .S(net284),
    .X(_01589_));
 sg13g2_mux2_1 _23958_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .S(net284),
    .X(_01590_));
 sg13g2_mux2_1 _23959_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .S(net284),
    .X(_01591_));
 sg13g2_mux2_1 _23960_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .S(net284),
    .X(_01592_));
 sg13g2_mux2_1 _23961_ (.A0(_06033_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(net284),
    .X(_01593_));
 sg13g2_mux2_1 _23962_ (.A0(_06034_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(_06046_),
    .X(_01594_));
 sg13g2_buf_1 _23963_ (.A(net714),
    .X(_06052_));
 sg13g2_nand2_1 _23964_ (.Y(_06053_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .B(_06046_));
 sg13g2_o21ai_1 _23965_ (.B1(_06053_),
    .Y(_01595_),
    .A1(net633),
    .A2(_06047_));
 sg13g2_buf_1 _23966_ (.A(net528),
    .X(_06054_));
 sg13g2_mux2_1 _23967_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(_06046_),
    .X(_01596_));
 sg13g2_nor2_1 _23968_ (.A(_05791_),
    .B(_05999_),
    .Y(_06055_));
 sg13g2_nand2_1 _23969_ (.Y(_06056_),
    .A(_06022_),
    .B(_06055_));
 sg13g2_buf_2 _23970_ (.A(_06056_),
    .X(_06057_));
 sg13g2_buf_1 _23971_ (.A(_06057_),
    .X(_06058_));
 sg13g2_nand2_1 _23972_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(_06057_));
 sg13g2_o21ai_1 _23973_ (.B1(_06059_),
    .Y(_01597_),
    .A1(_06043_),
    .A2(net283));
 sg13g2_mux2_1 _23974_ (.A0(_06049_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net283),
    .X(_01598_));
 sg13g2_mux2_1 _23975_ (.A0(_06050_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S(net283),
    .X(_01599_));
 sg13g2_nand2_1 _23976_ (.Y(_06060_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(_06057_));
 sg13g2_o21ai_1 _23977_ (.B1(_06060_),
    .Y(_01600_),
    .A1(_06027_),
    .A2(_06058_));
 sg13g2_mux2_1 _23978_ (.A0(_06029_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S(net283),
    .X(_01601_));
 sg13g2_mux2_1 _23979_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S(net283),
    .X(_01602_));
 sg13g2_mux2_1 _23980_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S(net283),
    .X(_01603_));
 sg13g2_mux2_1 _23981_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S(net283),
    .X(_01604_));
 sg13g2_mux2_1 _23982_ (.A0(_06033_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(net283),
    .X(_01605_));
 sg13g2_mux2_1 _23983_ (.A0(_06034_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(_06057_),
    .X(_01606_));
 sg13g2_nand2_1 _23984_ (.Y(_06061_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .B(_06057_));
 sg13g2_o21ai_1 _23985_ (.B1(_06061_),
    .Y(_01607_),
    .A1(_06052_),
    .A2(_06058_));
 sg13g2_mux2_1 _23986_ (.A0(_06054_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(_06057_),
    .X(_01608_));
 sg13g2_nor3_2 _23987_ (.A(net835),
    .B(net941),
    .C(net940),
    .Y(_06062_));
 sg13g2_nand3_1 _23988_ (.B(_06062_),
    .C(net392),
    .A(_05878_),
    .Y(_06063_));
 sg13g2_buf_2 _23989_ (.A(_06063_),
    .X(_06064_));
 sg13g2_buf_1 _23990_ (.A(_06064_),
    .X(_06065_));
 sg13g2_nand2_1 _23991_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(_06064_));
 sg13g2_o21ai_1 _23992_ (.B1(_06066_),
    .Y(_01609_),
    .A1(net573),
    .A2(net282));
 sg13g2_mux2_1 _23993_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(net282),
    .X(_01610_));
 sg13g2_mux2_1 _23994_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .S(net282),
    .X(_01611_));
 sg13g2_nand2_1 _23995_ (.Y(_06067_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(_06064_));
 sg13g2_o21ai_1 _23996_ (.B1(_06067_),
    .Y(_01612_),
    .A1(net706),
    .A2(_06065_));
 sg13g2_mux2_1 _23997_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .S(net282),
    .X(_01613_));
 sg13g2_mux2_1 _23998_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .S(net282),
    .X(_01614_));
 sg13g2_mux2_1 _23999_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .S(net282),
    .X(_01615_));
 sg13g2_mux2_1 _24000_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .S(net282),
    .X(_01616_));
 sg13g2_mux2_1 _24001_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net282),
    .X(_01617_));
 sg13g2_mux2_1 _24002_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(_06064_),
    .X(_01618_));
 sg13g2_nand2_1 _24003_ (.Y(_06068_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .B(_06064_));
 sg13g2_o21ai_1 _24004_ (.B1(_06068_),
    .Y(_01619_),
    .A1(net633),
    .A2(_06065_));
 sg13g2_mux2_1 _24005_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(_06064_),
    .X(_01620_));
 sg13g2_nor3_1 _24006_ (.A(net940),
    .B(_05781_),
    .C(_05999_),
    .Y(_06069_));
 sg13g2_nand2_1 _24007_ (.Y(_06070_),
    .A(_05878_),
    .B(_06069_));
 sg13g2_buf_2 _24008_ (.A(_06070_),
    .X(_06071_));
 sg13g2_buf_1 _24009_ (.A(_06071_),
    .X(_06072_));
 sg13g2_nand2_1 _24010_ (.Y(_06073_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(_06071_));
 sg13g2_o21ai_1 _24011_ (.B1(_06073_),
    .Y(_01621_),
    .A1(net573),
    .A2(net281));
 sg13g2_mux2_1 _24012_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(net281),
    .X(_01622_));
 sg13g2_mux2_1 _24013_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .S(net281),
    .X(_01623_));
 sg13g2_nand2_1 _24014_ (.Y(_06074_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(_06071_));
 sg13g2_o21ai_1 _24015_ (.B1(_06074_),
    .Y(_01624_),
    .A1(net706),
    .A2(_06072_));
 sg13g2_mux2_1 _24016_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .S(net281),
    .X(_01625_));
 sg13g2_mux2_1 _24017_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .S(net281),
    .X(_01626_));
 sg13g2_mux2_1 _24018_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .S(net281),
    .X(_01627_));
 sg13g2_mux2_1 _24019_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .S(net281),
    .X(_01628_));
 sg13g2_mux2_1 _24020_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net281),
    .X(_01629_));
 sg13g2_mux2_1 _24021_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(_06071_),
    .X(_01630_));
 sg13g2_nand2_1 _24022_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .B(_06071_));
 sg13g2_o21ai_1 _24023_ (.B1(_06075_),
    .Y(_01631_),
    .A1(net633),
    .A2(_06072_));
 sg13g2_mux2_1 _24024_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_06071_),
    .X(_01632_));
 sg13g2_nand2_1 _24025_ (.Y(_06076_),
    .A(_05888_),
    .B(net392));
 sg13g2_buf_2 _24026_ (.A(_06076_),
    .X(_06077_));
 sg13g2_buf_1 _24027_ (.A(_06077_),
    .X(_06078_));
 sg13g2_nand2_1 _24028_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24029_ (.B1(_06079_),
    .Y(_01633_),
    .A1(net573),
    .A2(net280));
 sg13g2_mux2_1 _24030_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(net280),
    .X(_01634_));
 sg13g2_mux2_1 _24031_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .S(net280),
    .X(_01635_));
 sg13g2_nand2_1 _24032_ (.Y(_06080_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24033_ (.B1(_06080_),
    .Y(_01636_),
    .A1(net706),
    .A2(_06078_));
 sg13g2_mux2_1 _24034_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .S(net280),
    .X(_01637_));
 sg13g2_mux2_1 _24035_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .S(net280),
    .X(_01638_));
 sg13g2_mux2_1 _24036_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .S(net280),
    .X(_01639_));
 sg13g2_mux2_1 _24037_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .S(net280),
    .X(_01640_));
 sg13g2_mux2_1 _24038_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net280),
    .X(_01641_));
 sg13g2_mux2_1 _24039_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(_06077_),
    .X(_01642_));
 sg13g2_nand2_1 _24040_ (.Y(_06081_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .B(_06077_));
 sg13g2_o21ai_1 _24041_ (.B1(_06081_),
    .Y(_01643_),
    .A1(net633),
    .A2(_06078_));
 sg13g2_mux2_1 _24042_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_06077_),
    .X(_01644_));
 sg13g2_nand2_1 _24043_ (.Y(_06082_),
    .A(_05894_),
    .B(net392));
 sg13g2_buf_2 _24044_ (.A(_06082_),
    .X(_06083_));
 sg13g2_buf_1 _24045_ (.A(_06083_),
    .X(_06084_));
 sg13g2_nand2_1 _24046_ (.Y(_06085_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(_06083_));
 sg13g2_o21ai_1 _24047_ (.B1(_06085_),
    .Y(_01645_),
    .A1(net573),
    .A2(net279));
 sg13g2_mux2_1 _24048_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(net279),
    .X(_01646_));
 sg13g2_mux2_1 _24049_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S(net279),
    .X(_01647_));
 sg13g2_nand2_1 _24050_ (.Y(_06086_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(_06083_));
 sg13g2_o21ai_1 _24051_ (.B1(_06086_),
    .Y(_01648_),
    .A1(net706),
    .A2(_06084_));
 sg13g2_mux2_1 _24052_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S(net279),
    .X(_01649_));
 sg13g2_mux2_1 _24053_ (.A0(net704),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S(net279),
    .X(_01650_));
 sg13g2_mux2_1 _24054_ (.A0(net703),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S(net279),
    .X(_01651_));
 sg13g2_mux2_1 _24055_ (.A0(net827),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S(net279),
    .X(_01652_));
 sg13g2_mux2_1 _24056_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net279),
    .X(_01653_));
 sg13g2_mux2_1 _24057_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(_06083_),
    .X(_01654_));
 sg13g2_nand2_1 _24058_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .B(_06083_));
 sg13g2_o21ai_1 _24059_ (.B1(_06087_),
    .Y(_01655_),
    .A1(net633),
    .A2(_06084_));
 sg13g2_mux2_1 _24060_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_06083_),
    .X(_01656_));
 sg13g2_nand2_1 _24061_ (.Y(_06088_),
    .A(_05997_),
    .B(_06036_));
 sg13g2_buf_2 _24062_ (.A(_06088_),
    .X(_06089_));
 sg13g2_buf_1 _24063_ (.A(_06089_),
    .X(_06090_));
 sg13g2_nand2_1 _24064_ (.Y(_06091_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(_06089_));
 sg13g2_o21ai_1 _24065_ (.B1(_06091_),
    .Y(_01657_),
    .A1(_06043_),
    .A2(net278));
 sg13g2_mux2_1 _24066_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(net278),
    .X(_01658_));
 sg13g2_mux2_1 _24067_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .S(net278),
    .X(_01659_));
 sg13g2_nand2_1 _24068_ (.Y(_06092_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(_06089_));
 sg13g2_o21ai_1 _24069_ (.B1(_06092_),
    .Y(_01660_),
    .A1(net706),
    .A2(_06090_));
 sg13g2_mux2_1 _24070_ (.A0(_06029_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .S(net278),
    .X(_01661_));
 sg13g2_mux2_1 _24071_ (.A0(_06030_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .S(net278),
    .X(_01662_));
 sg13g2_mux2_1 _24072_ (.A0(_06031_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .S(net278),
    .X(_01663_));
 sg13g2_mux2_1 _24073_ (.A0(_06032_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .S(net278),
    .X(_01664_));
 sg13g2_mux2_1 _24074_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(net278),
    .X(_01665_));
 sg13g2_mux2_1 _24075_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(_06089_),
    .X(_01666_));
 sg13g2_nand2_1 _24076_ (.Y(_06093_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .B(_06089_));
 sg13g2_o21ai_1 _24077_ (.B1(_06093_),
    .Y(_01667_),
    .A1(_06052_),
    .A2(_06090_));
 sg13g2_mux2_1 _24078_ (.A0(_06054_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(_06089_),
    .X(_01668_));
 sg13g2_nor2_1 _24079_ (.A(_05815_),
    .B(_05867_),
    .Y(_06094_));
 sg13g2_nand2_1 _24080_ (.Y(_06095_),
    .A(_06094_),
    .B(_06000_));
 sg13g2_buf_2 _24081_ (.A(_06095_),
    .X(_06096_));
 sg13g2_buf_1 _24082_ (.A(_06096_),
    .X(_06097_));
 sg13g2_nand2_1 _24083_ (.Y(_06098_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(_06096_));
 sg13g2_o21ai_1 _24084_ (.B1(_06098_),
    .Y(_01669_),
    .A1(net573),
    .A2(net277));
 sg13g2_mux2_1 _24085_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(net277),
    .X(_01670_));
 sg13g2_mux2_1 _24086_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .S(net277),
    .X(_01671_));
 sg13g2_nand2_1 _24087_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(_06096_));
 sg13g2_o21ai_1 _24088_ (.B1(_06099_),
    .Y(_01672_),
    .A1(net706),
    .A2(_06097_));
 sg13g2_mux2_1 _24089_ (.A0(net705),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .S(net277),
    .X(_01673_));
 sg13g2_mux2_1 _24090_ (.A0(_06030_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .S(net277),
    .X(_01674_));
 sg13g2_mux2_1 _24091_ (.A0(_06031_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .S(net277),
    .X(_01675_));
 sg13g2_mux2_1 _24092_ (.A0(_06032_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .S(net277),
    .X(_01676_));
 sg13g2_mux2_1 _24093_ (.A0(net826),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(net277),
    .X(_01677_));
 sg13g2_mux2_1 _24094_ (.A0(net825),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(_06096_),
    .X(_01678_));
 sg13g2_nand2_1 _24095_ (.Y(_06100_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .B(_06096_));
 sg13g2_o21ai_1 _24096_ (.B1(_06100_),
    .Y(_01679_),
    .A1(net633),
    .A2(_06097_));
 sg13g2_mux2_1 _24097_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(_06096_),
    .X(_01680_));
 sg13g2_nand2_1 _24098_ (.Y(_06101_),
    .A(_06094_),
    .B(_06036_));
 sg13g2_buf_2 _24099_ (.A(_06101_),
    .X(_06102_));
 sg13g2_buf_1 _24100_ (.A(_06102_),
    .X(_06103_));
 sg13g2_nand2_1 _24101_ (.Y(_06104_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(_06102_));
 sg13g2_o21ai_1 _24102_ (.B1(_06104_),
    .Y(_01681_),
    .A1(net573),
    .A2(net276));
 sg13g2_mux2_1 _24103_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(net276),
    .X(_01682_));
 sg13g2_mux2_1 _24104_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .S(net276),
    .X(_01683_));
 sg13g2_buf_1 _24105_ (.A(_11715_),
    .X(_06105_));
 sg13g2_nand2_1 _24106_ (.Y(_06106_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(_06102_));
 sg13g2_o21ai_1 _24107_ (.B1(_06106_),
    .Y(_01684_),
    .A1(net702),
    .A2(_06103_));
 sg13g2_buf_1 _24108_ (.A(net853),
    .X(_06107_));
 sg13g2_mux2_1 _24109_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .S(net276),
    .X(_01685_));
 sg13g2_buf_1 _24110_ (.A(net852),
    .X(_06108_));
 sg13g2_mux2_1 _24111_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .S(net276),
    .X(_01686_));
 sg13g2_buf_1 _24112_ (.A(net851),
    .X(_06109_));
 sg13g2_mux2_1 _24113_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .S(net276),
    .X(_01687_));
 sg13g2_buf_1 _24114_ (.A(net952),
    .X(_06110_));
 sg13g2_mux2_1 _24115_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .S(net276),
    .X(_01688_));
 sg13g2_buf_1 _24116_ (.A(net951),
    .X(_06111_));
 sg13g2_mux2_1 _24117_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(net276),
    .X(_01689_));
 sg13g2_buf_1 _24118_ (.A(net950),
    .X(_06112_));
 sg13g2_mux2_1 _24119_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(_06102_),
    .X(_01690_));
 sg13g2_nand2_1 _24120_ (.Y(_06113_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .B(_06102_));
 sg13g2_o21ai_1 _24121_ (.B1(_06113_),
    .Y(_01691_),
    .A1(net633),
    .A2(_06103_));
 sg13g2_mux2_1 _24122_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(_06102_),
    .X(_01692_));
 sg13g2_nand2_1 _24123_ (.Y(_06114_),
    .A(_06094_),
    .B(_06044_));
 sg13g2_buf_2 _24124_ (.A(_06114_),
    .X(_06115_));
 sg13g2_buf_1 _24125_ (.A(_06115_),
    .X(_06116_));
 sg13g2_nand2_1 _24126_ (.Y(_06117_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(_06115_));
 sg13g2_o21ai_1 _24127_ (.B1(_06117_),
    .Y(_01693_),
    .A1(net573),
    .A2(net275));
 sg13g2_mux2_1 _24128_ (.A0(net508),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(net275),
    .X(_01694_));
 sg13g2_mux2_1 _24129_ (.A0(net634),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .S(net275),
    .X(_01695_));
 sg13g2_nand2_1 _24130_ (.Y(_06118_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(_06115_));
 sg13g2_o21ai_1 _24131_ (.B1(_06118_),
    .Y(_01696_),
    .A1(_06105_),
    .A2(_06116_));
 sg13g2_mux2_1 _24132_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .S(net275),
    .X(_01697_));
 sg13g2_mux2_1 _24133_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .S(net275),
    .X(_01698_));
 sg13g2_mux2_1 _24134_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .S(net275),
    .X(_01699_));
 sg13g2_mux2_1 _24135_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .S(net275),
    .X(_01700_));
 sg13g2_mux2_1 _24136_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(net275),
    .X(_01701_));
 sg13g2_mux2_1 _24137_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(_06115_),
    .X(_01702_));
 sg13g2_nand2_1 _24138_ (.Y(_06119_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .B(_06115_));
 sg13g2_o21ai_1 _24139_ (.B1(_06119_),
    .Y(_01703_),
    .A1(net633),
    .A2(_06116_));
 sg13g2_mux2_1 _24140_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(_06115_),
    .X(_01704_));
 sg13g2_buf_1 _24141_ (.A(net712),
    .X(_06120_));
 sg13g2_nand2_1 _24142_ (.Y(_06121_),
    .A(_06094_),
    .B(_06055_));
 sg13g2_buf_2 _24143_ (.A(_06121_),
    .X(_06122_));
 sg13g2_buf_1 _24144_ (.A(_06122_),
    .X(_06123_));
 sg13g2_nand2_1 _24145_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24146_ (.B1(_06124_),
    .Y(_01705_),
    .A1(net632),
    .A2(net274));
 sg13g2_buf_1 _24147_ (.A(net594),
    .X(_06125_));
 sg13g2_mux2_1 _24148_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(net274),
    .X(_01706_));
 sg13g2_buf_1 _24149_ (.A(net717),
    .X(_06126_));
 sg13g2_mux2_1 _24150_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S(net274),
    .X(_01707_));
 sg13g2_nand2_1 _24151_ (.Y(_06127_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24152_ (.B1(_06127_),
    .Y(_01708_),
    .A1(_06105_),
    .A2(_06123_));
 sg13g2_mux2_1 _24153_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S(net274),
    .X(_01709_));
 sg13g2_mux2_1 _24154_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S(net274),
    .X(_01710_));
 sg13g2_mux2_1 _24155_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S(net274),
    .X(_01711_));
 sg13g2_mux2_1 _24156_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S(net274),
    .X(_01712_));
 sg13g2_mux2_1 _24157_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(net274),
    .X(_01713_));
 sg13g2_mux2_1 _24158_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(_06122_),
    .X(_01714_));
 sg13g2_buf_1 _24159_ (.A(net714),
    .X(_06128_));
 sg13g2_nand2_1 _24160_ (.Y(_06129_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .B(_06122_));
 sg13g2_o21ai_1 _24161_ (.B1(_06129_),
    .Y(_01715_),
    .A1(net630),
    .A2(_06123_));
 sg13g2_buf_1 _24162_ (.A(net528),
    .X(_06130_));
 sg13g2_mux2_1 _24163_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(_06122_),
    .X(_01716_));
 sg13g2_nand4_1 _24164_ (.B(net834),
    .C(_06062_),
    .A(net938),
    .Y(_06131_),
    .D(_06008_));
 sg13g2_buf_2 _24165_ (.A(_06131_),
    .X(_06132_));
 sg13g2_buf_1 _24166_ (.A(_06132_),
    .X(_06133_));
 sg13g2_nand2_1 _24167_ (.Y(_06134_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24168_ (.B1(_06134_),
    .Y(_01717_),
    .A1(net632),
    .A2(net329));
 sg13g2_mux2_1 _24169_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(net329),
    .X(_01718_));
 sg13g2_mux2_1 _24170_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .S(net329),
    .X(_01719_));
 sg13g2_nand2_1 _24171_ (.Y(_06135_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24172_ (.B1(_06135_),
    .Y(_01720_),
    .A1(net702),
    .A2(net329));
 sg13g2_mux2_1 _24173_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .S(_06133_),
    .X(_01721_));
 sg13g2_mux2_1 _24174_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .S(net329),
    .X(_01722_));
 sg13g2_mux2_1 _24175_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .S(net329),
    .X(_01723_));
 sg13g2_mux2_1 _24176_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .S(net329),
    .X(_01724_));
 sg13g2_mux2_1 _24177_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(net329),
    .X(_01725_));
 sg13g2_mux2_1 _24178_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(_06132_),
    .X(_01726_));
 sg13g2_nand2_1 _24179_ (.Y(_06136_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24180_ (.B1(_06136_),
    .Y(_01727_),
    .A1(net630),
    .A2(_06133_));
 sg13g2_mux2_1 _24181_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(_06132_),
    .X(_01728_));
 sg13g2_nand2b_1 _24182_ (.Y(_06137_),
    .B(_06069_),
    .A_N(_05919_));
 sg13g2_buf_2 _24183_ (.A(_06137_),
    .X(_06138_));
 sg13g2_buf_1 _24184_ (.A(_06138_),
    .X(_06139_));
 sg13g2_nand2_1 _24185_ (.Y(_06140_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(_06138_));
 sg13g2_o21ai_1 _24186_ (.B1(_06140_),
    .Y(_01729_),
    .A1(net632),
    .A2(net273));
 sg13g2_mux2_1 _24187_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(net273),
    .X(_01730_));
 sg13g2_mux2_1 _24188_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .S(net273),
    .X(_01731_));
 sg13g2_nand2_1 _24189_ (.Y(_06141_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(_06138_));
 sg13g2_o21ai_1 _24190_ (.B1(_06141_),
    .Y(_01732_),
    .A1(net702),
    .A2(net273));
 sg13g2_mux2_1 _24191_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .S(_06139_),
    .X(_01733_));
 sg13g2_mux2_1 _24192_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .S(net273),
    .X(_01734_));
 sg13g2_mux2_1 _24193_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .S(net273),
    .X(_01735_));
 sg13g2_mux2_1 _24194_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .S(net273),
    .X(_01736_));
 sg13g2_mux2_1 _24195_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(net273),
    .X(_01737_));
 sg13g2_mux2_1 _24196_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(_06138_),
    .X(_01738_));
 sg13g2_nand2_1 _24197_ (.Y(_06142_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .B(_06138_));
 sg13g2_o21ai_1 _24198_ (.B1(_06142_),
    .Y(_01739_),
    .A1(net630),
    .A2(_06139_));
 sg13g2_mux2_1 _24199_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(_06138_),
    .X(_01740_));
 sg13g2_nand2_1 _24200_ (.Y(_06143_),
    .A(_05930_),
    .B(net392));
 sg13g2_buf_2 _24201_ (.A(_06143_),
    .X(_06144_));
 sg13g2_buf_1 _24202_ (.A(_06144_),
    .X(_06145_));
 sg13g2_nand2_1 _24203_ (.Y(_06146_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24204_ (.B1(_06146_),
    .Y(_01741_),
    .A1(net632),
    .A2(net272));
 sg13g2_mux2_1 _24205_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(net272),
    .X(_01742_));
 sg13g2_mux2_1 _24206_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .S(net272),
    .X(_01743_));
 sg13g2_nand2_1 _24207_ (.Y(_06147_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24208_ (.B1(_06147_),
    .Y(_01744_),
    .A1(net702),
    .A2(net272));
 sg13g2_mux2_1 _24209_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .S(_06145_),
    .X(_01745_));
 sg13g2_mux2_1 _24210_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .S(net272),
    .X(_01746_));
 sg13g2_mux2_1 _24211_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .S(net272),
    .X(_01747_));
 sg13g2_mux2_1 _24212_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .S(net272),
    .X(_01748_));
 sg13g2_mux2_1 _24213_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(net272),
    .X(_01749_));
 sg13g2_mux2_1 _24214_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(_06144_),
    .X(_01750_));
 sg13g2_nand2_1 _24215_ (.Y(_06148_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24216_ (.B1(_06148_),
    .Y(_01751_),
    .A1(net630),
    .A2(_06145_));
 sg13g2_mux2_1 _24217_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(_06144_),
    .X(_01752_));
 sg13g2_nand2_1 _24218_ (.Y(_06149_),
    .A(_05938_),
    .B(net392));
 sg13g2_buf_2 _24219_ (.A(_06149_),
    .X(_06150_));
 sg13g2_buf_1 _24220_ (.A(_06150_),
    .X(_06151_));
 sg13g2_nand2_1 _24221_ (.Y(_06152_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24222_ (.B1(_06152_),
    .Y(_01753_),
    .A1(_06120_),
    .A2(net271));
 sg13g2_mux2_1 _24223_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net271),
    .X(_01754_));
 sg13g2_mux2_1 _24224_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S(net271),
    .X(_01755_));
 sg13g2_nand2_1 _24225_ (.Y(_06153_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24226_ (.B1(_06153_),
    .Y(_01756_),
    .A1(net702),
    .A2(net271));
 sg13g2_mux2_1 _24227_ (.A0(_06107_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S(_06151_),
    .X(_01757_));
 sg13g2_mux2_1 _24228_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S(net271),
    .X(_01758_));
 sg13g2_mux2_1 _24229_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S(net271),
    .X(_01759_));
 sg13g2_mux2_1 _24230_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S(net271),
    .X(_01760_));
 sg13g2_mux2_1 _24231_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(net271),
    .X(_01761_));
 sg13g2_mux2_1 _24232_ (.A0(_06112_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(_06150_),
    .X(_01762_));
 sg13g2_nand2_1 _24233_ (.Y(_06154_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .B(_06150_));
 sg13g2_o21ai_1 _24234_ (.B1(_06154_),
    .Y(_01763_),
    .A1(_06128_),
    .A2(_06151_));
 sg13g2_mux2_1 _24235_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(_06150_),
    .X(_01764_));
 sg13g2_nor2_1 _24236_ (.A(_05815_),
    .B(_05919_),
    .Y(_06155_));
 sg13g2_nand2_1 _24237_ (.Y(_06156_),
    .A(_06155_),
    .B(_06000_));
 sg13g2_buf_2 _24238_ (.A(_06156_),
    .X(_06157_));
 sg13g2_buf_1 _24239_ (.A(_06157_),
    .X(_06158_));
 sg13g2_nand2_1 _24240_ (.Y(_06159_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24241_ (.B1(_06159_),
    .Y(_01765_),
    .A1(net632),
    .A2(net270));
 sg13g2_mux2_1 _24242_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(net270),
    .X(_01766_));
 sg13g2_mux2_1 _24243_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .S(net270),
    .X(_01767_));
 sg13g2_nand2_1 _24244_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24245_ (.B1(_06160_),
    .Y(_01768_),
    .A1(net702),
    .A2(_06158_));
 sg13g2_mux2_1 _24246_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .S(net270),
    .X(_01769_));
 sg13g2_mux2_1 _24247_ (.A0(_06108_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .S(net270),
    .X(_01770_));
 sg13g2_mux2_1 _24248_ (.A0(_06109_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .S(net270),
    .X(_01771_));
 sg13g2_mux2_1 _24249_ (.A0(_06110_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .S(net270),
    .X(_01772_));
 sg13g2_mux2_1 _24250_ (.A0(_06111_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(net270),
    .X(_01773_));
 sg13g2_mux2_1 _24251_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(_06157_),
    .X(_01774_));
 sg13g2_nand2_1 _24252_ (.Y(_06161_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .B(_06157_));
 sg13g2_o21ai_1 _24253_ (.B1(_06161_),
    .Y(_01775_),
    .A1(net630),
    .A2(_06158_));
 sg13g2_mux2_1 _24254_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(_06157_),
    .X(_01776_));
 sg13g2_nand2_1 _24255_ (.Y(_06162_),
    .A(_06155_),
    .B(_06036_));
 sg13g2_buf_2 _24256_ (.A(_06162_),
    .X(_06163_));
 sg13g2_buf_1 _24257_ (.A(_06163_),
    .X(_06164_));
 sg13g2_nand2_1 _24258_ (.Y(_06165_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(_06163_));
 sg13g2_o21ai_1 _24259_ (.B1(_06165_),
    .Y(_01777_),
    .A1(net632),
    .A2(net269));
 sg13g2_mux2_1 _24260_ (.A0(_06125_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(net269),
    .X(_01778_));
 sg13g2_mux2_1 _24261_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .S(net269),
    .X(_01779_));
 sg13g2_nand2_1 _24262_ (.Y(_06166_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(_06163_));
 sg13g2_o21ai_1 _24263_ (.B1(_06166_),
    .Y(_01780_),
    .A1(net702),
    .A2(_06164_));
 sg13g2_mux2_1 _24264_ (.A0(net701),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .S(net269),
    .X(_01781_));
 sg13g2_mux2_1 _24265_ (.A0(net700),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .S(net269),
    .X(_01782_));
 sg13g2_mux2_1 _24266_ (.A0(net699),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .S(net269),
    .X(_01783_));
 sg13g2_mux2_1 _24267_ (.A0(net824),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .S(net269),
    .X(_01784_));
 sg13g2_mux2_1 _24268_ (.A0(_06111_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(net269),
    .X(_01785_));
 sg13g2_mux2_1 _24269_ (.A0(net822),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(_06163_),
    .X(_01786_));
 sg13g2_nand2_1 _24270_ (.Y(_06167_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .B(_06163_));
 sg13g2_o21ai_1 _24271_ (.B1(_06167_),
    .Y(_01787_),
    .A1(net630),
    .A2(_06164_));
 sg13g2_mux2_1 _24272_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(_06163_),
    .X(_01788_));
 sg13g2_nand2_1 _24273_ (.Y(_06168_),
    .A(_05997_),
    .B(_06044_));
 sg13g2_buf_2 _24274_ (.A(_06168_),
    .X(_06169_));
 sg13g2_buf_1 _24275_ (.A(_06169_),
    .X(_06170_));
 sg13g2_nand2_1 _24276_ (.Y(_06171_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(_06169_));
 sg13g2_o21ai_1 _24277_ (.B1(_06171_),
    .Y(_01789_),
    .A1(_06120_),
    .A2(net268));
 sg13g2_mux2_1 _24278_ (.A0(_06125_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(net268),
    .X(_01790_));
 sg13g2_mux2_1 _24279_ (.A0(net631),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .S(net268),
    .X(_01791_));
 sg13g2_nand2_1 _24280_ (.Y(_06172_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(_06169_));
 sg13g2_o21ai_1 _24281_ (.B1(_06172_),
    .Y(_01792_),
    .A1(net702),
    .A2(_06170_));
 sg13g2_mux2_1 _24282_ (.A0(_06107_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .S(net268),
    .X(_01793_));
 sg13g2_mux2_1 _24283_ (.A0(_06108_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .S(net268),
    .X(_01794_));
 sg13g2_mux2_1 _24284_ (.A0(_06109_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .S(net268),
    .X(_01795_));
 sg13g2_mux2_1 _24285_ (.A0(_06110_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .S(net268),
    .X(_01796_));
 sg13g2_mux2_1 _24286_ (.A0(net823),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(net268),
    .X(_01797_));
 sg13g2_mux2_1 _24287_ (.A0(_06112_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(_06169_),
    .X(_01798_));
 sg13g2_nand2_1 _24288_ (.Y(_06173_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .B(_06169_));
 sg13g2_o21ai_1 _24289_ (.B1(_06173_),
    .Y(_01799_),
    .A1(_06128_),
    .A2(_06170_));
 sg13g2_mux2_1 _24290_ (.A0(_06130_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(_06169_),
    .X(_01800_));
 sg13g2_nand2_1 _24291_ (.Y(_06174_),
    .A(_06155_),
    .B(_06044_));
 sg13g2_buf_2 _24292_ (.A(_06174_),
    .X(_06175_));
 sg13g2_buf_1 _24293_ (.A(_06175_),
    .X(_06176_));
 sg13g2_nand2_1 _24294_ (.Y(_06177_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(_06175_));
 sg13g2_o21ai_1 _24295_ (.B1(_06177_),
    .Y(_01801_),
    .A1(net632),
    .A2(net267));
 sg13g2_mux2_1 _24296_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(net267),
    .X(_01802_));
 sg13g2_mux2_1 _24297_ (.A0(_06126_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .S(_06176_),
    .X(_01803_));
 sg13g2_buf_1 _24298_ (.A(net865),
    .X(_06178_));
 sg13g2_nand2_1 _24299_ (.Y(_06179_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(_06175_));
 sg13g2_o21ai_1 _24300_ (.B1(_06179_),
    .Y(_01804_),
    .A1(net698),
    .A2(_06176_));
 sg13g2_mux2_1 _24301_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .S(net267),
    .X(_01805_));
 sg13g2_mux2_1 _24302_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .S(net267),
    .X(_01806_));
 sg13g2_mux2_1 _24303_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .S(net267),
    .X(_01807_));
 sg13g2_mux2_1 _24304_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .S(net267),
    .X(_01808_));
 sg13g2_mux2_1 _24305_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(net267),
    .X(_01809_));
 sg13g2_mux2_1 _24306_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(_06175_),
    .X(_01810_));
 sg13g2_nand2_1 _24307_ (.Y(_06180_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .B(_06175_));
 sg13g2_o21ai_1 _24308_ (.B1(_06180_),
    .Y(_01811_),
    .A1(net630),
    .A2(net267));
 sg13g2_mux2_1 _24309_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(_06175_),
    .X(_01812_));
 sg13g2_nand2_1 _24310_ (.Y(_06181_),
    .A(_06155_),
    .B(_06055_));
 sg13g2_buf_2 _24311_ (.A(_06181_),
    .X(_06182_));
 sg13g2_buf_1 _24312_ (.A(_06182_),
    .X(_06183_));
 sg13g2_nand2_1 _24313_ (.Y(_06184_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(_06182_));
 sg13g2_o21ai_1 _24314_ (.B1(_06184_),
    .Y(_01813_),
    .A1(net632),
    .A2(net266));
 sg13g2_mux2_1 _24315_ (.A0(net507),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(net266),
    .X(_01814_));
 sg13g2_mux2_1 _24316_ (.A0(_06126_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S(_06183_),
    .X(_01815_));
 sg13g2_nand2_1 _24317_ (.Y(_06185_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(_06182_));
 sg13g2_o21ai_1 _24318_ (.B1(_06185_),
    .Y(_01816_),
    .A1(net698),
    .A2(_06183_));
 sg13g2_mux2_1 _24319_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S(net266),
    .X(_01817_));
 sg13g2_mux2_1 _24320_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S(net266),
    .X(_01818_));
 sg13g2_mux2_1 _24321_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S(net266),
    .X(_01819_));
 sg13g2_mux2_1 _24322_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S(net266),
    .X(_01820_));
 sg13g2_mux2_1 _24323_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(net266),
    .X(_01821_));
 sg13g2_mux2_1 _24324_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(_06182_),
    .X(_01822_));
 sg13g2_nand2_1 _24325_ (.Y(_06186_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .B(_06182_));
 sg13g2_o21ai_1 _24326_ (.B1(_06186_),
    .Y(_01823_),
    .A1(net630),
    .A2(net266));
 sg13g2_mux2_1 _24327_ (.A0(_06130_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(_06182_),
    .X(_01824_));
 sg13g2_nand2_1 _24328_ (.Y(_06187_),
    .A(_05997_),
    .B(_06055_));
 sg13g2_buf_2 _24329_ (.A(_06187_),
    .X(_06188_));
 sg13g2_buf_1 _24330_ (.A(_06188_),
    .X(_06189_));
 sg13g2_nand2_1 _24331_ (.Y(_06190_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(_06188_));
 sg13g2_o21ai_1 _24332_ (.B1(_06190_),
    .Y(_01825_),
    .A1(net637),
    .A2(_06189_));
 sg13g2_mux2_1 _24333_ (.A0(net527),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(net265),
    .X(_01826_));
 sg13g2_mux2_1 _24334_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S(_06189_),
    .X(_01827_));
 sg13g2_nand2_1 _24335_ (.Y(_06191_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(_06188_));
 sg13g2_o21ai_1 _24336_ (.B1(_06191_),
    .Y(_01828_),
    .A1(_06178_),
    .A2(net265));
 sg13g2_mux2_1 _24337_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S(net265),
    .X(_01829_));
 sg13g2_mux2_1 _24338_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S(net265),
    .X(_01830_));
 sg13g2_mux2_1 _24339_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S(net265),
    .X(_01831_));
 sg13g2_mux2_1 _24340_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S(net265),
    .X(_01832_));
 sg13g2_mux2_1 _24341_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(net265),
    .X(_01833_));
 sg13g2_mux2_1 _24342_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(_06188_),
    .X(_01834_));
 sg13g2_nand2_1 _24343_ (.Y(_06192_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .B(_06188_));
 sg13g2_o21ai_1 _24344_ (.B1(_06192_),
    .Y(_01835_),
    .A1(net714),
    .A2(net265));
 sg13g2_mux2_1 _24345_ (.A0(net470),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(_06188_),
    .X(_01836_));
 sg13g2_nand3_1 _24346_ (.B(_05975_),
    .C(_06000_),
    .A(_05835_),
    .Y(_06193_));
 sg13g2_buf_2 _24347_ (.A(_06193_),
    .X(_06194_));
 sg13g2_buf_1 _24348_ (.A(_06194_),
    .X(_06195_));
 sg13g2_nand2_1 _24349_ (.Y(_06196_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24350_ (.B1(_06196_),
    .Y(_01837_),
    .A1(net637),
    .A2(_06195_));
 sg13g2_mux2_1 _24351_ (.A0(net527),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net264),
    .X(_01838_));
 sg13g2_mux2_1 _24352_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .S(_06195_),
    .X(_01839_));
 sg13g2_nand2_1 _24353_ (.Y(_06197_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24354_ (.B1(_06197_),
    .Y(_01840_),
    .A1(net698),
    .A2(net264));
 sg13g2_mux2_1 _24355_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .S(net264),
    .X(_01841_));
 sg13g2_mux2_1 _24356_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .S(net264),
    .X(_01842_));
 sg13g2_mux2_1 _24357_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .S(net264),
    .X(_01843_));
 sg13g2_mux2_1 _24358_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .S(net264),
    .X(_01844_));
 sg13g2_mux2_1 _24359_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(net264),
    .X(_01845_));
 sg13g2_mux2_1 _24360_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(_06194_),
    .X(_01846_));
 sg13g2_nand2_1 _24361_ (.Y(_06198_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .B(_06194_));
 sg13g2_o21ai_1 _24362_ (.B1(_06198_),
    .Y(_01847_),
    .A1(net714),
    .A2(net264));
 sg13g2_mux2_1 _24363_ (.A0(net470),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(_06194_),
    .X(_01848_));
 sg13g2_nand2_1 _24364_ (.Y(_06199_),
    .A(_05971_),
    .B(net392));
 sg13g2_buf_2 _24365_ (.A(_06199_),
    .X(_06200_));
 sg13g2_buf_1 _24366_ (.A(_06200_),
    .X(_06201_));
 sg13g2_nand2_1 _24367_ (.Y(_06202_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(_06200_));
 sg13g2_o21ai_1 _24368_ (.B1(_06202_),
    .Y(_01849_),
    .A1(net637),
    .A2(_06201_));
 sg13g2_mux2_1 _24369_ (.A0(net527),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net263),
    .X(_01850_));
 sg13g2_mux2_1 _24370_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .S(_06201_),
    .X(_01851_));
 sg13g2_nand2_1 _24371_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(_06200_));
 sg13g2_o21ai_1 _24372_ (.B1(_06203_),
    .Y(_01852_),
    .A1(net698),
    .A2(net263));
 sg13g2_mux2_1 _24373_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .S(net263),
    .X(_01853_));
 sg13g2_mux2_1 _24374_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .S(net263),
    .X(_01854_));
 sg13g2_mux2_1 _24375_ (.A0(_02933_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .S(net263),
    .X(_01855_));
 sg13g2_mux2_1 _24376_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .S(net263),
    .X(_01856_));
 sg13g2_mux2_1 _24377_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(net263),
    .X(_01857_));
 sg13g2_mux2_1 _24378_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(_06200_),
    .X(_01858_));
 sg13g2_nand2_1 _24379_ (.Y(_06204_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .B(_06200_));
 sg13g2_o21ai_1 _24380_ (.B1(_06204_),
    .Y(_01859_),
    .A1(net714),
    .A2(net263));
 sg13g2_mux2_1 _24381_ (.A0(net470),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(_06200_),
    .X(_01860_));
 sg13g2_nand2_1 _24382_ (.Y(_06205_),
    .A(_05977_),
    .B(_06009_));
 sg13g2_buf_2 _24383_ (.A(_06205_),
    .X(_06206_));
 sg13g2_buf_1 _24384_ (.A(_06206_),
    .X(_06207_));
 sg13g2_nand2_1 _24385_ (.Y(_06208_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24386_ (.B1(_06208_),
    .Y(_01861_),
    .A1(net637),
    .A2(_06207_));
 sg13g2_mux2_1 _24387_ (.A0(net527),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net262),
    .X(_01862_));
 sg13g2_mux2_1 _24388_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .S(_06207_),
    .X(_01863_));
 sg13g2_nand2_1 _24389_ (.Y(_06209_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24390_ (.B1(_06209_),
    .Y(_01864_),
    .A1(net698),
    .A2(net262));
 sg13g2_mux2_1 _24391_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .S(net262),
    .X(_01865_));
 sg13g2_mux2_1 _24392_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .S(net262),
    .X(_01866_));
 sg13g2_mux2_1 _24393_ (.A0(_02933_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .S(net262),
    .X(_01867_));
 sg13g2_mux2_1 _24394_ (.A0(_02934_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .S(net262),
    .X(_01868_));
 sg13g2_mux2_1 _24395_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net262),
    .X(_01869_));
 sg13g2_mux2_1 _24396_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(_06206_),
    .X(_01870_));
 sg13g2_nand2_1 _24397_ (.Y(_06210_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24398_ (.B1(_06210_),
    .Y(_01871_),
    .A1(net714),
    .A2(net262));
 sg13g2_mux2_1 _24399_ (.A0(net470),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(_06206_),
    .X(_01872_));
 sg13g2_nand2_1 _24400_ (.Y(_06211_),
    .A(_05982_),
    .B(net392));
 sg13g2_buf_2 _24401_ (.A(_06211_),
    .X(_06212_));
 sg13g2_buf_1 _24402_ (.A(_06212_),
    .X(_06213_));
 sg13g2_nand2_1 _24403_ (.Y(_06214_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(_06212_));
 sg13g2_o21ai_1 _24404_ (.B1(_06214_),
    .Y(_01873_),
    .A1(net637),
    .A2(_06213_));
 sg13g2_mux2_1 _24405_ (.A0(_03391_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net261),
    .X(_01874_));
 sg13g2_mux2_1 _24406_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S(_06213_),
    .X(_01875_));
 sg13g2_nand2_1 _24407_ (.Y(_06215_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(_06212_));
 sg13g2_o21ai_1 _24408_ (.B1(_06215_),
    .Y(_01876_),
    .A1(net698),
    .A2(net261));
 sg13g2_mux2_1 _24409_ (.A0(net725),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S(net261),
    .X(_01877_));
 sg13g2_mux2_1 _24410_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S(net261),
    .X(_01878_));
 sg13g2_mux2_1 _24411_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S(net261),
    .X(_01879_));
 sg13g2_mux2_1 _24412_ (.A0(_02934_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S(net261),
    .X(_01880_));
 sg13g2_mux2_1 _24413_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net261),
    .X(_01881_));
 sg13g2_mux2_1 _24414_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(_06212_),
    .X(_01882_));
 sg13g2_nand2_1 _24415_ (.Y(_06216_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .B(_06212_));
 sg13g2_o21ai_1 _24416_ (.B1(_06216_),
    .Y(_01883_),
    .A1(net714),
    .A2(net261));
 sg13g2_mux2_1 _24417_ (.A0(net470),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06212_),
    .X(_01884_));
 sg13g2_nand3_1 _24418_ (.B(_06062_),
    .C(_06008_),
    .A(_05843_),
    .Y(_06217_));
 sg13g2_buf_2 _24419_ (.A(_06217_),
    .X(_06218_));
 sg13g2_buf_1 _24420_ (.A(_06218_),
    .X(_06219_));
 sg13g2_nand2_1 _24421_ (.Y(_06220_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(_06218_));
 sg13g2_o21ai_1 _24422_ (.B1(_06220_),
    .Y(_01885_),
    .A1(net637),
    .A2(net328));
 sg13g2_mux2_1 _24423_ (.A0(net527),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(_06219_),
    .X(_01886_));
 sg13g2_mux2_1 _24424_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .S(_06219_),
    .X(_01887_));
 sg13g2_nand2_1 _24425_ (.Y(_06221_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(_06218_));
 sg13g2_o21ai_1 _24426_ (.B1(_06221_),
    .Y(_01888_),
    .A1(net698),
    .A2(net328));
 sg13g2_mux2_1 _24427_ (.A0(_02930_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .S(net328),
    .X(_01889_));
 sg13g2_mux2_1 _24428_ (.A0(net724),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .S(net328),
    .X(_01890_));
 sg13g2_mux2_1 _24429_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .S(net328),
    .X(_01891_));
 sg13g2_mux2_1 _24430_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .S(net328),
    .X(_01892_));
 sg13g2_mux2_1 _24431_ (.A0(_02935_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net328),
    .X(_01893_));
 sg13g2_mux2_1 _24432_ (.A0(_02936_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(_06218_),
    .X(_01894_));
 sg13g2_nand2_1 _24433_ (.Y(_06222_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .B(_06218_));
 sg13g2_o21ai_1 _24434_ (.B1(_06222_),
    .Y(_01895_),
    .A1(net714),
    .A2(net328));
 sg13g2_mux2_1 _24435_ (.A0(_03389_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(_06218_),
    .X(_01896_));
 sg13g2_nand2_1 _24436_ (.Y(_06223_),
    .A(_05843_),
    .B(_06069_));
 sg13g2_buf_2 _24437_ (.A(_06223_),
    .X(_06224_));
 sg13g2_buf_1 _24438_ (.A(_06224_),
    .X(_06225_));
 sg13g2_nand2_1 _24439_ (.Y(_06226_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(_06224_));
 sg13g2_o21ai_1 _24440_ (.B1(_06226_),
    .Y(_01897_),
    .A1(_03703_),
    .A2(net260));
 sg13g2_mux2_1 _24441_ (.A0(net527),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(_06225_),
    .X(_01898_));
 sg13g2_mux2_1 _24442_ (.A0(net642),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .S(_06225_),
    .X(_01899_));
 sg13g2_nand2_1 _24443_ (.Y(_06227_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(_06224_));
 sg13g2_o21ai_1 _24444_ (.B1(_06227_),
    .Y(_01900_),
    .A1(net698),
    .A2(net260));
 sg13g2_mux2_1 _24445_ (.A0(_02930_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .S(net260),
    .X(_01901_));
 sg13g2_mux2_1 _24446_ (.A0(_02932_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .S(net260),
    .X(_01902_));
 sg13g2_mux2_1 _24447_ (.A0(net723),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .S(net260),
    .X(_01903_));
 sg13g2_mux2_1 _24448_ (.A0(net847),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .S(net260),
    .X(_01904_));
 sg13g2_mux2_1 _24449_ (.A0(_02935_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net260),
    .X(_01905_));
 sg13g2_mux2_1 _24450_ (.A0(net845),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(_06224_),
    .X(_01906_));
 sg13g2_nand2_1 _24451_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .B(_06224_));
 sg13g2_o21ai_1 _24452_ (.B1(_06228_),
    .Y(_01907_),
    .A1(_03692_),
    .A2(net260));
 sg13g2_mux2_1 _24453_ (.A0(_03389_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(_06224_),
    .X(_01908_));
 sg13g2_mux2_1 _24454_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(_03395_),
    .S(_05824_),
    .X(_01909_));
 sg13g2_mux2_1 _24455_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(_03395_),
    .S(_05831_),
    .X(_01910_));
 sg13g2_buf_1 _24456_ (.A(net551),
    .X(_06229_));
 sg13g2_mux2_1 _24457_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net455),
    .S(_05840_),
    .X(_01911_));
 sg13g2_mux2_1 _24458_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net455),
    .S(_05847_),
    .X(_01912_));
 sg13g2_mux2_1 _24459_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net455),
    .S(_05852_),
    .X(_01913_));
 sg13g2_mux2_1 _24460_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(_06229_),
    .S(_05858_),
    .X(_01914_));
 sg13g2_mux2_1 _24461_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(_06229_),
    .S(_05862_),
    .X(_01915_));
 sg13g2_mux2_1 _24462_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net455),
    .S(_05872_),
    .X(_01916_));
 sg13g2_nand2_1 _24463_ (.Y(_06230_),
    .A(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .B(_05881_));
 sg13g2_o21ai_1 _24464_ (.B1(_06230_),
    .Y(_01917_),
    .A1(net638),
    .A2(net197));
 sg13g2_mux2_1 _24465_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net455),
    .S(_05890_),
    .X(_01918_));
 sg13g2_mux2_1 _24466_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net455),
    .S(_05896_),
    .X(_01919_));
 sg13g2_mux2_1 _24467_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(net455),
    .S(_05899_),
    .X(_01920_));
 sg13g2_mux2_1 _24468_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net455),
    .S(_05904_),
    .X(_01921_));
 sg13g2_buf_1 _24469_ (.A(_09119_),
    .X(_06231_));
 sg13g2_mux2_1 _24470_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net454),
    .S(_05909_),
    .X(_01922_));
 sg13g2_mux2_1 _24471_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(net454),
    .S(_05912_),
    .X(_01923_));
 sg13g2_mux2_1 _24472_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net454),
    .S(_05915_),
    .X(_01924_));
 sg13g2_mux2_1 _24473_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net454),
    .S(_05921_),
    .X(_01925_));
 sg13g2_nand2_1 _24474_ (.Y(_06232_),
    .A(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .B(_05925_));
 sg13g2_o21ai_1 _24475_ (.B1(_06232_),
    .Y(_01926_),
    .A1(_03699_),
    .A2(net196));
 sg13g2_mux2_1 _24476_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(_06231_),
    .S(_05932_),
    .X(_01927_));
 sg13g2_mux2_1 _24477_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(_06231_),
    .S(_05940_),
    .X(_01928_));
 sg13g2_mux2_1 _24478_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net454),
    .S(_05949_),
    .X(_01929_));
 sg13g2_mux2_1 _24479_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net454),
    .S(_05952_),
    .X(_01930_));
 sg13g2_mux2_1 _24480_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(net454),
    .S(_05955_),
    .X(_01931_));
 sg13g2_mux2_1 _24481_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net454),
    .S(_05958_),
    .X(_01932_));
 sg13g2_mux2_1 _24482_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net469),
    .S(_05961_),
    .X(_01933_));
 sg13g2_mux2_1 _24483_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net469),
    .S(_05964_),
    .X(_01934_));
 sg13g2_mux2_1 _24484_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net469),
    .S(_05968_),
    .X(_01935_));
 sg13g2_mux2_1 _24485_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net469),
    .S(_05973_),
    .X(_01936_));
 sg13g2_mux2_1 _24486_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net469),
    .S(_05979_),
    .X(_01937_));
 sg13g2_mux2_1 _24487_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(_03394_),
    .S(_05984_),
    .X(_01938_));
 sg13g2_mux2_1 _24488_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(_03394_),
    .S(_05988_),
    .X(_01939_));
 sg13g2_nand2_1 _24489_ (.Y(_06233_),
    .A(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .B(_05991_));
 sg13g2_o21ai_1 _24490_ (.B1(_06233_),
    .Y(_01940_),
    .A1(_03699_),
    .A2(net195));
 sg13g2_nor2_2 _24491_ (.A(net953),
    .B(_09109_),
    .Y(_06234_));
 sg13g2_nand3_1 _24492_ (.B(_00235_),
    .C(_06234_),
    .A(net1037),
    .Y(_06235_));
 sg13g2_buf_2 _24493_ (.A(_06235_),
    .X(_06236_));
 sg13g2_nor2_1 _24494_ (.A(net896),
    .B(_06236_),
    .Y(_06237_));
 sg13g2_buf_2 _24495_ (.A(_06237_),
    .X(_06238_));
 sg13g2_nand3_1 _24496_ (.B(_09963_),
    .C(_06238_),
    .A(net837),
    .Y(_06239_));
 sg13g2_buf_1 _24497_ (.A(_06239_),
    .X(_06240_));
 sg13g2_mux2_1 _24498_ (.A0(net989),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .S(_06240_),
    .X(_01957_));
 sg13g2_mux2_1 _24499_ (.A0(net988),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .S(_06240_),
    .X(_01958_));
 sg13g2_mux2_1 _24500_ (.A0(net987),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .S(_06240_),
    .X(_01959_));
 sg13g2_mux2_1 _24501_ (.A0(net1013),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .S(_06240_),
    .X(_01960_));
 sg13g2_nand3_1 _24502_ (.B(_04860_),
    .C(_06238_),
    .A(net837),
    .Y(_06241_));
 sg13g2_buf_2 _24503_ (.A(_06241_),
    .X(_06242_));
 sg13g2_mux2_1 _24504_ (.A0(net990),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .S(_06242_),
    .X(_01961_));
 sg13g2_mux2_1 _24505_ (.A0(net989),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06242_),
    .X(_01962_));
 sg13g2_mux2_1 _24506_ (.A0(net988),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06242_),
    .X(_01963_));
 sg13g2_mux2_1 _24507_ (.A0(net987),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .S(_06242_),
    .X(_01964_));
 sg13g2_mux2_1 _24508_ (.A0(net1013),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .S(_06242_),
    .X(_01965_));
 sg13g2_nand2b_1 _24509_ (.Y(_06243_),
    .B(_06238_),
    .A_N(_05327_));
 sg13g2_buf_4 _24510_ (.X(_06244_),
    .A(_06243_));
 sg13g2_mux2_1 _24511_ (.A0(net884),
    .A1(_04933_),
    .S(_06244_),
    .X(_01966_));
 sg13g2_buf_1 _24512_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06245_));
 sg13g2_mux2_1 _24513_ (.A0(net883),
    .A1(_06245_),
    .S(_06244_),
    .X(_01967_));
 sg13g2_mux2_1 _24514_ (.A0(net862),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(_06244_),
    .X(_01968_));
 sg13g2_buf_1 _24515_ (.A(\cpu.gpio.r_spi_miso_src[0][3] ),
    .X(_06246_));
 sg13g2_mux2_1 _24516_ (.A0(net990),
    .A1(_06246_),
    .S(_06244_),
    .X(_01969_));
 sg13g2_mux2_1 _24517_ (.A0(_11866_),
    .A1(_05503_),
    .S(_06244_),
    .X(_01970_));
 sg13g2_mux2_1 _24518_ (.A0(net988),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .S(_06244_),
    .X(_01971_));
 sg13g2_mux2_1 _24519_ (.A0(net987),
    .A1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .S(_06244_),
    .X(_01972_));
 sg13g2_buf_1 _24520_ (.A(\cpu.gpio.r_spi_miso_src[1][3] ),
    .X(_06247_));
 sg13g2_mux2_1 _24521_ (.A0(net1013),
    .A1(_06247_),
    .S(_06244_),
    .X(_01973_));
 sg13g2_nand2_1 _24522_ (.Y(_06248_),
    .A(net398),
    .B(_06238_));
 sg13g2_buf_4 _24523_ (.X(_06249_),
    .A(_06248_));
 sg13g2_mux2_1 _24524_ (.A0(net884),
    .A1(_04919_),
    .S(_06249_),
    .X(_01974_));
 sg13g2_mux2_1 _24525_ (.A0(net883),
    .A1(_05323_),
    .S(_06249_),
    .X(_01975_));
 sg13g2_mux2_1 _24526_ (.A0(net862),
    .A1(_05389_),
    .S(_06249_),
    .X(_01976_));
 sg13g2_mux2_1 _24527_ (.A0(net990),
    .A1(_05425_),
    .S(_06249_),
    .X(_01977_));
 sg13g2_mux2_1 _24528_ (.A0(net989),
    .A1(_05509_),
    .S(_06249_),
    .X(_01978_));
 sg13g2_mux2_1 _24529_ (.A0(net988),
    .A1(_05572_),
    .S(_06249_),
    .X(_01979_));
 sg13g2_mux2_1 _24530_ (.A0(net987),
    .A1(_05661_),
    .S(_06249_),
    .X(_01980_));
 sg13g2_mux2_1 _24531_ (.A0(net1013),
    .A1(_05003_),
    .S(_06249_),
    .X(_01981_));
 sg13g2_nand2_1 _24532_ (.Y(_06250_),
    .A(net397),
    .B(_06238_));
 sg13g2_buf_4 _24533_ (.X(_06251_),
    .A(_06250_));
 sg13g2_mux2_1 _24534_ (.A0(_09897_),
    .A1(_04925_),
    .S(_06251_),
    .X(_01982_));
 sg13g2_buf_1 _24535_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06252_));
 sg13g2_mux2_1 _24536_ (.A0(_09951_),
    .A1(_06252_),
    .S(_06251_),
    .X(_01983_));
 sg13g2_mux2_1 _24537_ (.A0(_11856_),
    .A1(\cpu.gpio.r_src_io[6][2] ),
    .S(_06251_),
    .X(_01984_));
 sg13g2_mux2_1 _24538_ (.A0(_11858_),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .S(_06251_),
    .X(_01985_));
 sg13g2_mux2_1 _24539_ (.A0(net989),
    .A1(_05496_),
    .S(_06251_),
    .X(_01986_));
 sg13g2_buf_1 _24540_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06253_));
 sg13g2_mux2_1 _24541_ (.A0(net988),
    .A1(_06253_),
    .S(_06251_),
    .X(_01987_));
 sg13g2_mux2_1 _24542_ (.A0(net987),
    .A1(\cpu.gpio.r_src_io[7][2] ),
    .S(_06251_),
    .X(_01988_));
 sg13g2_mux2_1 _24543_ (.A0(net1013),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .S(_06251_),
    .X(_01989_));
 sg13g2_nor4_2 _24544_ (.A(net865),
    .B(net896),
    .C(_05489_),
    .Y(_06254_),
    .D(_06236_));
 sg13g2_mux2_1 _24545_ (.A0(_05493_),
    .A1(net989),
    .S(_06254_),
    .X(_01990_));
 sg13g2_buf_1 _24546_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06255_));
 sg13g2_mux2_1 _24547_ (.A0(_06255_),
    .A1(net988),
    .S(_06254_),
    .X(_01991_));
 sg13g2_mux2_1 _24548_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(net987),
    .S(_06254_),
    .X(_01992_));
 sg13g2_mux2_1 _24549_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(_12006_),
    .S(_06254_),
    .X(_01993_));
 sg13g2_nand2_1 _24550_ (.Y(_06256_),
    .A(_04942_),
    .B(_06238_));
 sg13g2_buf_4 _24551_ (.X(_06257_),
    .A(_06256_));
 sg13g2_mux2_1 _24552_ (.A0(_09897_),
    .A1(_04943_),
    .S(_06257_),
    .X(_01994_));
 sg13g2_buf_1 _24553_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06258_));
 sg13g2_mux2_1 _24554_ (.A0(_09951_),
    .A1(_06258_),
    .S(_06257_),
    .X(_01995_));
 sg13g2_mux2_1 _24555_ (.A0(_11856_),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(_06257_),
    .X(_01996_));
 sg13g2_mux2_1 _24556_ (.A0(_11858_),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .S(_06257_),
    .X(_01997_));
 sg13g2_mux2_1 _24557_ (.A0(net989),
    .A1(_05511_),
    .S(_06257_),
    .X(_01998_));
 sg13g2_buf_1 _24558_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06259_));
 sg13g2_mux2_1 _24559_ (.A0(net988),
    .A1(_06259_),
    .S(_06257_),
    .X(_01999_));
 sg13g2_mux2_1 _24560_ (.A0(net987),
    .A1(\cpu.gpio.r_src_o[5][2] ),
    .S(_06257_),
    .X(_02000_));
 sg13g2_mux2_1 _24561_ (.A0(net1013),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .S(_06257_),
    .X(_02001_));
 sg13g2_nand2_2 _24562_ (.Y(_06260_),
    .A(_04940_),
    .B(_06238_));
 sg13g2_mux2_1 _24563_ (.A0(net989),
    .A1(_05498_),
    .S(_06260_),
    .X(_02006_));
 sg13g2_buf_1 _24564_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06261_));
 sg13g2_mux2_1 _24565_ (.A0(net988),
    .A1(_06261_),
    .S(_06260_),
    .X(_02007_));
 sg13g2_mux2_1 _24566_ (.A0(net987),
    .A1(\cpu.gpio.r_src_o[7][2] ),
    .S(_06260_),
    .X(_02008_));
 sg13g2_mux2_1 _24567_ (.A0(net1013),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .S(_06260_),
    .X(_02009_));
 sg13g2_buf_1 _24568_ (.A(net958),
    .X(_06262_));
 sg13g2_and2_1 _24569_ (.A(net691),
    .B(_08229_),
    .X(_06263_));
 sg13g2_buf_4 _24570_ (.X(_06264_),
    .A(_06263_));
 sg13g2_buf_1 _24571_ (.A(\cpu.icache.r_offset[2] ),
    .X(_06265_));
 sg13g2_buf_2 _24572_ (.A(_00253_),
    .X(_06266_));
 sg13g2_buf_1 _24573_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06267_));
 sg13g2_buf_1 _24574_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06268_));
 sg13g2_nand2b_1 _24575_ (.Y(_06269_),
    .B(_06268_),
    .A_N(_06267_));
 sg13g2_nor3_1 _24576_ (.A(_06265_),
    .B(_06266_),
    .C(_06269_),
    .Y(_06270_));
 sg13g2_buf_2 _24577_ (.A(_06270_),
    .X(_06271_));
 sg13g2_nand2_2 _24578_ (.Y(_06272_),
    .A(_06264_),
    .B(_06271_));
 sg13g2_mux2_1 _24579_ (.A0(net821),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06272_),
    .X(_02013_));
 sg13g2_buf_1 _24580_ (.A(net957),
    .X(_06273_));
 sg13g2_buf_1 _24581_ (.A(_00254_),
    .X(_06274_));
 sg13g2_inv_1 _24582_ (.Y(_06275_),
    .A(_06274_));
 sg13g2_nand2_1 _24583_ (.Y(_06276_),
    .A(_06267_),
    .B(_06268_));
 sg13g2_nor3_1 _24584_ (.A(_06266_),
    .B(_06275_),
    .C(_06276_),
    .Y(_06277_));
 sg13g2_buf_2 _24585_ (.A(_06277_),
    .X(_06278_));
 sg13g2_nand2_2 _24586_ (.Y(_06279_),
    .A(_06264_),
    .B(_06278_));
 sg13g2_mux2_1 _24587_ (.A0(_06273_),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06279_),
    .X(_02014_));
 sg13g2_buf_1 _24588_ (.A(net956),
    .X(_06280_));
 sg13g2_mux2_1 _24589_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06279_),
    .X(_02015_));
 sg13g2_nand2b_1 _24590_ (.Y(_06281_),
    .B(_06267_),
    .A_N(_06268_));
 sg13g2_nor3_1 _24591_ (.A(_06265_),
    .B(_06266_),
    .C(_06281_),
    .Y(_06282_));
 sg13g2_buf_2 _24592_ (.A(_06282_),
    .X(_06283_));
 sg13g2_nand2_2 _24593_ (.Y(_06284_),
    .A(_06264_),
    .B(_06283_));
 sg13g2_mux2_1 _24594_ (.A0(net821),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06284_),
    .X(_02016_));
 sg13g2_buf_1 _24595_ (.A(net955),
    .X(_06285_));
 sg13g2_mux2_1 _24596_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06284_),
    .X(_02017_));
 sg13g2_mux2_1 _24597_ (.A0(net820),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06284_),
    .X(_02018_));
 sg13g2_mux2_1 _24598_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06284_),
    .X(_02019_));
 sg13g2_nor3_1 _24599_ (.A(_06266_),
    .B(_06274_),
    .C(_06269_),
    .Y(_06286_));
 sg13g2_buf_2 _24600_ (.A(_06286_),
    .X(_06287_));
 sg13g2_nand2_2 _24601_ (.Y(_06288_),
    .A(_06264_),
    .B(_06287_));
 sg13g2_mux2_1 _24602_ (.A0(net821),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06288_),
    .X(_02020_));
 sg13g2_mux2_1 _24603_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06288_),
    .X(_02021_));
 sg13g2_mux2_1 _24604_ (.A0(net820),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06288_),
    .X(_02022_));
 sg13g2_mux2_1 _24605_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06288_),
    .X(_02023_));
 sg13g2_mux2_1 _24606_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06272_),
    .X(_02024_));
 sg13g2_nor4_1 _24607_ (.A(_06267_),
    .B(_06268_),
    .C(_06266_),
    .D(_06274_),
    .Y(_06289_));
 sg13g2_buf_2 _24608_ (.A(_06289_),
    .X(_06290_));
 sg13g2_nand2_2 _24609_ (.Y(_06291_),
    .A(_06264_),
    .B(_06290_));
 sg13g2_mux2_1 _24610_ (.A0(net821),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06291_),
    .X(_02025_));
 sg13g2_mux2_1 _24611_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06291_),
    .X(_02026_));
 sg13g2_mux2_1 _24612_ (.A0(net820),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06291_),
    .X(_02027_));
 sg13g2_mux2_1 _24613_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06291_),
    .X(_02028_));
 sg13g2_inv_1 _24614_ (.Y(_06292_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_1 _24615_ (.A(_06274_),
    .B(_06292_),
    .C(_06276_),
    .Y(_06293_));
 sg13g2_buf_2 _24616_ (.A(_06293_),
    .X(_06294_));
 sg13g2_nand2_1 _24617_ (.Y(_06295_),
    .A(_06264_),
    .B(_06294_));
 sg13g2_buf_1 _24618_ (.A(_06295_),
    .X(_06296_));
 sg13g2_buf_1 _24619_ (.A(_06296_),
    .X(_06297_));
 sg13g2_mux2_1 _24620_ (.A0(_06262_),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(_06297_),
    .X(_02029_));
 sg13g2_mux2_1 _24621_ (.A0(_06285_),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(_06297_),
    .X(_02030_));
 sg13g2_buf_1 _24622_ (.A(_06296_),
    .X(_06298_));
 sg13g2_mux2_1 _24623_ (.A0(_06273_),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(_06298_),
    .X(_02031_));
 sg13g2_mux2_1 _24624_ (.A0(_06280_),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(_06298_),
    .X(_02032_));
 sg13g2_nor3_1 _24625_ (.A(_06266_),
    .B(_06274_),
    .C(_06281_),
    .Y(_06299_));
 sg13g2_buf_2 _24626_ (.A(_06299_),
    .X(_06300_));
 sg13g2_nand2_2 _24627_ (.Y(_06301_),
    .A(_06264_),
    .B(_06300_));
 sg13g2_mux2_1 _24628_ (.A0(net821),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06301_),
    .X(_02033_));
 sg13g2_mux2_1 _24629_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06301_),
    .X(_02034_));
 sg13g2_mux2_1 _24630_ (.A0(net820),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06272_),
    .X(_02035_));
 sg13g2_mux2_1 _24631_ (.A0(net820),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06301_),
    .X(_02036_));
 sg13g2_mux2_1 _24632_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06301_),
    .X(_02037_));
 sg13g2_mux2_1 _24633_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06272_),
    .X(_02038_));
 sg13g2_nor4_1 _24634_ (.A(_06267_),
    .B(_06268_),
    .C(_06265_),
    .D(_06266_),
    .Y(_06302_));
 sg13g2_buf_2 _24635_ (.A(_06302_),
    .X(_06303_));
 sg13g2_nand2_2 _24636_ (.Y(_06304_),
    .A(_06264_),
    .B(_06303_));
 sg13g2_mux2_1 _24637_ (.A0(net821),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06304_),
    .X(_02039_));
 sg13g2_mux2_1 _24638_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06304_),
    .X(_02040_));
 sg13g2_mux2_1 _24639_ (.A0(net820),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06304_),
    .X(_02041_));
 sg13g2_mux2_1 _24640_ (.A0(net819),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06304_),
    .X(_02042_));
 sg13g2_mux2_1 _24641_ (.A0(_06262_),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06279_),
    .X(_02043_));
 sg13g2_mux2_1 _24642_ (.A0(net818),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06279_),
    .X(_02044_));
 sg13g2_buf_1 _24643_ (.A(net958),
    .X(_06305_));
 sg13g2_and2_1 _24644_ (.A(net441),
    .B(_06271_),
    .X(_06306_));
 sg13g2_buf_1 _24645_ (.A(_06306_),
    .X(_06307_));
 sg13g2_mux2_1 _24646_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net817),
    .S(_06307_),
    .X(_02045_));
 sg13g2_buf_1 _24647_ (.A(net957),
    .X(_06308_));
 sg13g2_and2_1 _24648_ (.A(_08909_),
    .B(_06278_),
    .X(_06309_));
 sg13g2_buf_1 _24649_ (.A(_06309_),
    .X(_06310_));
 sg13g2_mux2_1 _24650_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net816),
    .S(_06310_),
    .X(_02046_));
 sg13g2_buf_1 _24651_ (.A(net956),
    .X(_06311_));
 sg13g2_mux2_1 _24652_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net815),
    .S(_06310_),
    .X(_02047_));
 sg13g2_and2_1 _24653_ (.A(net441),
    .B(_06283_),
    .X(_06312_));
 sg13g2_buf_1 _24654_ (.A(_06312_),
    .X(_06313_));
 sg13g2_mux2_1 _24655_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net817),
    .S(_06313_),
    .X(_02048_));
 sg13g2_buf_1 _24656_ (.A(net955),
    .X(_06314_));
 sg13g2_mux2_1 _24657_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net814),
    .S(_06313_),
    .X(_02049_));
 sg13g2_mux2_1 _24658_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net816),
    .S(_06313_),
    .X(_02050_));
 sg13g2_mux2_1 _24659_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net815),
    .S(_06313_),
    .X(_02051_));
 sg13g2_and2_1 _24660_ (.A(net441),
    .B(_06287_),
    .X(_06315_));
 sg13g2_buf_1 _24661_ (.A(_06315_),
    .X(_06316_));
 sg13g2_mux2_1 _24662_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net817),
    .S(_06316_),
    .X(_02052_));
 sg13g2_mux2_1 _24663_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net814),
    .S(_06316_),
    .X(_02053_));
 sg13g2_mux2_1 _24664_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net816),
    .S(_06316_),
    .X(_02054_));
 sg13g2_mux2_1 _24665_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net815),
    .S(_06316_),
    .X(_02055_));
 sg13g2_mux2_1 _24666_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net814),
    .S(_06307_),
    .X(_02056_));
 sg13g2_buf_1 _24667_ (.A(net958),
    .X(_06317_));
 sg13g2_and2_1 _24668_ (.A(net441),
    .B(_06290_),
    .X(_06318_));
 sg13g2_buf_2 _24669_ (.A(_06318_),
    .X(_06319_));
 sg13g2_mux2_1 _24670_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net813),
    .S(_06319_),
    .X(_02057_));
 sg13g2_buf_1 _24671_ (.A(net955),
    .X(_06320_));
 sg13g2_mux2_1 _24672_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net812),
    .S(_06319_),
    .X(_02058_));
 sg13g2_buf_1 _24673_ (.A(net957),
    .X(_06321_));
 sg13g2_mux2_1 _24674_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net811),
    .S(_06319_),
    .X(_02059_));
 sg13g2_buf_1 _24675_ (.A(net956),
    .X(_06322_));
 sg13g2_mux2_1 _24676_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net810),
    .S(_06319_),
    .X(_02060_));
 sg13g2_and2_1 _24677_ (.A(net441),
    .B(_06294_),
    .X(_06323_));
 sg13g2_buf_2 _24678_ (.A(_06323_),
    .X(_06324_));
 sg13g2_mux2_1 _24679_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net813),
    .S(_06324_),
    .X(_02061_));
 sg13g2_mux2_1 _24680_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net812),
    .S(_06324_),
    .X(_02062_));
 sg13g2_mux2_1 _24681_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(net811),
    .S(_06324_),
    .X(_02063_));
 sg13g2_mux2_1 _24682_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net810),
    .S(_06324_),
    .X(_02064_));
 sg13g2_and2_1 _24683_ (.A(net441),
    .B(_06300_),
    .X(_06325_));
 sg13g2_buf_1 _24684_ (.A(_06325_),
    .X(_06326_));
 sg13g2_mux2_1 _24685_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net813),
    .S(_06326_),
    .X(_02065_));
 sg13g2_mux2_1 _24686_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net812),
    .S(_06326_),
    .X(_02066_));
 sg13g2_mux2_1 _24687_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net811),
    .S(_06307_),
    .X(_02067_));
 sg13g2_mux2_1 _24688_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net811),
    .S(_06326_),
    .X(_02068_));
 sg13g2_mux2_1 _24689_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net810),
    .S(_06326_),
    .X(_02069_));
 sg13g2_mux2_1 _24690_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net810),
    .S(_06307_),
    .X(_02070_));
 sg13g2_and2_1 _24691_ (.A(net441),
    .B(_06303_),
    .X(_06327_));
 sg13g2_buf_1 _24692_ (.A(_06327_),
    .X(_06328_));
 sg13g2_mux2_1 _24693_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(_06317_),
    .S(_06328_),
    .X(_02071_));
 sg13g2_mux2_1 _24694_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net812),
    .S(_06328_),
    .X(_02072_));
 sg13g2_mux2_1 _24695_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(_06321_),
    .S(_06328_),
    .X(_02073_));
 sg13g2_mux2_1 _24696_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net810),
    .S(_06328_),
    .X(_02074_));
 sg13g2_mux2_1 _24697_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(net813),
    .S(_06310_),
    .X(_02075_));
 sg13g2_mux2_1 _24698_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(net812),
    .S(_06310_),
    .X(_02076_));
 sg13g2_and2_1 _24699_ (.A(net378),
    .B(_06271_),
    .X(_06329_));
 sg13g2_buf_1 _24700_ (.A(_06329_),
    .X(_06330_));
 sg13g2_mux2_1 _24701_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(_06317_),
    .S(_06330_),
    .X(_02077_));
 sg13g2_and2_1 _24702_ (.A(net378),
    .B(_06278_),
    .X(_06331_));
 sg13g2_buf_1 _24703_ (.A(_06331_),
    .X(_06332_));
 sg13g2_mux2_1 _24704_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(net811),
    .S(_06332_),
    .X(_02078_));
 sg13g2_mux2_1 _24705_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(_06322_),
    .S(_06332_),
    .X(_02079_));
 sg13g2_and2_1 _24706_ (.A(net378),
    .B(_06283_),
    .X(_06333_));
 sg13g2_buf_1 _24707_ (.A(_06333_),
    .X(_06334_));
 sg13g2_mux2_1 _24708_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net813),
    .S(_06334_),
    .X(_02080_));
 sg13g2_mux2_1 _24709_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(net812),
    .S(_06334_),
    .X(_02081_));
 sg13g2_mux2_1 _24710_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net811),
    .S(_06334_),
    .X(_02082_));
 sg13g2_mux2_1 _24711_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net810),
    .S(_06334_),
    .X(_02083_));
 sg13g2_and2_1 _24712_ (.A(net378),
    .B(_06287_),
    .X(_06335_));
 sg13g2_buf_2 _24713_ (.A(_06335_),
    .X(_06336_));
 sg13g2_mux2_1 _24714_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net813),
    .S(_06336_),
    .X(_02084_));
 sg13g2_mux2_1 _24715_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(net812),
    .S(_06336_),
    .X(_02085_));
 sg13g2_mux2_1 _24716_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net811),
    .S(_06336_),
    .X(_02086_));
 sg13g2_mux2_1 _24717_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net810),
    .S(_06336_),
    .X(_02087_));
 sg13g2_mux2_1 _24718_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(_06320_),
    .S(_06330_),
    .X(_02088_));
 sg13g2_and2_1 _24719_ (.A(net378),
    .B(_06290_),
    .X(_06337_));
 sg13g2_buf_2 _24720_ (.A(_06337_),
    .X(_06338_));
 sg13g2_mux2_1 _24721_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net813),
    .S(_06338_),
    .X(_02089_));
 sg13g2_mux2_1 _24722_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net812),
    .S(_06338_),
    .X(_02090_));
 sg13g2_mux2_1 _24723_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net811),
    .S(_06338_),
    .X(_02091_));
 sg13g2_mux2_1 _24724_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(_06322_),
    .S(_06338_),
    .X(_02092_));
 sg13g2_and2_1 _24725_ (.A(net378),
    .B(_06294_),
    .X(_06339_));
 sg13g2_buf_2 _24726_ (.A(_06339_),
    .X(_06340_));
 sg13g2_mux2_1 _24727_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net813),
    .S(_06340_),
    .X(_02093_));
 sg13g2_mux2_1 _24728_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(_06320_),
    .S(_06340_),
    .X(_02094_));
 sg13g2_mux2_1 _24729_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(_06321_),
    .S(_06340_),
    .X(_02095_));
 sg13g2_mux2_1 _24730_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net810),
    .S(_06340_),
    .X(_02096_));
 sg13g2_buf_1 _24731_ (.A(_11761_),
    .X(_06341_));
 sg13g2_and2_1 _24732_ (.A(net378),
    .B(_06300_),
    .X(_06342_));
 sg13g2_buf_1 _24733_ (.A(_06342_),
    .X(_06343_));
 sg13g2_mux2_1 _24734_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net931),
    .S(_06343_),
    .X(_02097_));
 sg13g2_buf_1 _24735_ (.A(_11832_),
    .X(_06344_));
 sg13g2_mux2_1 _24736_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net930),
    .S(_06343_),
    .X(_02098_));
 sg13g2_buf_1 _24737_ (.A(_11795_),
    .X(_06345_));
 sg13g2_mux2_1 _24738_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(_06345_),
    .S(_06330_),
    .X(_02099_));
 sg13g2_mux2_1 _24739_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net929),
    .S(_06343_),
    .X(_02100_));
 sg13g2_buf_1 _24740_ (.A(_11812_),
    .X(_06346_));
 sg13g2_mux2_1 _24741_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net928),
    .S(_06343_),
    .X(_02101_));
 sg13g2_mux2_1 _24742_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net928),
    .S(_06330_),
    .X(_02102_));
 sg13g2_and2_1 _24743_ (.A(_08908_),
    .B(_06303_),
    .X(_06347_));
 sg13g2_buf_1 _24744_ (.A(_06347_),
    .X(_06348_));
 sg13g2_mux2_1 _24745_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(_06341_),
    .S(_06348_),
    .X(_02103_));
 sg13g2_mux2_1 _24746_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(_06344_),
    .S(_06348_),
    .X(_02104_));
 sg13g2_mux2_1 _24747_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(_06345_),
    .S(_06348_),
    .X(_02105_));
 sg13g2_mux2_1 _24748_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(_06346_),
    .S(_06348_),
    .X(_02106_));
 sg13g2_mux2_1 _24749_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net931),
    .S(_06332_),
    .X(_02107_));
 sg13g2_mux2_1 _24750_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net930),
    .S(_06332_),
    .X(_02108_));
 sg13g2_nand2_2 _24751_ (.Y(_06349_),
    .A(net386),
    .B(_06271_));
 sg13g2_mux2_1 _24752_ (.A0(net821),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06349_),
    .X(_02109_));
 sg13g2_and2_1 _24753_ (.A(_08341_),
    .B(_06278_),
    .X(_06350_));
 sg13g2_buf_1 _24754_ (.A(_06350_),
    .X(_06351_));
 sg13g2_mux2_1 _24755_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net929),
    .S(_06351_),
    .X(_02110_));
 sg13g2_mux2_1 _24756_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net928),
    .S(_06351_),
    .X(_02111_));
 sg13g2_nand2_2 _24757_ (.Y(_06352_),
    .A(net386),
    .B(_06283_));
 sg13g2_mux2_1 _24758_ (.A0(net821),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06352_),
    .X(_02112_));
 sg13g2_mux2_1 _24759_ (.A0(net818),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06352_),
    .X(_02113_));
 sg13g2_mux2_1 _24760_ (.A0(net820),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06352_),
    .X(_02114_));
 sg13g2_mux2_1 _24761_ (.A0(_06280_),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06352_),
    .X(_02115_));
 sg13g2_buf_1 _24762_ (.A(_02788_),
    .X(_06353_));
 sg13g2_nand2_2 _24763_ (.Y(_06354_),
    .A(net386),
    .B(_06287_));
 sg13g2_mux2_1 _24764_ (.A0(net809),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06354_),
    .X(_02116_));
 sg13g2_mux2_1 _24765_ (.A0(_06285_),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06354_),
    .X(_02117_));
 sg13g2_mux2_1 _24766_ (.A0(net820),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06354_),
    .X(_02118_));
 sg13g2_mux2_1 _24767_ (.A0(net819),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06354_),
    .X(_02119_));
 sg13g2_buf_1 _24768_ (.A(_02805_),
    .X(_06355_));
 sg13g2_mux2_1 _24769_ (.A0(net808),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06349_),
    .X(_02120_));
 sg13g2_nand2_2 _24770_ (.Y(_06356_),
    .A(net386),
    .B(_06290_));
 sg13g2_mux2_1 _24771_ (.A0(net809),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06356_),
    .X(_02121_));
 sg13g2_mux2_1 _24772_ (.A0(net808),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06356_),
    .X(_02122_));
 sg13g2_buf_1 _24773_ (.A(_02797_),
    .X(_06357_));
 sg13g2_mux2_1 _24774_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06356_),
    .X(_02123_));
 sg13g2_buf_1 _24775_ (.A(_02801_),
    .X(_06358_));
 sg13g2_mux2_1 _24776_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06356_),
    .X(_02124_));
 sg13g2_nand2_1 _24777_ (.Y(_06359_),
    .A(_08341_),
    .B(_06294_));
 sg13g2_buf_1 _24778_ (.A(_06359_),
    .X(_06360_));
 sg13g2_buf_1 _24779_ (.A(_06360_),
    .X(_06361_));
 sg13g2_mux2_1 _24780_ (.A0(_06353_),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(_06361_),
    .X(_02125_));
 sg13g2_mux2_1 _24781_ (.A0(net808),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net221),
    .X(_02126_));
 sg13g2_buf_1 _24782_ (.A(_06360_),
    .X(_06362_));
 sg13g2_mux2_1 _24783_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net220),
    .X(_02127_));
 sg13g2_mux2_1 _24784_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net220),
    .X(_02128_));
 sg13g2_nand2_2 _24785_ (.Y(_06363_),
    .A(net386),
    .B(_06300_));
 sg13g2_mux2_1 _24786_ (.A0(net809),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06363_),
    .X(_02129_));
 sg13g2_mux2_1 _24787_ (.A0(net808),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06363_),
    .X(_02130_));
 sg13g2_mux2_1 _24788_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06349_),
    .X(_02131_));
 sg13g2_mux2_1 _24789_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06363_),
    .X(_02132_));
 sg13g2_mux2_1 _24790_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06363_),
    .X(_02133_));
 sg13g2_mux2_1 _24791_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06349_),
    .X(_02134_));
 sg13g2_nand2_2 _24792_ (.Y(_06364_),
    .A(net386),
    .B(_06303_));
 sg13g2_mux2_1 _24793_ (.A0(_06353_),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06364_),
    .X(_02135_));
 sg13g2_mux2_1 _24794_ (.A0(_06355_),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06364_),
    .X(_02136_));
 sg13g2_mux2_1 _24795_ (.A0(net807),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06364_),
    .X(_02137_));
 sg13g2_mux2_1 _24796_ (.A0(net806),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06364_),
    .X(_02138_));
 sg13g2_mux2_1 _24797_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(net931),
    .S(_06351_),
    .X(_02139_));
 sg13g2_mux2_1 _24798_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net930),
    .S(_06351_),
    .X(_02140_));
 sg13g2_nand2_2 _24799_ (.Y(_06365_),
    .A(net554),
    .B(_06271_));
 sg13g2_mux2_1 _24800_ (.A0(net809),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06365_),
    .X(_02141_));
 sg13g2_and2_1 _24801_ (.A(net554),
    .B(_06278_),
    .X(_06366_));
 sg13g2_buf_1 _24802_ (.A(_06366_),
    .X(_06367_));
 sg13g2_mux2_1 _24803_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(net929),
    .S(_06367_),
    .X(_02142_));
 sg13g2_mux2_1 _24804_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net928),
    .S(_06367_),
    .X(_02143_));
 sg13g2_nand2_2 _24805_ (.Y(_06368_),
    .A(net554),
    .B(_06283_));
 sg13g2_mux2_1 _24806_ (.A0(net809),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06368_),
    .X(_02144_));
 sg13g2_mux2_1 _24807_ (.A0(net808),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06368_),
    .X(_02145_));
 sg13g2_mux2_1 _24808_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06368_),
    .X(_02146_));
 sg13g2_mux2_1 _24809_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06368_),
    .X(_02147_));
 sg13g2_nand2_2 _24810_ (.Y(_06369_),
    .A(net554),
    .B(_06287_));
 sg13g2_mux2_1 _24811_ (.A0(net809),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06369_),
    .X(_02148_));
 sg13g2_mux2_1 _24812_ (.A0(net808),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06369_),
    .X(_02149_));
 sg13g2_mux2_1 _24813_ (.A0(_06357_),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06369_),
    .X(_02150_));
 sg13g2_mux2_1 _24814_ (.A0(_06358_),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06369_),
    .X(_02151_));
 sg13g2_mux2_1 _24815_ (.A0(_06355_),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06365_),
    .X(_02152_));
 sg13g2_nand2_2 _24816_ (.Y(_06370_),
    .A(_08894_),
    .B(_06290_));
 sg13g2_mux2_1 _24817_ (.A0(net809),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06370_),
    .X(_02153_));
 sg13g2_mux2_1 _24818_ (.A0(net808),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06370_),
    .X(_02154_));
 sg13g2_mux2_1 _24819_ (.A0(_06357_),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06370_),
    .X(_02155_));
 sg13g2_mux2_1 _24820_ (.A0(_06358_),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06370_),
    .X(_02156_));
 sg13g2_and2_1 _24821_ (.A(_08894_),
    .B(_06294_),
    .X(_06371_));
 sg13g2_buf_2 _24822_ (.A(_06371_),
    .X(_06372_));
 sg13g2_mux2_1 _24823_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net931),
    .S(_06372_),
    .X(_02157_));
 sg13g2_mux2_1 _24824_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net930),
    .S(_06372_),
    .X(_02158_));
 sg13g2_mux2_1 _24825_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net929),
    .S(_06372_),
    .X(_02159_));
 sg13g2_mux2_1 _24826_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(net928),
    .S(_06372_),
    .X(_02160_));
 sg13g2_nand2_2 _24827_ (.Y(_06373_),
    .A(net554),
    .B(_06300_));
 sg13g2_mux2_1 _24828_ (.A0(net809),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06373_),
    .X(_02161_));
 sg13g2_mux2_1 _24829_ (.A0(net808),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06373_),
    .X(_02162_));
 sg13g2_mux2_1 _24830_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06365_),
    .X(_02163_));
 sg13g2_mux2_1 _24831_ (.A0(net807),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06373_),
    .X(_02164_));
 sg13g2_mux2_1 _24832_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06373_),
    .X(_02165_));
 sg13g2_mux2_1 _24833_ (.A0(net806),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06365_),
    .X(_02166_));
 sg13g2_buf_1 _24834_ (.A(_02788_),
    .X(_06374_));
 sg13g2_nand2_2 _24835_ (.Y(_06375_),
    .A(net554),
    .B(_06303_));
 sg13g2_mux2_1 _24836_ (.A0(_06374_),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06375_),
    .X(_02167_));
 sg13g2_buf_1 _24837_ (.A(_02805_),
    .X(_06376_));
 sg13g2_mux2_1 _24838_ (.A0(net804),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06375_),
    .X(_02168_));
 sg13g2_buf_1 _24839_ (.A(_02797_),
    .X(_06377_));
 sg13g2_mux2_1 _24840_ (.A0(net803),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06375_),
    .X(_02169_));
 sg13g2_buf_1 _24841_ (.A(_02801_),
    .X(_06378_));
 sg13g2_mux2_1 _24842_ (.A0(net802),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06375_),
    .X(_02170_));
 sg13g2_mux2_1 _24843_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(net931),
    .S(_06367_),
    .X(_02171_));
 sg13g2_mux2_1 _24844_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(_06344_),
    .S(_06367_),
    .X(_02172_));
 sg13g2_nand2_2 _24845_ (.Y(_06379_),
    .A(net446),
    .B(_06271_));
 sg13g2_mux2_1 _24846_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][0] ),
    .S(_06379_),
    .X(_02173_));
 sg13g2_nand2_2 _24847_ (.Y(_06380_),
    .A(net446),
    .B(_06278_));
 sg13g2_mux2_1 _24848_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][10] ),
    .S(_06380_),
    .X(_02174_));
 sg13g2_mux2_1 _24849_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][11] ),
    .S(_06380_),
    .X(_02175_));
 sg13g2_nand2_2 _24850_ (.Y(_06381_),
    .A(net446),
    .B(_06283_));
 sg13g2_mux2_1 _24851_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][12] ),
    .S(_06381_),
    .X(_02176_));
 sg13g2_mux2_1 _24852_ (.A0(net804),
    .A1(\cpu.icache.r_data[5][13] ),
    .S(_06381_),
    .X(_02177_));
 sg13g2_mux2_1 _24853_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][14] ),
    .S(_06381_),
    .X(_02178_));
 sg13g2_mux2_1 _24854_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][15] ),
    .S(_06381_),
    .X(_02179_));
 sg13g2_nand2_2 _24855_ (.Y(_06382_),
    .A(net446),
    .B(_06287_));
 sg13g2_mux2_1 _24856_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][16] ),
    .S(_06382_),
    .X(_02180_));
 sg13g2_mux2_1 _24857_ (.A0(net804),
    .A1(\cpu.icache.r_data[5][17] ),
    .S(_06382_),
    .X(_02181_));
 sg13g2_mux2_1 _24858_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][18] ),
    .S(_06382_),
    .X(_02182_));
 sg13g2_mux2_1 _24859_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][19] ),
    .S(_06382_),
    .X(_02183_));
 sg13g2_mux2_1 _24860_ (.A0(net804),
    .A1(\cpu.icache.r_data[5][1] ),
    .S(_06379_),
    .X(_02184_));
 sg13g2_nand2_2 _24861_ (.Y(_06383_),
    .A(_08346_),
    .B(_06290_));
 sg13g2_mux2_1 _24862_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][20] ),
    .S(_06383_),
    .X(_02185_));
 sg13g2_mux2_1 _24863_ (.A0(_06376_),
    .A1(\cpu.icache.r_data[5][21] ),
    .S(_06383_),
    .X(_02186_));
 sg13g2_mux2_1 _24864_ (.A0(_06377_),
    .A1(\cpu.icache.r_data[5][22] ),
    .S(_06383_),
    .X(_02187_));
 sg13g2_mux2_1 _24865_ (.A0(_06378_),
    .A1(\cpu.icache.r_data[5][23] ),
    .S(_06383_),
    .X(_02188_));
 sg13g2_nand2_1 _24866_ (.Y(_06384_),
    .A(_08346_),
    .B(_06294_));
 sg13g2_buf_2 _24867_ (.A(_06384_),
    .X(_06385_));
 sg13g2_mux2_1 _24868_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][24] ),
    .S(_06385_),
    .X(_02189_));
 sg13g2_mux2_1 _24869_ (.A0(net804),
    .A1(\cpu.icache.r_data[5][25] ),
    .S(_06385_),
    .X(_02190_));
 sg13g2_mux2_1 _24870_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][26] ),
    .S(_06385_),
    .X(_02191_));
 sg13g2_mux2_1 _24871_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][27] ),
    .S(_06385_),
    .X(_02192_));
 sg13g2_nand2_2 _24872_ (.Y(_06386_),
    .A(net446),
    .B(_06300_));
 sg13g2_mux2_1 _24873_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][28] ),
    .S(_06386_),
    .X(_02193_));
 sg13g2_mux2_1 _24874_ (.A0(net804),
    .A1(\cpu.icache.r_data[5][29] ),
    .S(_06386_),
    .X(_02194_));
 sg13g2_mux2_1 _24875_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][2] ),
    .S(_06379_),
    .X(_02195_));
 sg13g2_mux2_1 _24876_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][30] ),
    .S(_06386_),
    .X(_02196_));
 sg13g2_mux2_1 _24877_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][31] ),
    .S(_06386_),
    .X(_02197_));
 sg13g2_mux2_1 _24878_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][3] ),
    .S(_06379_),
    .X(_02198_));
 sg13g2_nand2_2 _24879_ (.Y(_06387_),
    .A(net446),
    .B(_06303_));
 sg13g2_mux2_1 _24880_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][4] ),
    .S(_06387_),
    .X(_02199_));
 sg13g2_mux2_1 _24881_ (.A0(net804),
    .A1(\cpu.icache.r_data[5][5] ),
    .S(_06387_),
    .X(_02200_));
 sg13g2_mux2_1 _24882_ (.A0(net803),
    .A1(\cpu.icache.r_data[5][6] ),
    .S(_06387_),
    .X(_02201_));
 sg13g2_mux2_1 _24883_ (.A0(net802),
    .A1(\cpu.icache.r_data[5][7] ),
    .S(_06387_),
    .X(_02202_));
 sg13g2_mux2_1 _24884_ (.A0(net805),
    .A1(\cpu.icache.r_data[5][8] ),
    .S(_06380_),
    .X(_02203_));
 sg13g2_mux2_1 _24885_ (.A0(_06376_),
    .A1(\cpu.icache.r_data[5][9] ),
    .S(_06380_),
    .X(_02204_));
 sg13g2_nand2_2 _24886_ (.Y(_06388_),
    .A(net553),
    .B(_06271_));
 sg13g2_mux2_1 _24887_ (.A0(_06374_),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_06388_),
    .X(_02205_));
 sg13g2_nand2_2 _24888_ (.Y(_06389_),
    .A(net553),
    .B(_06278_));
 sg13g2_mux2_1 _24889_ (.A0(_06377_),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(_06389_),
    .X(_02206_));
 sg13g2_mux2_1 _24890_ (.A0(_06378_),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(_06389_),
    .X(_02207_));
 sg13g2_nand2_2 _24891_ (.Y(_06390_),
    .A(net553),
    .B(_06283_));
 sg13g2_mux2_1 _24892_ (.A0(net817),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_06390_),
    .X(_02208_));
 sg13g2_mux2_1 _24893_ (.A0(net804),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(_06390_),
    .X(_02209_));
 sg13g2_mux2_1 _24894_ (.A0(net816),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(_06390_),
    .X(_02210_));
 sg13g2_mux2_1 _24895_ (.A0(net815),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(_06390_),
    .X(_02211_));
 sg13g2_nand2_2 _24896_ (.Y(_06391_),
    .A(net553),
    .B(_06287_));
 sg13g2_mux2_1 _24897_ (.A0(net817),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(_06391_),
    .X(_02212_));
 sg13g2_mux2_1 _24898_ (.A0(net814),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(_06391_),
    .X(_02213_));
 sg13g2_mux2_1 _24899_ (.A0(net816),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(_06391_),
    .X(_02214_));
 sg13g2_mux2_1 _24900_ (.A0(net815),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(_06391_),
    .X(_02215_));
 sg13g2_mux2_1 _24901_ (.A0(_06314_),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_06388_),
    .X(_02216_));
 sg13g2_nand2_2 _24902_ (.Y(_06392_),
    .A(net553),
    .B(_06290_));
 sg13g2_mux2_1 _24903_ (.A0(net817),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_06392_),
    .X(_02217_));
 sg13g2_mux2_1 _24904_ (.A0(net814),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_06392_),
    .X(_02218_));
 sg13g2_mux2_1 _24905_ (.A0(_06308_),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_06392_),
    .X(_02219_));
 sg13g2_mux2_1 _24906_ (.A0(_06311_),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_06392_),
    .X(_02220_));
 sg13g2_nand2_1 _24907_ (.Y(_06393_),
    .A(_08899_),
    .B(_06294_));
 sg13g2_buf_2 _24908_ (.A(_06393_),
    .X(_06394_));
 sg13g2_mux2_1 _24909_ (.A0(net817),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_06394_),
    .X(_02221_));
 sg13g2_mux2_1 _24910_ (.A0(net814),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_06394_),
    .X(_02222_));
 sg13g2_mux2_1 _24911_ (.A0(net816),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(_06394_),
    .X(_02223_));
 sg13g2_mux2_1 _24912_ (.A0(net815),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_06394_),
    .X(_02224_));
 sg13g2_nand2_2 _24913_ (.Y(_06395_),
    .A(net553),
    .B(_06300_));
 sg13g2_mux2_1 _24914_ (.A0(net817),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_06395_),
    .X(_02225_));
 sg13g2_mux2_1 _24915_ (.A0(net814),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(_06395_),
    .X(_02226_));
 sg13g2_mux2_1 _24916_ (.A0(net816),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_06388_),
    .X(_02227_));
 sg13g2_mux2_1 _24917_ (.A0(net816),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_06395_),
    .X(_02228_));
 sg13g2_mux2_1 _24918_ (.A0(net815),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(_06395_),
    .X(_02229_));
 sg13g2_mux2_1 _24919_ (.A0(net815),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(_06388_),
    .X(_02230_));
 sg13g2_nand2_2 _24920_ (.Y(_06396_),
    .A(_08899_),
    .B(_06303_));
 sg13g2_mux2_1 _24921_ (.A0(_06305_),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(_06396_),
    .X(_02231_));
 sg13g2_mux2_1 _24922_ (.A0(net814),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_06396_),
    .X(_02232_));
 sg13g2_mux2_1 _24923_ (.A0(_06308_),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(_06396_),
    .X(_02233_));
 sg13g2_mux2_1 _24924_ (.A0(_06311_),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(_06396_),
    .X(_02234_));
 sg13g2_mux2_1 _24925_ (.A0(_06305_),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_06389_),
    .X(_02235_));
 sg13g2_mux2_1 _24926_ (.A0(_06314_),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(_06389_),
    .X(_02236_));
 sg13g2_and2_1 _24927_ (.A(net440),
    .B(_06271_),
    .X(_06397_));
 sg13g2_buf_2 _24928_ (.A(_06397_),
    .X(_06398_));
 sg13g2_mux2_1 _24929_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(_06341_),
    .S(_06398_),
    .X(_02237_));
 sg13g2_and2_1 _24930_ (.A(net440),
    .B(_06278_),
    .X(_06399_));
 sg13g2_buf_1 _24931_ (.A(_06399_),
    .X(_06400_));
 sg13g2_mux2_1 _24932_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net929),
    .S(_06400_),
    .X(_02238_));
 sg13g2_mux2_1 _24933_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net928),
    .S(_06400_),
    .X(_02239_));
 sg13g2_and2_1 _24934_ (.A(net440),
    .B(_06283_),
    .X(_06401_));
 sg13g2_buf_1 _24935_ (.A(_06401_),
    .X(_06402_));
 sg13g2_mux2_1 _24936_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(net931),
    .S(_06402_),
    .X(_02240_));
 sg13g2_mux2_1 _24937_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net930),
    .S(_06402_),
    .X(_02241_));
 sg13g2_mux2_1 _24938_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net929),
    .S(_06402_),
    .X(_02242_));
 sg13g2_mux2_1 _24939_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(net928),
    .S(_06402_),
    .X(_02243_));
 sg13g2_and2_1 _24940_ (.A(net440),
    .B(_06287_),
    .X(_06403_));
 sg13g2_buf_2 _24941_ (.A(_06403_),
    .X(_06404_));
 sg13g2_mux2_1 _24942_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(net931),
    .S(_06404_),
    .X(_02244_));
 sg13g2_mux2_1 _24943_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net930),
    .S(_06404_),
    .X(_02245_));
 sg13g2_mux2_1 _24944_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(net929),
    .S(_06404_),
    .X(_02246_));
 sg13g2_mux2_1 _24945_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(net928),
    .S(_06404_),
    .X(_02247_));
 sg13g2_mux2_1 _24946_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net930),
    .S(_06398_),
    .X(_02248_));
 sg13g2_and2_1 _24947_ (.A(net440),
    .B(_06290_),
    .X(_06405_));
 sg13g2_buf_2 _24948_ (.A(_06405_),
    .X(_06406_));
 sg13g2_mux2_1 _24949_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net931),
    .S(_06406_),
    .X(_02249_));
 sg13g2_mux2_1 _24950_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(net930),
    .S(_06406_),
    .X(_02250_));
 sg13g2_mux2_1 _24951_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net929),
    .S(_06406_),
    .X(_02251_));
 sg13g2_mux2_1 _24952_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(_06346_),
    .S(_06406_),
    .X(_02252_));
 sg13g2_and2_1 _24953_ (.A(net440),
    .B(_06294_),
    .X(_06407_));
 sg13g2_buf_2 _24954_ (.A(_06407_),
    .X(_06408_));
 sg13g2_mux2_1 _24955_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net986),
    .S(_06408_),
    .X(_02253_));
 sg13g2_mux2_1 _24956_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net983),
    .S(_06408_),
    .X(_02254_));
 sg13g2_mux2_1 _24957_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net985),
    .S(_06408_),
    .X(_02255_));
 sg13g2_mux2_1 _24958_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net984),
    .S(_06408_),
    .X(_02256_));
 sg13g2_and2_1 _24959_ (.A(net440),
    .B(_06300_),
    .X(_06409_));
 sg13g2_buf_1 _24960_ (.A(_06409_),
    .X(_06410_));
 sg13g2_mux2_1 _24961_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net986),
    .S(_06410_),
    .X(_02257_));
 sg13g2_mux2_1 _24962_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net983),
    .S(_06410_),
    .X(_02258_));
 sg13g2_mux2_1 _24963_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net985),
    .S(_06398_),
    .X(_02259_));
 sg13g2_mux2_1 _24964_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_11938_),
    .S(_06410_),
    .X(_02260_));
 sg13g2_mux2_1 _24965_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net984),
    .S(_06410_),
    .X(_02261_));
 sg13g2_mux2_1 _24966_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_11945_),
    .S(_06398_),
    .X(_02262_));
 sg13g2_and2_1 _24967_ (.A(_08911_),
    .B(_06303_),
    .X(_06411_));
 sg13g2_buf_1 _24968_ (.A(_06411_),
    .X(_06412_));
 sg13g2_mux2_1 _24969_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_11925_),
    .S(_06412_),
    .X(_02263_));
 sg13g2_mux2_1 _24970_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_11974_),
    .S(_06412_),
    .X(_02264_));
 sg13g2_mux2_1 _24971_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_11938_),
    .S(_06412_),
    .X(_02265_));
 sg13g2_mux2_1 _24972_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_11945_),
    .S(_06412_),
    .X(_02266_));
 sg13g2_mux2_1 _24973_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_11925_),
    .S(_06400_),
    .X(_02267_));
 sg13g2_mux2_1 _24974_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_11974_),
    .S(_06400_),
    .X(_02268_));
 sg13g2_mux2_1 _24975_ (.A0(net947),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(net358),
    .X(_02272_));
 sg13g2_buf_1 _24976_ (.A(_06296_),
    .X(_06413_));
 sg13g2_nand2_1 _24977_ (.Y(_06414_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net358));
 sg13g2_o21ai_1 _24978_ (.B1(_06414_),
    .Y(_02273_),
    .A1(net382),
    .A2(net357));
 sg13g2_nand2_1 _24979_ (.Y(_06415_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net358));
 sg13g2_o21ai_1 _24980_ (.B1(_06415_),
    .Y(_02274_),
    .A1(net383),
    .A2(net357));
 sg13g2_nand2_1 _24981_ (.Y(_06416_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net358));
 sg13g2_o21ai_1 _24982_ (.B1(_06416_),
    .Y(_02275_),
    .A1(net381),
    .A2(_06413_));
 sg13g2_nand2_1 _24983_ (.Y(_06417_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net358));
 sg13g2_o21ai_1 _24984_ (.B1(_06417_),
    .Y(_02276_),
    .A1(net380),
    .A2(net357));
 sg13g2_nand2_1 _24985_ (.Y(_06418_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(net358));
 sg13g2_o21ai_1 _24986_ (.B1(_06418_),
    .Y(_02277_),
    .A1(net442),
    .A2(net357));
 sg13g2_nand2_1 _24987_ (.Y(_06419_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net358));
 sg13g2_o21ai_1 _24988_ (.B1(_06419_),
    .Y(_02278_),
    .A1(net443),
    .A2(net357));
 sg13g2_buf_1 _24989_ (.A(_06296_),
    .X(_06420_));
 sg13g2_nand2_1 _24990_ (.Y(_06421_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net356));
 sg13g2_o21ai_1 _24991_ (.B1(_06421_),
    .Y(_02279_),
    .A1(_08477_),
    .A2(net357));
 sg13g2_nand2_1 _24992_ (.Y(_06422_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net356));
 sg13g2_o21ai_1 _24993_ (.B1(_06422_),
    .Y(_02280_),
    .A1(net445),
    .A2(net357));
 sg13g2_nand2_1 _24994_ (.Y(_06423_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net356));
 sg13g2_o21ai_1 _24995_ (.B1(_06423_),
    .Y(_02281_),
    .A1(net498),
    .A2(net357));
 sg13g2_nand2_1 _24996_ (.Y(_06424_),
    .A(\cpu.icache.r_tag[0][6] ),
    .B(net356));
 sg13g2_o21ai_1 _24997_ (.B1(_06424_),
    .Y(_02282_),
    .A1(net1046),
    .A2(net359));
 sg13g2_nand2_1 _24998_ (.Y(_06425_),
    .A(\cpu.icache.r_tag[0][7] ),
    .B(net356));
 sg13g2_o21ai_1 _24999_ (.B1(_06425_),
    .Y(_02283_),
    .A1(net1045),
    .A2(net359));
 sg13g2_nand2_1 _25000_ (.Y(_06426_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(_06420_));
 sg13g2_o21ai_1 _25001_ (.B1(_06426_),
    .Y(_02284_),
    .A1(net948),
    .A2(net359));
 sg13g2_nand2_1 _25002_ (.Y(_06427_),
    .A(\cpu.icache.r_tag[0][9] ),
    .B(net356));
 sg13g2_o21ai_1 _25003_ (.B1(_06427_),
    .Y(_02285_),
    .A1(net903),
    .A2(net359));
 sg13g2_mux2_1 _25004_ (.A0(net946),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net358),
    .X(_02286_));
 sg13g2_nand2_1 _25005_ (.Y(_06428_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net356));
 sg13g2_o21ai_1 _25006_ (.B1(_06428_),
    .Y(_02287_),
    .A1(net1047),
    .A2(net359));
 sg13g2_nand2_1 _25007_ (.Y(_06429_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(net356));
 sg13g2_o21ai_1 _25008_ (.B1(_06429_),
    .Y(_02288_),
    .A1(net348),
    .A2(net359));
 sg13g2_nand2_1 _25009_ (.Y(_06430_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(_06420_));
 sg13g2_o21ai_1 _25010_ (.B1(_06430_),
    .Y(_02289_),
    .A1(net385),
    .A2(net359));
 sg13g2_nand2_1 _25011_ (.Y(_06431_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(_06296_));
 sg13g2_o21ai_1 _25012_ (.B1(_06431_),
    .Y(_02290_),
    .A1(net444),
    .A2(net359));
 sg13g2_nor3_1 _25013_ (.A(_06266_),
    .B(_06274_),
    .C(_06276_),
    .Y(_06432_));
 sg13g2_buf_1 _25014_ (.A(_06432_),
    .X(_06433_));
 sg13g2_nand2_1 _25015_ (.Y(_06434_),
    .A(_08909_),
    .B(_06433_));
 sg13g2_buf_1 _25016_ (.A(_06434_),
    .X(_06435_));
 sg13g2_buf_1 _25017_ (.A(net327),
    .X(_06436_));
 sg13g2_mux2_1 _25018_ (.A0(net947),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(net259),
    .X(_02291_));
 sg13g2_buf_1 _25019_ (.A(net327),
    .X(_06437_));
 sg13g2_nand2_1 _25020_ (.Y(_06438_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(_06436_));
 sg13g2_o21ai_1 _25021_ (.B1(_06438_),
    .Y(_02292_),
    .A1(net382),
    .A2(_06437_));
 sg13g2_buf_1 _25022_ (.A(net327),
    .X(_06439_));
 sg13g2_nand2_1 _25023_ (.Y(_06440_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net257));
 sg13g2_o21ai_1 _25024_ (.B1(_06440_),
    .Y(_02293_),
    .A1(net383),
    .A2(net258));
 sg13g2_nand2_1 _25025_ (.Y(_06441_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(_06439_));
 sg13g2_o21ai_1 _25026_ (.B1(_06441_),
    .Y(_02294_),
    .A1(net381),
    .A2(_06437_));
 sg13g2_nand2_1 _25027_ (.Y(_06442_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(_06439_));
 sg13g2_o21ai_1 _25028_ (.B1(_06442_),
    .Y(_02295_),
    .A1(net380),
    .A2(net258));
 sg13g2_nand2_1 _25029_ (.Y(_06443_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net257));
 sg13g2_o21ai_1 _25030_ (.B1(_06443_),
    .Y(_02296_),
    .A1(net442),
    .A2(net258));
 sg13g2_nand2_1 _25031_ (.Y(_06444_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net257));
 sg13g2_o21ai_1 _25032_ (.B1(_06444_),
    .Y(_02297_),
    .A1(net443),
    .A2(net258));
 sg13g2_nand2_1 _25033_ (.Y(_06445_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net257));
 sg13g2_o21ai_1 _25034_ (.B1(_06445_),
    .Y(_02298_),
    .A1(net384),
    .A2(net258));
 sg13g2_nand2_1 _25035_ (.Y(_06446_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(net257));
 sg13g2_o21ai_1 _25036_ (.B1(_06446_),
    .Y(_02299_),
    .A1(net445),
    .A2(net258));
 sg13g2_nand2_1 _25037_ (.Y(_06447_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net257));
 sg13g2_o21ai_1 _25038_ (.B1(_06447_),
    .Y(_02300_),
    .A1(net498),
    .A2(net258));
 sg13g2_nand2_1 _25039_ (.Y(_06448_),
    .A(\cpu.icache.r_tag[1][6] ),
    .B(net257));
 sg13g2_o21ai_1 _25040_ (.B1(_06448_),
    .Y(_02301_),
    .A1(net1046),
    .A2(net258));
 sg13g2_nand2_1 _25041_ (.Y(_06449_),
    .A(\cpu.icache.r_tag[1][7] ),
    .B(net257));
 sg13g2_o21ai_1 _25042_ (.B1(_06449_),
    .Y(_02302_),
    .A1(net1045),
    .A2(net259));
 sg13g2_nand2_1 _25043_ (.Y(_06450_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net327));
 sg13g2_o21ai_1 _25044_ (.B1(_06450_),
    .Y(_02303_),
    .A1(net948),
    .A2(net259));
 sg13g2_nand2_1 _25045_ (.Y(_06451_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(net327));
 sg13g2_o21ai_1 _25046_ (.B1(_06451_),
    .Y(_02304_),
    .A1(net903),
    .A2(net259));
 sg13g2_mux2_1 _25047_ (.A0(net946),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net259),
    .X(_02305_));
 sg13g2_nand2_1 _25048_ (.Y(_06452_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(net327));
 sg13g2_o21ai_1 _25049_ (.B1(_06452_),
    .Y(_02306_),
    .A1(net1047),
    .A2(net259));
 sg13g2_nand2_1 _25050_ (.Y(_06453_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(net327));
 sg13g2_o21ai_1 _25051_ (.B1(_06453_),
    .Y(_02307_),
    .A1(net348),
    .A2(net259));
 sg13g2_nand2_1 _25052_ (.Y(_06454_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(net327));
 sg13g2_o21ai_1 _25053_ (.B1(_06454_),
    .Y(_02308_),
    .A1(net385),
    .A2(net259));
 sg13g2_nand2_1 _25054_ (.Y(_06455_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06435_));
 sg13g2_o21ai_1 _25055_ (.B1(_06455_),
    .Y(_02309_),
    .A1(net444),
    .A2(_06436_));
 sg13g2_nand2_1 _25056_ (.Y(_06456_),
    .A(_08908_),
    .B(_06433_));
 sg13g2_buf_1 _25057_ (.A(_06456_),
    .X(_06457_));
 sg13g2_buf_1 _25058_ (.A(net256),
    .X(_06458_));
 sg13g2_mux2_1 _25059_ (.A0(net947),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net219),
    .X(_02310_));
 sg13g2_buf_1 _25060_ (.A(net256),
    .X(_06459_));
 sg13g2_nand2_1 _25061_ (.Y(_06460_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net219));
 sg13g2_o21ai_1 _25062_ (.B1(_06460_),
    .Y(_02311_),
    .A1(net382),
    .A2(net218));
 sg13g2_buf_1 _25063_ (.A(net256),
    .X(_06461_));
 sg13g2_nand2_1 _25064_ (.Y(_06462_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net217));
 sg13g2_o21ai_1 _25065_ (.B1(_06462_),
    .Y(_02312_),
    .A1(net383),
    .A2(net218));
 sg13g2_nand2_1 _25066_ (.Y(_06463_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net217));
 sg13g2_o21ai_1 _25067_ (.B1(_06463_),
    .Y(_02313_),
    .A1(net381),
    .A2(net218));
 sg13g2_nand2_1 _25068_ (.Y(_06464_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net217));
 sg13g2_o21ai_1 _25069_ (.B1(_06464_),
    .Y(_02314_),
    .A1(net380),
    .A2(_06459_));
 sg13g2_nand2_1 _25070_ (.Y(_06465_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net217));
 sg13g2_o21ai_1 _25071_ (.B1(_06465_),
    .Y(_02315_),
    .A1(net442),
    .A2(net218));
 sg13g2_nand2_1 _25072_ (.Y(_06466_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net217));
 sg13g2_o21ai_1 _25073_ (.B1(_06466_),
    .Y(_02316_),
    .A1(net443),
    .A2(net218));
 sg13g2_nand2_1 _25074_ (.Y(_06467_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(_06461_));
 sg13g2_o21ai_1 _25075_ (.B1(_06467_),
    .Y(_02317_),
    .A1(net384),
    .A2(_06459_));
 sg13g2_nand2_1 _25076_ (.Y(_06468_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(net217));
 sg13g2_o21ai_1 _25077_ (.B1(_06468_),
    .Y(_02318_),
    .A1(net445),
    .A2(net218));
 sg13g2_nand2_1 _25078_ (.Y(_06469_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(_06461_));
 sg13g2_o21ai_1 _25079_ (.B1(_06469_),
    .Y(_02319_),
    .A1(net498),
    .A2(net218));
 sg13g2_nand2_1 _25080_ (.Y(_06470_),
    .A(\cpu.icache.r_tag[2][6] ),
    .B(net217));
 sg13g2_o21ai_1 _25081_ (.B1(_06470_),
    .Y(_02320_),
    .A1(net1046),
    .A2(net218));
 sg13g2_nand2_1 _25082_ (.Y(_06471_),
    .A(\cpu.icache.r_tag[2][7] ),
    .B(net217));
 sg13g2_o21ai_1 _25083_ (.B1(_06471_),
    .Y(_02321_),
    .A1(net1045),
    .A2(net219));
 sg13g2_nand2_1 _25084_ (.Y(_06472_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(_06457_));
 sg13g2_o21ai_1 _25085_ (.B1(_06472_),
    .Y(_02322_),
    .A1(net948),
    .A2(net219));
 sg13g2_nand2_1 _25086_ (.Y(_06473_),
    .A(\cpu.icache.r_tag[2][9] ),
    .B(net256));
 sg13g2_o21ai_1 _25087_ (.B1(_06473_),
    .Y(_02323_),
    .A1(net903),
    .A2(net219));
 sg13g2_mux2_1 _25088_ (.A0(net946),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net219),
    .X(_02324_));
 sg13g2_nand2_1 _25089_ (.Y(_06474_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(net256));
 sg13g2_o21ai_1 _25090_ (.B1(_06474_),
    .Y(_02325_),
    .A1(net1047),
    .A2(net219));
 sg13g2_nand2_1 _25091_ (.Y(_06475_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(net256));
 sg13g2_o21ai_1 _25092_ (.B1(_06475_),
    .Y(_02326_),
    .A1(net348),
    .A2(_06458_));
 sg13g2_nand2_1 _25093_ (.Y(_06476_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(net256));
 sg13g2_o21ai_1 _25094_ (.B1(_06476_),
    .Y(_02327_),
    .A1(net385),
    .A2(_06458_));
 sg13g2_nand2_1 _25095_ (.Y(_06477_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(net256));
 sg13g2_o21ai_1 _25096_ (.B1(_06477_),
    .Y(_02328_),
    .A1(net444),
    .A2(net219));
 sg13g2_mux2_1 _25097_ (.A0(net947),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net220),
    .X(_02329_));
 sg13g2_buf_1 _25098_ (.A(_06360_),
    .X(_06478_));
 sg13g2_nand2_1 _25099_ (.Y(_06479_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net220));
 sg13g2_o21ai_1 _25100_ (.B1(_06479_),
    .Y(_02330_),
    .A1(net382),
    .A2(net216));
 sg13g2_nand2_1 _25101_ (.Y(_06480_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net220));
 sg13g2_o21ai_1 _25102_ (.B1(_06480_),
    .Y(_02331_),
    .A1(net383),
    .A2(net216));
 sg13g2_nand2_1 _25103_ (.Y(_06481_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(_06362_));
 sg13g2_o21ai_1 _25104_ (.B1(_06481_),
    .Y(_02332_),
    .A1(net381),
    .A2(_06478_));
 sg13g2_nand2_1 _25105_ (.Y(_06482_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(_06362_));
 sg13g2_o21ai_1 _25106_ (.B1(_06482_),
    .Y(_02333_),
    .A1(_08564_),
    .A2(_06478_));
 sg13g2_nand2_1 _25107_ (.Y(_06483_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net220));
 sg13g2_o21ai_1 _25108_ (.B1(_06483_),
    .Y(_02334_),
    .A1(net442),
    .A2(net216));
 sg13g2_nand2_1 _25109_ (.Y(_06484_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net220));
 sg13g2_o21ai_1 _25110_ (.B1(_06484_),
    .Y(_02335_),
    .A1(net443),
    .A2(net216));
 sg13g2_buf_1 _25111_ (.A(_06360_),
    .X(_06485_));
 sg13g2_nand2_1 _25112_ (.Y(_06486_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net215));
 sg13g2_o21ai_1 _25113_ (.B1(_06486_),
    .Y(_02336_),
    .A1(net384),
    .A2(net216));
 sg13g2_nand2_1 _25114_ (.Y(_06487_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(net215));
 sg13g2_o21ai_1 _25115_ (.B1(_06487_),
    .Y(_02337_),
    .A1(net445),
    .A2(net216));
 sg13g2_nand2_1 _25116_ (.Y(_06488_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net215));
 sg13g2_o21ai_1 _25117_ (.B1(_06488_),
    .Y(_02338_),
    .A1(net498),
    .A2(net216));
 sg13g2_nand2_1 _25118_ (.Y(_06489_),
    .A(\cpu.icache.r_tag[3][6] ),
    .B(net215));
 sg13g2_o21ai_1 _25119_ (.B1(_06489_),
    .Y(_02339_),
    .A1(net1046),
    .A2(net221));
 sg13g2_nand2_1 _25120_ (.Y(_06490_),
    .A(\cpu.icache.r_tag[3][7] ),
    .B(net215));
 sg13g2_o21ai_1 _25121_ (.B1(_06490_),
    .Y(_02340_),
    .A1(_08680_),
    .A2(net221));
 sg13g2_nand2_1 _25122_ (.Y(_06491_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(net215));
 sg13g2_o21ai_1 _25123_ (.B1(_06491_),
    .Y(_02341_),
    .A1(net948),
    .A2(net221));
 sg13g2_nand2_1 _25124_ (.Y(_06492_),
    .A(\cpu.icache.r_tag[3][9] ),
    .B(net215));
 sg13g2_o21ai_1 _25125_ (.B1(_06492_),
    .Y(_02342_),
    .A1(net903),
    .A2(net221));
 sg13g2_mux2_1 _25126_ (.A0(net946),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net220),
    .X(_02343_));
 sg13g2_nand2_1 _25127_ (.Y(_06493_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(_06485_));
 sg13g2_o21ai_1 _25128_ (.B1(_06493_),
    .Y(_02344_),
    .A1(net1047),
    .A2(net221));
 sg13g2_nand2_1 _25129_ (.Y(_06494_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(_06485_));
 sg13g2_o21ai_1 _25130_ (.B1(_06494_),
    .Y(_02345_),
    .A1(net348),
    .A2(_06361_));
 sg13g2_nand2_1 _25131_ (.Y(_06495_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(net215));
 sg13g2_o21ai_1 _25132_ (.B1(_06495_),
    .Y(_02346_),
    .A1(net385),
    .A2(net221));
 sg13g2_nand2_1 _25133_ (.Y(_06496_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(_06360_));
 sg13g2_o21ai_1 _25134_ (.B1(_06496_),
    .Y(_02347_),
    .A1(net444),
    .A2(net221));
 sg13g2_nand2_1 _25135_ (.Y(_06497_),
    .A(net554),
    .B(_06433_));
 sg13g2_buf_1 _25136_ (.A(_06497_),
    .X(_06498_));
 sg13g2_buf_1 _25137_ (.A(net391),
    .X(_06499_));
 sg13g2_mux2_1 _25138_ (.A0(net947),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net355),
    .X(_02348_));
 sg13g2_buf_1 _25139_ (.A(net391),
    .X(_06500_));
 sg13g2_nand2_1 _25140_ (.Y(_06501_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net355));
 sg13g2_o21ai_1 _25141_ (.B1(_06501_),
    .Y(_02349_),
    .A1(net382),
    .A2(net354));
 sg13g2_buf_1 _25142_ (.A(_06498_),
    .X(_06502_));
 sg13g2_nand2_1 _25143_ (.Y(_06503_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net353));
 sg13g2_o21ai_1 _25144_ (.B1(_06503_),
    .Y(_02350_),
    .A1(net383),
    .A2(net354));
 sg13g2_nand2_1 _25145_ (.Y(_06504_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net353));
 sg13g2_o21ai_1 _25146_ (.B1(_06504_),
    .Y(_02351_),
    .A1(net381),
    .A2(net354));
 sg13g2_nand2_1 _25147_ (.Y(_06505_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net353));
 sg13g2_o21ai_1 _25148_ (.B1(_06505_),
    .Y(_02352_),
    .A1(net380),
    .A2(net354));
 sg13g2_nand2_1 _25149_ (.Y(_06506_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net353));
 sg13g2_o21ai_1 _25150_ (.B1(_06506_),
    .Y(_02353_),
    .A1(net442),
    .A2(net354));
 sg13g2_nand2_1 _25151_ (.Y(_06507_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net353));
 sg13g2_o21ai_1 _25152_ (.B1(_06507_),
    .Y(_02354_),
    .A1(net443),
    .A2(net354));
 sg13g2_nand2_1 _25153_ (.Y(_06508_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(_06502_));
 sg13g2_o21ai_1 _25154_ (.B1(_06508_),
    .Y(_02355_),
    .A1(net384),
    .A2(_06500_));
 sg13g2_nand2_1 _25155_ (.Y(_06509_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net353));
 sg13g2_o21ai_1 _25156_ (.B1(_06509_),
    .Y(_02356_),
    .A1(net445),
    .A2(net354));
 sg13g2_nand2_1 _25157_ (.Y(_06510_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(_06502_));
 sg13g2_o21ai_1 _25158_ (.B1(_06510_),
    .Y(_02357_),
    .A1(net498),
    .A2(_06500_));
 sg13g2_nand2_1 _25159_ (.Y(_06511_),
    .A(\cpu.icache.r_tag[4][6] ),
    .B(net353));
 sg13g2_o21ai_1 _25160_ (.B1(_06511_),
    .Y(_02358_),
    .A1(net1046),
    .A2(net354));
 sg13g2_nand2_1 _25161_ (.Y(_06512_),
    .A(\cpu.icache.r_tag[4][7] ),
    .B(net353));
 sg13g2_o21ai_1 _25162_ (.B1(_06512_),
    .Y(_02359_),
    .A1(net1045),
    .A2(net355));
 sg13g2_nand2_1 _25163_ (.Y(_06513_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(net391));
 sg13g2_o21ai_1 _25164_ (.B1(_06513_),
    .Y(_02360_),
    .A1(net948),
    .A2(net355));
 sg13g2_nand2_1 _25165_ (.Y(_06514_),
    .A(\cpu.icache.r_tag[4][9] ),
    .B(net391));
 sg13g2_o21ai_1 _25166_ (.B1(_06514_),
    .Y(_02361_),
    .A1(net903),
    .A2(_06499_));
 sg13g2_mux2_1 _25167_ (.A0(net946),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net355),
    .X(_02362_));
 sg13g2_nand2_1 _25168_ (.Y(_06515_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(net391));
 sg13g2_o21ai_1 _25169_ (.B1(_06515_),
    .Y(_02363_),
    .A1(net1047),
    .A2(net355));
 sg13g2_nand2_1 _25170_ (.Y(_06516_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(net391));
 sg13g2_o21ai_1 _25171_ (.B1(_06516_),
    .Y(_02364_),
    .A1(net348),
    .A2(_06499_));
 sg13g2_nand2_1 _25172_ (.Y(_06517_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(net391));
 sg13g2_o21ai_1 _25173_ (.B1(_06517_),
    .Y(_02365_),
    .A1(net385),
    .A2(net355));
 sg13g2_nand2_1 _25174_ (.Y(_06518_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(net391));
 sg13g2_o21ai_1 _25175_ (.B1(_06518_),
    .Y(_02366_),
    .A1(_08607_),
    .A2(net355));
 sg13g2_nand2_1 _25176_ (.Y(_06519_),
    .A(net446),
    .B(_06433_));
 sg13g2_buf_1 _25177_ (.A(_06519_),
    .X(_06520_));
 sg13g2_buf_1 _25178_ (.A(_06520_),
    .X(_06521_));
 sg13g2_mux2_1 _25179_ (.A0(net947),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net255),
    .X(_02367_));
 sg13g2_buf_1 _25180_ (.A(net326),
    .X(_06522_));
 sg13g2_nand2_1 _25181_ (.Y(_06523_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(_06521_));
 sg13g2_o21ai_1 _25182_ (.B1(_06523_),
    .Y(_02368_),
    .A1(net382),
    .A2(_06522_));
 sg13g2_buf_1 _25183_ (.A(net326),
    .X(_06524_));
 sg13g2_nand2_1 _25184_ (.Y(_06525_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net253));
 sg13g2_o21ai_1 _25185_ (.B1(_06525_),
    .Y(_02369_),
    .A1(net383),
    .A2(net254));
 sg13g2_nand2_1 _25186_ (.Y(_06526_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net253));
 sg13g2_o21ai_1 _25187_ (.B1(_06526_),
    .Y(_02370_),
    .A1(net381),
    .A2(net254));
 sg13g2_nand2_1 _25188_ (.Y(_06527_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(_06524_));
 sg13g2_o21ai_1 _25189_ (.B1(_06527_),
    .Y(_02371_),
    .A1(net380),
    .A2(net254));
 sg13g2_nand2_1 _25190_ (.Y(_06528_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net253));
 sg13g2_o21ai_1 _25191_ (.B1(_06528_),
    .Y(_02372_),
    .A1(net442),
    .A2(net254));
 sg13g2_nand2_1 _25192_ (.Y(_06529_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(net253));
 sg13g2_o21ai_1 _25193_ (.B1(_06529_),
    .Y(_02373_),
    .A1(_08628_),
    .A2(net254));
 sg13g2_nand2_1 _25194_ (.Y(_06530_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(net253));
 sg13g2_o21ai_1 _25195_ (.B1(_06530_),
    .Y(_02374_),
    .A1(net384),
    .A2(net254));
 sg13g2_nand2_1 _25196_ (.Y(_06531_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(net253));
 sg13g2_o21ai_1 _25197_ (.B1(_06531_),
    .Y(_02375_),
    .A1(net445),
    .A2(net254));
 sg13g2_nand2_1 _25198_ (.Y(_06532_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net253));
 sg13g2_o21ai_1 _25199_ (.B1(_06532_),
    .Y(_02376_),
    .A1(net498),
    .A2(net254));
 sg13g2_nand2_1 _25200_ (.Y(_06533_),
    .A(\cpu.icache.r_tag[5][6] ),
    .B(_06524_));
 sg13g2_o21ai_1 _25201_ (.B1(_06533_),
    .Y(_02377_),
    .A1(_08670_),
    .A2(_06522_));
 sg13g2_nand2_1 _25202_ (.Y(_06534_),
    .A(\cpu.icache.r_tag[5][7] ),
    .B(net253));
 sg13g2_o21ai_1 _25203_ (.B1(_06534_),
    .Y(_02378_),
    .A1(net1045),
    .A2(net255));
 sg13g2_nand2_1 _25204_ (.Y(_06535_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net326));
 sg13g2_o21ai_1 _25205_ (.B1(_06535_),
    .Y(_02379_),
    .A1(net948),
    .A2(net255));
 sg13g2_nand2_1 _25206_ (.Y(_06536_),
    .A(\cpu.icache.r_tag[5][9] ),
    .B(net326));
 sg13g2_o21ai_1 _25207_ (.B1(_06536_),
    .Y(_02380_),
    .A1(net903),
    .A2(net255));
 sg13g2_mux2_1 _25208_ (.A0(net946),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net255),
    .X(_02381_));
 sg13g2_nand2_1 _25209_ (.Y(_06537_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(net326));
 sg13g2_o21ai_1 _25210_ (.B1(_06537_),
    .Y(_02382_),
    .A1(_08659_),
    .A2(net255));
 sg13g2_nand2_1 _25211_ (.Y(_06538_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(net326));
 sg13g2_o21ai_1 _25212_ (.B1(_06538_),
    .Y(_02383_),
    .A1(net348),
    .A2(net255));
 sg13g2_nand2_1 _25213_ (.Y(_06539_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(net326));
 sg13g2_o21ai_1 _25214_ (.B1(_06539_),
    .Y(_02384_),
    .A1(_08426_),
    .A2(net255));
 sg13g2_nand2_1 _25215_ (.Y(_06540_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(net326));
 sg13g2_o21ai_1 _25216_ (.B1(_06540_),
    .Y(_02385_),
    .A1(net444),
    .A2(_06521_));
 sg13g2_nand2_1 _25217_ (.Y(_06541_),
    .A(net553),
    .B(_06433_));
 sg13g2_buf_1 _25218_ (.A(_06541_),
    .X(_06542_));
 sg13g2_buf_1 _25219_ (.A(_06542_),
    .X(_06543_));
 sg13g2_mux2_1 _25220_ (.A0(_04570_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net352),
    .X(_02386_));
 sg13g2_buf_1 _25221_ (.A(net390),
    .X(_06544_));
 sg13g2_nand2_1 _25222_ (.Y(_06545_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net352));
 sg13g2_o21ai_1 _25223_ (.B1(_06545_),
    .Y(_02387_),
    .A1(net382),
    .A2(net351));
 sg13g2_buf_1 _25224_ (.A(net390),
    .X(_06546_));
 sg13g2_nand2_1 _25225_ (.Y(_06547_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net350));
 sg13g2_o21ai_1 _25226_ (.B1(_06547_),
    .Y(_02388_),
    .A1(net383),
    .A2(net351));
 sg13g2_nand2_1 _25227_ (.Y(_06548_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net350));
 sg13g2_o21ai_1 _25228_ (.B1(_06548_),
    .Y(_02389_),
    .A1(net381),
    .A2(net351));
 sg13g2_nand2_1 _25229_ (.Y(_06549_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net350));
 sg13g2_o21ai_1 _25230_ (.B1(_06549_),
    .Y(_02390_),
    .A1(net380),
    .A2(net351));
 sg13g2_nand2_1 _25231_ (.Y(_06550_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net350));
 sg13g2_o21ai_1 _25232_ (.B1(_06550_),
    .Y(_02391_),
    .A1(net442),
    .A2(net351));
 sg13g2_nand2_1 _25233_ (.Y(_06551_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(net350));
 sg13g2_o21ai_1 _25234_ (.B1(_06551_),
    .Y(_02392_),
    .A1(net443),
    .A2(net351));
 sg13g2_nand2_1 _25235_ (.Y(_06552_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(_06546_));
 sg13g2_o21ai_1 _25236_ (.B1(_06552_),
    .Y(_02393_),
    .A1(net384),
    .A2(_06544_));
 sg13g2_nand2_1 _25237_ (.Y(_06553_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net350));
 sg13g2_o21ai_1 _25238_ (.B1(_06553_),
    .Y(_02394_),
    .A1(_08585_),
    .A2(net351));
 sg13g2_nand2_1 _25239_ (.Y(_06554_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(_06546_));
 sg13g2_o21ai_1 _25240_ (.B1(_06554_),
    .Y(_02395_),
    .A1(net498),
    .A2(_06544_));
 sg13g2_nand2_1 _25241_ (.Y(_06555_),
    .A(\cpu.icache.r_tag[6][6] ),
    .B(net350));
 sg13g2_o21ai_1 _25242_ (.B1(_06555_),
    .Y(_02396_),
    .A1(net1046),
    .A2(net351));
 sg13g2_nand2_1 _25243_ (.Y(_06556_),
    .A(\cpu.icache.r_tag[6][7] ),
    .B(net350));
 sg13g2_o21ai_1 _25244_ (.B1(_06556_),
    .Y(_02397_),
    .A1(net1045),
    .A2(net352));
 sg13g2_nand2_1 _25245_ (.Y(_06557_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(net390));
 sg13g2_o21ai_1 _25246_ (.B1(_06557_),
    .Y(_02398_),
    .A1(_04212_),
    .A2(net352));
 sg13g2_nand2_1 _25247_ (.Y(_06558_),
    .A(\cpu.icache.r_tag[6][9] ),
    .B(net390));
 sg13g2_o21ai_1 _25248_ (.B1(_06558_),
    .Y(_02399_),
    .A1(net903),
    .A2(_06543_));
 sg13g2_mux2_1 _25249_ (.A0(_04720_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net352),
    .X(_02400_));
 sg13g2_nand2_1 _25250_ (.Y(_06559_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(net390));
 sg13g2_o21ai_1 _25251_ (.B1(_06559_),
    .Y(_02401_),
    .A1(net1047),
    .A2(_06543_));
 sg13g2_nand2_1 _25252_ (.Y(_06560_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(net390));
 sg13g2_o21ai_1 _25253_ (.B1(_06560_),
    .Y(_02402_),
    .A1(net348),
    .A2(net352));
 sg13g2_nand2_1 _25254_ (.Y(_06561_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(net390));
 sg13g2_o21ai_1 _25255_ (.B1(_06561_),
    .Y(_02403_),
    .A1(net385),
    .A2(net352));
 sg13g2_nand2_1 _25256_ (.Y(_06562_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(net390));
 sg13g2_o21ai_1 _25257_ (.B1(_06562_),
    .Y(_02404_),
    .A1(net444),
    .A2(net352));
 sg13g2_nand2_1 _25258_ (.Y(_06563_),
    .A(_08911_),
    .B(_06433_));
 sg13g2_buf_1 _25259_ (.A(_06563_),
    .X(_06564_));
 sg13g2_buf_1 _25260_ (.A(net325),
    .X(_06565_));
 sg13g2_mux2_1 _25261_ (.A0(_04570_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net252),
    .X(_02405_));
 sg13g2_buf_1 _25262_ (.A(net325),
    .X(_06566_));
 sg13g2_nand2_1 _25263_ (.Y(_06567_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(_06565_));
 sg13g2_o21ai_1 _25264_ (.B1(_06567_),
    .Y(_02406_),
    .A1(_08522_),
    .A2(net251));
 sg13g2_buf_1 _25265_ (.A(net325),
    .X(_06568_));
 sg13g2_nand2_1 _25266_ (.Y(_06569_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net250));
 sg13g2_o21ai_1 _25267_ (.B1(_06569_),
    .Y(_02407_),
    .A1(net383),
    .A2(net251));
 sg13g2_nand2_1 _25268_ (.Y(_06570_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net250));
 sg13g2_o21ai_1 _25269_ (.B1(_06570_),
    .Y(_02408_),
    .A1(_08543_),
    .A2(_06566_));
 sg13g2_nand2_1 _25270_ (.Y(_06571_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(net250));
 sg13g2_o21ai_1 _25271_ (.B1(_06571_),
    .Y(_02409_),
    .A1(net380),
    .A2(net251));
 sg13g2_nand2_1 _25272_ (.Y(_06572_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net250));
 sg13g2_o21ai_1 _25273_ (.B1(_06572_),
    .Y(_02410_),
    .A1(net442),
    .A2(net251));
 sg13g2_nand2_1 _25274_ (.Y(_06573_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(_06568_));
 sg13g2_o21ai_1 _25275_ (.B1(_06573_),
    .Y(_02411_),
    .A1(net443),
    .A2(net251));
 sg13g2_nand2_1 _25276_ (.Y(_06574_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net250));
 sg13g2_o21ai_1 _25277_ (.B1(_06574_),
    .Y(_02412_),
    .A1(net384),
    .A2(net251));
 sg13g2_nand2_1 _25278_ (.Y(_06575_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(_06568_));
 sg13g2_o21ai_1 _25279_ (.B1(_06575_),
    .Y(_02413_),
    .A1(net445),
    .A2(_06566_));
 sg13g2_nand2_1 _25280_ (.Y(_06576_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net250));
 sg13g2_o21ai_1 _25281_ (.B1(_06576_),
    .Y(_02414_),
    .A1(_08450_),
    .A2(net251));
 sg13g2_nand2_1 _25282_ (.Y(_06577_),
    .A(\cpu.icache.r_tag[7][6] ),
    .B(net250));
 sg13g2_o21ai_1 _25283_ (.B1(_06577_),
    .Y(_02415_),
    .A1(net1046),
    .A2(net251));
 sg13g2_nand2_1 _25284_ (.Y(_06578_),
    .A(\cpu.icache.r_tag[7][7] ),
    .B(net250));
 sg13g2_o21ai_1 _25285_ (.B1(_06578_),
    .Y(_02416_),
    .A1(net1045),
    .A2(net252));
 sg13g2_nand2_1 _25286_ (.Y(_06579_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net325));
 sg13g2_o21ai_1 _25287_ (.B1(_06579_),
    .Y(_02417_),
    .A1(_04212_),
    .A2(net252));
 sg13g2_nand2_1 _25288_ (.Y(_06580_),
    .A(\cpu.icache.r_tag[7][9] ),
    .B(net325));
 sg13g2_o21ai_1 _25289_ (.B1(_06580_),
    .Y(_02418_),
    .A1(_08721_),
    .A2(net252));
 sg13g2_mux2_1 _25290_ (.A0(_04720_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net252),
    .X(_02419_));
 sg13g2_nand2_1 _25291_ (.Y(_06581_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(net325));
 sg13g2_o21ai_1 _25292_ (.B1(_06581_),
    .Y(_02420_),
    .A1(net1047),
    .A2(net252));
 sg13g2_nand2_1 _25293_ (.Y(_06582_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(net325));
 sg13g2_o21ai_1 _25294_ (.B1(_06582_),
    .Y(_02421_),
    .A1(_08401_),
    .A2(net252));
 sg13g2_nand2_1 _25295_ (.Y(_06583_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(net325));
 sg13g2_o21ai_1 _25296_ (.B1(_06583_),
    .Y(_02422_),
    .A1(net385),
    .A2(net252));
 sg13g2_nand2_1 _25297_ (.Y(_06584_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06564_));
 sg13g2_o21ai_1 _25298_ (.B1(_06584_),
    .Y(_02423_),
    .A1(net444),
    .A2(_06565_));
 sg13g2_and2_1 _25299_ (.A(_09957_),
    .B(net458),
    .X(_06585_));
 sg13g2_buf_2 _25300_ (.A(_06585_),
    .X(_06586_));
 sg13g2_buf_1 _25301_ (.A(_06586_),
    .X(_06587_));
 sg13g2_mux2_1 _25302_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(net861),
    .S(net75),
    .X(_02433_));
 sg13g2_mux2_1 _25303_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(_10018_),
    .S(net75),
    .X(_02434_));
 sg13g2_mux2_1 _25304_ (.A0(\cpu.intr.r_clock_cmp[11] ),
    .A1(_10025_),
    .S(net75),
    .X(_02435_));
 sg13g2_mux2_1 _25305_ (.A0(\cpu.intr.r_clock_cmp[12] ),
    .A1(_10030_),
    .S(net75),
    .X(_02436_));
 sg13g2_mux2_1 _25306_ (.A0(\cpu.intr.r_clock_cmp[13] ),
    .A1(_10036_),
    .S(net75),
    .X(_02437_));
 sg13g2_mux2_1 _25307_ (.A0(\cpu.intr.r_clock_cmp[14] ),
    .A1(_10043_),
    .S(_06587_),
    .X(_02438_));
 sg13g2_mux2_1 _25308_ (.A0(\cpu.intr.r_clock_cmp[15] ),
    .A1(_10048_),
    .S(_06587_),
    .X(_02439_));
 sg13g2_nor3_1 _25309_ (.A(_09109_),
    .B(_09821_),
    .C(_05421_),
    .Y(_06588_));
 sg13g2_buf_2 _25310_ (.A(_06588_),
    .X(_06589_));
 sg13g2_buf_1 _25311_ (.A(_06589_),
    .X(_06590_));
 sg13g2_mux2_1 _25312_ (.A0(\cpu.intr.r_clock_cmp[16] ),
    .A1(net861),
    .S(net96),
    .X(_02440_));
 sg13g2_mux2_1 _25313_ (.A0(\cpu.intr.r_clock_cmp[17] ),
    .A1(net883),
    .S(net96),
    .X(_02441_));
 sg13g2_mux2_1 _25314_ (.A0(\cpu.intr.r_clock_cmp[18] ),
    .A1(net862),
    .S(net96),
    .X(_02442_));
 sg13g2_mux2_1 _25315_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(net990),
    .S(net96),
    .X(_02443_));
 sg13g2_mux2_1 _25316_ (.A0(\cpu.intr.r_clock_cmp[1] ),
    .A1(net859),
    .S(net75),
    .X(_02444_));
 sg13g2_mux2_1 _25317_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(net981),
    .S(net96),
    .X(_02445_));
 sg13g2_mux2_1 _25318_ (.A0(\cpu.intr.r_clock_cmp[21] ),
    .A1(net980),
    .S(net96),
    .X(_02446_));
 sg13g2_mux2_1 _25319_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(net979),
    .S(net96),
    .X(_02447_));
 sg13g2_mux2_1 _25320_ (.A0(\cpu.intr.r_clock_cmp[23] ),
    .A1(net978),
    .S(net96),
    .X(_02448_));
 sg13g2_mux2_1 _25321_ (.A0(\cpu.intr.r_clock_cmp[24] ),
    .A1(_10008_),
    .S(_06590_),
    .X(_02449_));
 sg13g2_mux2_1 _25322_ (.A0(\cpu.intr.r_clock_cmp[25] ),
    .A1(_10013_),
    .S(_06590_),
    .X(_02450_));
 sg13g2_mux2_1 _25323_ (.A0(\cpu.intr.r_clock_cmp[26] ),
    .A1(_10018_),
    .S(_06589_),
    .X(_02451_));
 sg13g2_mux2_1 _25324_ (.A0(\cpu.intr.r_clock_cmp[27] ),
    .A1(_10025_),
    .S(_06589_),
    .X(_02452_));
 sg13g2_mux2_1 _25325_ (.A0(\cpu.intr.r_clock_cmp[28] ),
    .A1(_10030_),
    .S(_06589_),
    .X(_02453_));
 sg13g2_mux2_1 _25326_ (.A0(\cpu.intr.r_clock_cmp[29] ),
    .A1(_10036_),
    .S(_06589_),
    .X(_02454_));
 sg13g2_mux2_1 _25327_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(net858),
    .S(net75),
    .X(_02455_));
 sg13g2_mux2_1 _25328_ (.A0(\cpu.intr.r_clock_cmp[30] ),
    .A1(_10043_),
    .S(_06589_),
    .X(_02456_));
 sg13g2_mux2_1 _25329_ (.A0(\cpu.intr.r_clock_cmp[31] ),
    .A1(_10048_),
    .S(_06589_),
    .X(_02457_));
 sg13g2_mux2_1 _25330_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(net990),
    .S(net75),
    .X(_02458_));
 sg13g2_mux2_1 _25331_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(net981),
    .S(_06586_),
    .X(_02459_));
 sg13g2_mux2_1 _25332_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(net980),
    .S(_06586_),
    .X(_02460_));
 sg13g2_mux2_1 _25333_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(_12002_),
    .S(_06586_),
    .X(_02461_));
 sg13g2_mux2_1 _25334_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(net978),
    .S(_06586_),
    .X(_02462_));
 sg13g2_mux2_1 _25335_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(_10008_),
    .S(_06586_),
    .X(_02463_));
 sg13g2_mux2_1 _25336_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(_10013_),
    .S(_06586_),
    .X(_02464_));
 sg13g2_and2_1 _25337_ (.A(net123),
    .B(net361),
    .X(_06591_));
 sg13g2_buf_2 _25338_ (.A(_06591_),
    .X(_06592_));
 sg13g2_buf_1 _25339_ (.A(_06592_),
    .X(_06593_));
 sg13g2_mux2_1 _25340_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(net861),
    .S(net74),
    .X(_02488_));
 sg13g2_mux2_1 _25341_ (.A0(\cpu.intr.r_timer_reload[10] ),
    .A1(_10018_),
    .S(net74),
    .X(_02489_));
 sg13g2_mux2_1 _25342_ (.A0(\cpu.intr.r_timer_reload[11] ),
    .A1(_10025_),
    .S(net74),
    .X(_02490_));
 sg13g2_mux2_1 _25343_ (.A0(\cpu.intr.r_timer_reload[12] ),
    .A1(_10030_),
    .S(net74),
    .X(_02491_));
 sg13g2_mux2_1 _25344_ (.A0(\cpu.intr.r_timer_reload[13] ),
    .A1(_10036_),
    .S(net74),
    .X(_02492_));
 sg13g2_mux2_1 _25345_ (.A0(\cpu.intr.r_timer_reload[14] ),
    .A1(_10043_),
    .S(_06593_),
    .X(_02493_));
 sg13g2_mux2_1 _25346_ (.A0(\cpu.intr.r_timer_reload[15] ),
    .A1(_10048_),
    .S(_06593_),
    .X(_02494_));
 sg13g2_mux2_1 _25347_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net861),
    .S(net105),
    .X(_02495_));
 sg13g2_inv_1 _25348_ (.Y(_06594_),
    .A(\cpu.intr.r_timer_reload[17] ));
 sg13g2_o21ai_1 _25349_ (.B1(_09906_),
    .Y(_02496_),
    .A1(_06594_),
    .A2(net104));
 sg13g2_inv_1 _25350_ (.Y(_06595_),
    .A(\cpu.intr.r_timer_reload[18] ));
 sg13g2_o21ai_1 _25351_ (.B1(_09911_),
    .Y(_02497_),
    .A1(_06595_),
    .A2(net104));
 sg13g2_inv_1 _25352_ (.Y(_06596_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25353_ (.B1(_09917_),
    .Y(_02498_),
    .A1(_06596_),
    .A2(net104));
 sg13g2_mux2_1 _25354_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(net859),
    .S(net74),
    .X(_02499_));
 sg13g2_inv_1 _25355_ (.Y(_06597_),
    .A(\cpu.intr.r_timer_reload[20] ));
 sg13g2_o21ai_1 _25356_ (.B1(_09923_),
    .Y(_02500_),
    .A1(_06597_),
    .A2(net104));
 sg13g2_inv_1 _25357_ (.Y(_06598_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25358_ (.B1(_09929_),
    .Y(_02501_),
    .A1(_06598_),
    .A2(_09899_));
 sg13g2_inv_1 _25359_ (.Y(_06599_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25360_ (.B1(_09935_),
    .Y(_02502_),
    .A1(_06599_),
    .A2(_09899_));
 sg13g2_mux2_1 _25361_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net978),
    .S(net105),
    .X(_02503_));
 sg13g2_mux2_1 _25362_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(net858),
    .S(net74),
    .X(_02504_));
 sg13g2_mux2_1 _25363_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(net990),
    .S(net74),
    .X(_02505_));
 sg13g2_mux2_1 _25364_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(net981),
    .S(_06592_),
    .X(_02506_));
 sg13g2_mux2_1 _25365_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(net980),
    .S(_06592_),
    .X(_02507_));
 sg13g2_mux2_1 _25366_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(net979),
    .S(_06592_),
    .X(_02508_));
 sg13g2_mux2_1 _25367_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(net978),
    .S(_06592_),
    .X(_02509_));
 sg13g2_mux2_1 _25368_ (.A0(\cpu.intr.r_timer_reload[8] ),
    .A1(_10008_),
    .S(_06592_),
    .X(_02510_));
 sg13g2_mux2_1 _25369_ (.A0(\cpu.intr.r_timer_reload[9] ),
    .A1(_10013_),
    .S(_06592_),
    .X(_02511_));
 sg13g2_inv_1 _25370_ (.Y(_06600_),
    .A(_09664_));
 sg13g2_nor4_2 _25371_ (.A(_11666_),
    .B(_11665_),
    .C(_09683_),
    .Y(_06601_),
    .D(_11664_));
 sg13g2_or2_1 _25372_ (.X(_06602_),
    .B(_09662_),
    .A(\cpu.qspi.r_state[1] ));
 sg13g2_buf_1 _25373_ (.A(_06602_),
    .X(_06603_));
 sg13g2_nor3_1 _25374_ (.A(_11681_),
    .B(_11667_),
    .C(_11680_),
    .Y(_06604_));
 sg13g2_nor2b_1 _25375_ (.A(_06603_),
    .B_N(_06604_),
    .Y(_06605_));
 sg13g2_and4_1 _25376_ (.A(_09661_),
    .B(_11662_),
    .C(_06601_),
    .D(_06605_),
    .X(_06606_));
 sg13g2_buf_1 _25377_ (.A(_06606_),
    .X(_06607_));
 sg13g2_inv_1 _25378_ (.Y(_06608_),
    .A(_09738_));
 sg13g2_nor2_1 _25379_ (.A(net324),
    .B(net69),
    .Y(_06609_));
 sg13g2_and2_1 _25380_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(net69),
    .X(_06610_));
 sg13g2_a221oi_1 _25381_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06610_),
    .B1(_06609_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06611_),
    .A2(net324));
 sg13g2_nor2_1 _25382_ (.A(_09671_),
    .B(_09686_),
    .Y(_06612_));
 sg13g2_nor2_1 _25383_ (.A(_09682_),
    .B(_09673_),
    .Y(_06613_));
 sg13g2_nand2_2 _25384_ (.Y(_06614_),
    .A(_06612_),
    .B(_06613_));
 sg13g2_a221oi_1 _25385_ (.B2(_06614_),
    .C1(_09677_),
    .B1(_00183_),
    .A1(net1101),
    .Y(_06615_),
    .A2(_06600_));
 sg13g2_o21ai_1 _25386_ (.B1(_06615_),
    .Y(_06616_),
    .A1(_06608_),
    .A2(_06611_));
 sg13g2_nand2_1 _25387_ (.Y(_06617_),
    .A(net27),
    .B(_06616_));
 sg13g2_o21ai_1 _25388_ (.B1(_06617_),
    .Y(_02512_),
    .A1(_06600_),
    .A2(net27));
 sg13g2_or3_1 _25389_ (.A(_06608_),
    .B(net1101),
    .C(_06614_),
    .X(_06618_));
 sg13g2_xor2_1 _25390_ (.B(_09665_),
    .A(_09664_),
    .X(_06619_));
 sg13g2_o21ai_1 _25391_ (.B1(_06619_),
    .Y(_06620_),
    .A1(net1101),
    .A2(_06614_));
 sg13g2_inv_1 _25392_ (.Y(_06621_),
    .A(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_a22oi_1 _25393_ (.Y(_06622_),
    .B1(net69),
    .B2(\cpu.qspi.r_read_delay[1][1] ),
    .A2(net324),
    .A1(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_o21ai_1 _25394_ (.B1(_06622_),
    .Y(_06623_),
    .A1(_06621_),
    .A2(_09700_));
 sg13g2_a221oi_1 _25395_ (.B2(_09738_),
    .C1(_09677_),
    .B1(_06623_),
    .A1(_06618_),
    .Y(_06624_),
    .A2(_06620_));
 sg13g2_nor2_1 _25396_ (.A(_09665_),
    .B(net27),
    .Y(_06625_));
 sg13g2_a21oi_1 _25397_ (.A1(net27),
    .A2(_06624_),
    .Y(_02513_),
    .B1(_06625_));
 sg13g2_inv_1 _25398_ (.Y(_06626_),
    .A(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_a22oi_1 _25399_ (.Y(_06627_),
    .B1(_09698_),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(_09694_),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_o21ai_1 _25400_ (.B1(_06627_),
    .Y(_06628_),
    .A1(_06626_),
    .A2(_09700_));
 sg13g2_nor2_1 _25401_ (.A(_09664_),
    .B(_09665_),
    .Y(_06629_));
 sg13g2_xor2_1 _25402_ (.B(_06629_),
    .A(_00184_),
    .X(_06630_));
 sg13g2_mux2_1 _25403_ (.A0(_06614_),
    .A1(net671),
    .S(net1101),
    .X(_06631_));
 sg13g2_nand2_1 _25404_ (.Y(_06632_),
    .A(_06630_),
    .B(_06631_));
 sg13g2_a221oi_1 _25405_ (.B2(_06618_),
    .C1(_09677_),
    .B1(_06632_),
    .A1(_09738_),
    .Y(_06633_),
    .A2(_06628_));
 sg13g2_nor2_1 _25406_ (.A(_09666_),
    .B(net27),
    .Y(_06634_));
 sg13g2_a21oi_1 _25407_ (.A1(net27),
    .A2(_06633_),
    .Y(_02514_),
    .B1(_06634_));
 sg13g2_a21oi_1 _25408_ (.A1(net1101),
    .A2(net671),
    .Y(_06635_),
    .B1(_06614_));
 sg13g2_o21ai_1 _25409_ (.B1(net27),
    .Y(_06636_),
    .A1(_09667_),
    .A2(_06635_));
 sg13g2_inv_1 _25410_ (.Y(_06637_),
    .A(_06635_));
 sg13g2_inv_1 _25411_ (.Y(_06638_),
    .A(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_a22oi_1 _25412_ (.Y(_06639_),
    .B1(net69),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(net324),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_o21ai_1 _25413_ (.B1(_06639_),
    .Y(_06640_),
    .A1(_06638_),
    .A2(_09700_));
 sg13g2_a22oi_1 _25414_ (.Y(_06641_),
    .B1(_06640_),
    .B2(_09738_),
    .A2(_06637_),
    .A1(_09668_));
 sg13g2_nor2b_1 _25415_ (.A(_06641_),
    .B_N(_06607_),
    .Y(_06642_));
 sg13g2_a21o_1 _25416_ (.A2(_06636_),
    .A1(\cpu.qspi.r_count[3] ),
    .B1(_06642_),
    .X(_02515_));
 sg13g2_or2_1 _25417_ (.X(_06643_),
    .B(_09668_),
    .A(_00252_));
 sg13g2_a21oi_1 _25418_ (.A1(net671),
    .A2(_06643_),
    .Y(_06644_),
    .B1(_06635_));
 sg13g2_mux2_1 _25419_ (.A0(\cpu.qspi.r_count[4] ),
    .A1(_06644_),
    .S(net27),
    .X(_02516_));
 sg13g2_nand2_1 _25420_ (.Y(_06645_),
    .A(_09819_),
    .B(_06234_));
 sg13g2_buf_1 _25421_ (.A(_06645_),
    .X(_06646_));
 sg13g2_nor3_1 _25422_ (.A(net609),
    .B(net551),
    .C(net95),
    .Y(_06647_));
 sg13g2_buf_1 _25423_ (.A(_06647_),
    .X(_06648_));
 sg13g2_nand2_1 _25424_ (.Y(_06649_),
    .A(net959),
    .B(_06648_));
 sg13g2_nand3_1 _25425_ (.B(_09819_),
    .C(_06234_),
    .A(_09120_),
    .Y(_06650_));
 sg13g2_buf_1 _25426_ (.A(_06650_),
    .X(_06651_));
 sg13g2_nand2_1 _25427_ (.Y(_06652_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06651_));
 sg13g2_a21oi_1 _25428_ (.A1(_06649_),
    .A2(_06652_),
    .Y(_02527_),
    .B1(net610));
 sg13g2_nand2_1 _25429_ (.Y(_06653_),
    .A(net954),
    .B(_06648_));
 sg13g2_nand2_1 _25430_ (.Y(_06654_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06651_));
 sg13g2_a21oi_1 _25431_ (.A1(_06653_),
    .A2(_06654_),
    .Y(_02528_),
    .B1(net610));
 sg13g2_buf_1 _25432_ (.A(_09128_),
    .X(_06655_));
 sg13g2_nand2_1 _25433_ (.Y(_06656_),
    .A(_02848_),
    .B(_06648_));
 sg13g2_nand2_1 _25434_ (.Y(_06657_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06651_));
 sg13g2_nand3_1 _25435_ (.B(_06656_),
    .C(_06657_),
    .A(net629),
    .Y(_02529_));
 sg13g2_nand2_1 _25436_ (.Y(_06658_),
    .A(net1017),
    .B(_06648_));
 sg13g2_nand2_1 _25437_ (.Y(_06659_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06651_));
 sg13g2_a21oi_1 _25438_ (.A1(_06658_),
    .A2(_06659_),
    .Y(_02530_),
    .B1(net610));
 sg13g2_nor2_1 _25439_ (.A(_09959_),
    .B(net95),
    .Y(_06660_));
 sg13g2_nand2_1 _25440_ (.Y(_06661_),
    .A(net959),
    .B(_06660_));
 sg13g2_or2_1 _25441_ (.X(_06662_),
    .B(net95),
    .A(_09959_));
 sg13g2_buf_1 _25442_ (.A(_06662_),
    .X(_06663_));
 sg13g2_nand2_1 _25443_ (.Y(_06664_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06663_));
 sg13g2_a21oi_1 _25444_ (.A1(_06661_),
    .A2(_06664_),
    .Y(_02531_),
    .B1(net610));
 sg13g2_nand2_1 _25445_ (.Y(_06665_),
    .A(_02808_),
    .B(_06660_));
 sg13g2_nand2_1 _25446_ (.Y(_06666_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06663_));
 sg13g2_a21oi_1 _25447_ (.A1(_06665_),
    .A2(_06666_),
    .Y(_02532_),
    .B1(net610));
 sg13g2_nand2_1 _25448_ (.Y(_06667_),
    .A(_02848_),
    .B(_06660_));
 sg13g2_nand2_1 _25449_ (.Y(_06668_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06663_));
 sg13g2_nand3_1 _25450_ (.B(_06667_),
    .C(_06668_),
    .A(net629),
    .Y(_02533_));
 sg13g2_nand2_1 _25451_ (.Y(_06669_),
    .A(_09916_),
    .B(_06660_));
 sg13g2_nand2_1 _25452_ (.Y(_06670_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06663_));
 sg13g2_a21oi_1 _25453_ (.A1(_06669_),
    .A2(_06670_),
    .Y(_02534_),
    .B1(net610));
 sg13g2_nor2_1 _25454_ (.A(_04867_),
    .B(net95),
    .Y(_06671_));
 sg13g2_buf_1 _25455_ (.A(_06671_),
    .X(_06672_));
 sg13g2_nand2_1 _25456_ (.Y(_06673_),
    .A(net959),
    .B(_06672_));
 sg13g2_or2_1 _25457_ (.X(_06674_),
    .B(net95),
    .A(_04867_));
 sg13g2_buf_1 _25458_ (.A(_06674_),
    .X(_06675_));
 sg13g2_nand2_1 _25459_ (.Y(_06676_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06675_));
 sg13g2_a21oi_1 _25460_ (.A1(_06673_),
    .A2(_06676_),
    .Y(_02535_),
    .B1(net610));
 sg13g2_nand2_1 _25461_ (.Y(_06677_),
    .A(net954),
    .B(_06672_));
 sg13g2_nand2_1 _25462_ (.Y(_06678_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06675_));
 sg13g2_a21oi_1 _25463_ (.A1(_06677_),
    .A2(_06678_),
    .Y(_02536_),
    .B1(net610));
 sg13g2_nand2_1 _25464_ (.Y(_06679_),
    .A(net855),
    .B(_06672_));
 sg13g2_nand2_1 _25465_ (.Y(_06680_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06675_));
 sg13g2_nand3_1 _25466_ (.B(_06679_),
    .C(_06680_),
    .A(net680),
    .Y(_02537_));
 sg13g2_nand2_1 _25467_ (.Y(_06681_),
    .A(_09916_),
    .B(_06672_));
 sg13g2_nand2_1 _25468_ (.Y(_06682_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06675_));
 sg13g2_a21oi_1 _25469_ (.A1(_06681_),
    .A2(_06682_),
    .Y(_02538_),
    .B1(_09710_));
 sg13g2_buf_1 _25470_ (.A(_08830_),
    .X(_06683_));
 sg13g2_buf_1 _25471_ (.A(_06683_),
    .X(_06684_));
 sg13g2_buf_1 _25472_ (.A(_08830_),
    .X(_06685_));
 sg13g2_buf_1 _25473_ (.A(_09655_),
    .X(_06686_));
 sg13g2_mux2_1 _25474_ (.A0(net344),
    .A1(_09297_),
    .S(net94),
    .X(_06687_));
 sg13g2_nand2_1 _25475_ (.Y(_06688_),
    .A(net696),
    .B(_06687_));
 sg13g2_o21ai_1 _25476_ (.B1(_06688_),
    .Y(_06689_),
    .A1(net628),
    .A2(_08401_));
 sg13g2_nand2_1 _25477_ (.Y(_06690_),
    .A(_09378_),
    .B(net94));
 sg13g2_o21ai_1 _25478_ (.B1(_06690_),
    .Y(_06691_),
    .A1(_00235_),
    .A2(net94));
 sg13g2_nand2_1 _25479_ (.Y(_06692_),
    .A(net696),
    .B(_06691_));
 sg13g2_o21ai_1 _25480_ (.B1(_06692_),
    .Y(_06693_),
    .A1(net628),
    .A2(_10695_));
 sg13g2_mux2_1 _25481_ (.A0(net435),
    .A1(_09522_),
    .S(_09655_),
    .X(_06694_));
 sg13g2_nand2_1 _25482_ (.Y(_06695_),
    .A(net697),
    .B(_06694_));
 sg13g2_o21ai_1 _25483_ (.B1(_06695_),
    .Y(_06696_),
    .A1(net697),
    .A2(_08498_));
 sg13g2_nand2_1 _25484_ (.Y(_06697_),
    .A(_09683_),
    .B(net107));
 sg13g2_nand2b_1 _25485_ (.Y(_06698_),
    .B(_11771_),
    .A_N(_11770_));
 sg13g2_a22oi_1 _25486_ (.Y(_06699_),
    .B1(_05169_),
    .B2(_11821_),
    .A2(_04838_),
    .A1(net863));
 sg13g2_o21ai_1 _25487_ (.B1(_06699_),
    .Y(_06700_),
    .A1(_06698_),
    .A2(_04816_));
 sg13g2_nand2b_1 _25488_ (.Y(_06701_),
    .B(net992),
    .A_N(_11771_));
 sg13g2_nand2_1 _25489_ (.Y(_06702_),
    .A(_11772_),
    .B(_04809_));
 sg13g2_o21ai_1 _25490_ (.B1(_06702_),
    .Y(_06703_),
    .A1(_06701_),
    .A2(_05162_));
 sg13g2_nand3_1 _25491_ (.B(net863),
    .C(_04831_),
    .A(_11767_),
    .Y(_06704_));
 sg13g2_inv_1 _25492_ (.Y(_06705_),
    .A(_11767_));
 sg13g2_nor2_1 _25493_ (.A(_06705_),
    .B(_11860_),
    .Y(_06706_));
 sg13g2_nor2_2 _25494_ (.A(net1080),
    .B(_06706_),
    .Y(_06707_));
 sg13g2_a21oi_1 _25495_ (.A1(_11860_),
    .A2(_05542_),
    .Y(_06708_),
    .B1(_06707_));
 sg13g2_nand2_1 _25496_ (.Y(_06709_),
    .A(_06704_),
    .B(_06708_));
 sg13g2_a221oi_1 _25497_ (.B2(_11768_),
    .C1(_06709_),
    .B1(_06703_),
    .A1(net1080),
    .Y(_06710_),
    .A2(_06700_));
 sg13g2_nand2_1 _25498_ (.Y(_06711_),
    .A(_05533_),
    .B(_06707_));
 sg13g2_nand3b_1 _25499_ (.B(_06711_),
    .C(_09673_),
    .Y(_06712_),
    .A_N(_06710_));
 sg13g2_nand2_1 _25500_ (.Y(_06713_),
    .A(_06604_),
    .B(_06613_));
 sg13g2_nor2_1 _25501_ (.A(_09677_),
    .B(_06713_),
    .Y(_06714_));
 sg13g2_nor2b_1 _25502_ (.A(net1102),
    .B_N(_06601_),
    .Y(_06715_));
 sg13g2_and3_1 _25503_ (.X(_06716_),
    .A(_09685_),
    .B(_06714_),
    .C(_06715_));
 sg13g2_buf_1 _25504_ (.A(_06716_),
    .X(_06717_));
 sg13g2_nor2_1 _25505_ (.A(_11666_),
    .B(_06717_),
    .Y(_06718_));
 sg13g2_buf_1 _25506_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06719_));
 sg13g2_buf_1 _25507_ (.A(_08734_),
    .X(_06720_));
 sg13g2_nand2_1 _25508_ (.Y(_06721_),
    .A(net1116),
    .B(_08734_));
 sg13g2_o21ai_1 _25509_ (.B1(_06721_),
    .Y(_06722_),
    .A1(net927),
    .A2(_03702_));
 sg13g2_a22oi_1 _25510_ (.Y(_06723_),
    .B1(_06722_),
    .B2(_11680_),
    .A2(_06719_),
    .A1(_09711_));
 sg13g2_nand4_1 _25511_ (.B(_06712_),
    .C(_06718_),
    .A(_06697_),
    .Y(_06724_),
    .D(_06723_));
 sg13g2_a21o_1 _25512_ (.A2(_06696_),
    .A1(_11681_),
    .B1(_06724_),
    .X(_06725_));
 sg13g2_a221oi_1 _25513_ (.B2(_11665_),
    .C1(_06725_),
    .B1(_06693_),
    .A1(_11667_),
    .Y(_06726_),
    .A2(_06689_));
 sg13g2_nand2_1 _25514_ (.Y(_06727_),
    .A(net1102),
    .B(_09663_));
 sg13g2_nand3b_1 _25515_ (.B(_00183_),
    .C(_06727_),
    .Y(_06728_),
    .A_N(_09665_));
 sg13g2_nor2_1 _25516_ (.A(net1102),
    .B(net107),
    .Y(_06729_));
 sg13g2_o21ai_1 _25517_ (.B1(_09666_),
    .Y(_06730_),
    .A1(_06728_),
    .A2(_06729_));
 sg13g2_nand3_1 _25518_ (.B(_09665_),
    .C(_06727_),
    .A(_06600_),
    .Y(_06731_));
 sg13g2_o21ai_1 _25519_ (.B1(_06731_),
    .Y(_06732_),
    .A1(_06600_),
    .A2(_06727_));
 sg13g2_nor2_1 _25520_ (.A(_09666_),
    .B(_06732_),
    .Y(_06733_));
 sg13g2_o21ai_1 _25521_ (.B1(_06733_),
    .Y(_06734_),
    .A1(net1102),
    .A2(_09665_));
 sg13g2_o21ai_1 _25522_ (.B1(_06734_),
    .Y(_06735_),
    .A1(_09665_),
    .A2(_06730_));
 sg13g2_nor3_1 _25523_ (.A(net1102),
    .B(_09664_),
    .C(_06730_),
    .Y(_06736_));
 sg13g2_o21ai_1 _25524_ (.B1(net107),
    .Y(_06737_),
    .A1(_06733_),
    .A2(_06736_));
 sg13g2_nand2b_1 _25525_ (.Y(_06738_),
    .B(_06737_),
    .A_N(_06735_));
 sg13g2_o21ai_1 _25526_ (.B1(_06738_),
    .Y(_06739_),
    .A1(_09682_),
    .A2(net1102));
 sg13g2_xnor2_1 _25527_ (.Y(_06740_),
    .A(net107),
    .B(_09703_));
 sg13g2_a22oi_1 _25528_ (.Y(_06741_),
    .B1(_06740_),
    .B2(_06717_),
    .A2(_06739_),
    .A1(_06726_));
 sg13g2_and2_1 _25529_ (.A(\cpu.qspi.r_mask[1] ),
    .B(net69),
    .X(_06742_));
 sg13g2_a221oi_1 _25530_ (.B2(\cpu.qspi.r_mask[0] ),
    .C1(_06742_),
    .B1(_06609_),
    .A1(\cpu.qspi.r_mask[2] ),
    .Y(_06743_),
    .A2(net324));
 sg13g2_nor2_1 _25531_ (.A(_09671_),
    .B(_06603_),
    .Y(_06744_));
 sg13g2_nor2_1 _25532_ (.A(_09738_),
    .B(net1101),
    .Y(_06745_));
 sg13g2_nand3_1 _25533_ (.B(_06744_),
    .C(_06745_),
    .A(_09661_),
    .Y(_06746_));
 sg13g2_a21oi_1 _25534_ (.A1(_11666_),
    .A2(_06743_),
    .Y(_06747_),
    .B1(_06746_));
 sg13g2_buf_2 _25535_ (.A(_06747_),
    .X(_06748_));
 sg13g2_mux2_1 _25536_ (.A0(net11),
    .A1(_06741_),
    .S(_06748_),
    .X(_02543_));
 sg13g2_nand2_1 _25537_ (.Y(_06749_),
    .A(net927),
    .B(_10399_));
 sg13g2_nand2_1 _25538_ (.Y(_06750_),
    .A(_09400_),
    .B(_06686_));
 sg13g2_o21ai_1 _25539_ (.B1(_06750_),
    .Y(_06751_),
    .A1(_04932_),
    .A2(net94));
 sg13g2_nand2b_1 _25540_ (.Y(_06752_),
    .B(net628),
    .A_N(_06751_));
 sg13g2_nand3_1 _25541_ (.B(_06749_),
    .C(_06752_),
    .A(_11680_),
    .Y(_06753_));
 sg13g2_mux2_1 _25542_ (.A0(net376),
    .A1(_09323_),
    .S(_09655_),
    .X(_06754_));
 sg13g2_nand2_1 _25543_ (.Y(_06755_),
    .A(net697),
    .B(_06754_));
 sg13g2_o21ai_1 _25544_ (.B1(_06755_),
    .Y(_06756_),
    .A1(net696),
    .A2(_08426_));
 sg13g2_buf_1 _25545_ (.A(_09655_),
    .X(_06757_));
 sg13g2_mux2_1 _25546_ (.A0(_09586_),
    .A1(_09593_),
    .S(net93),
    .X(_06758_));
 sg13g2_nand2_1 _25547_ (.Y(_06759_),
    .A(net697),
    .B(_06758_));
 sg13g2_o21ai_1 _25548_ (.B1(_06759_),
    .Y(_06760_),
    .A1(net696),
    .A2(_08543_));
 sg13g2_a22oi_1 _25549_ (.Y(_06761_),
    .B1(_06760_),
    .B2(_11681_),
    .A2(_06756_),
    .A1(_11667_));
 sg13g2_mux2_1 _25550_ (.A0(_05264_),
    .A1(_05288_),
    .S(net992),
    .X(_06762_));
 sg13g2_buf_1 _25551_ (.A(_11771_),
    .X(_06763_));
 sg13g2_nand3b_1 _25552_ (.B(net993),
    .C(net926),
    .Y(_06764_),
    .A_N(_06762_));
 sg13g2_mux2_1 _25553_ (.A0(_05607_),
    .A1(_05271_),
    .S(net926),
    .X(_06765_));
 sg13g2_nor2b_1 _25554_ (.A(net992),
    .B_N(net1080),
    .Y(_06766_));
 sg13g2_nand2b_1 _25555_ (.Y(_06767_),
    .B(_06766_),
    .A_N(_06765_));
 sg13g2_nor3_1 _25556_ (.A(_06705_),
    .B(_06701_),
    .C(_05193_),
    .Y(_06768_));
 sg13g2_a21oi_1 _25557_ (.A1(_05599_),
    .A2(_06707_),
    .Y(_06769_),
    .B1(_06768_));
 sg13g2_nand2_1 _25558_ (.Y(_06770_),
    .A(net926),
    .B(_05280_));
 sg13g2_o21ai_1 _25559_ (.B1(_06770_),
    .Y(_06771_),
    .A1(net926),
    .A2(_05201_));
 sg13g2_nand3_1 _25560_ (.B(net977),
    .C(_06771_),
    .A(net992),
    .Y(_06772_));
 sg13g2_nand4_1 _25561_ (.B(_06767_),
    .C(_06769_),
    .A(_06764_),
    .Y(_06773_),
    .D(_06772_));
 sg13g2_a221oi_1 _25562_ (.B2(_09673_),
    .C1(_11666_),
    .B1(_06773_),
    .A1(_09683_),
    .Y(_06774_),
    .A2(net107));
 sg13g2_mux2_1 _25563_ (.A0(_09357_),
    .A1(_09368_),
    .S(_06757_),
    .X(_06775_));
 sg13g2_nand2_1 _25564_ (.Y(_06776_),
    .A(net697),
    .B(_06775_));
 sg13g2_o21ai_1 _25565_ (.B1(_06776_),
    .Y(_06777_),
    .A1(net628),
    .A2(_10626_));
 sg13g2_nand2_1 _25566_ (.Y(_06778_),
    .A(_11665_),
    .B(_06777_));
 sg13g2_nand4_1 _25567_ (.B(_06761_),
    .C(_06774_),
    .A(_06753_),
    .Y(_06779_),
    .D(_06778_));
 sg13g2_a21oi_1 _25568_ (.A1(_09703_),
    .A2(_06717_),
    .Y(_06780_),
    .B1(_06779_));
 sg13g2_nor2_1 _25569_ (.A(net12),
    .B(_06748_),
    .Y(_06781_));
 sg13g2_a21oi_1 _25570_ (.A1(_06748_),
    .A2(_06780_),
    .Y(_02544_),
    .B1(_06781_));
 sg13g2_inv_1 _25571_ (.Y(_06782_),
    .A(net13));
 sg13g2_nand2_1 _25572_ (.Y(_06783_),
    .A(net977),
    .B(_05641_));
 sg13g2_a22oi_1 _25573_ (.Y(_06784_),
    .B1(_05349_),
    .B2(net993),
    .A2(_05356_),
    .A1(net977));
 sg13g2_a22oi_1 _25574_ (.Y(_06785_),
    .B1(_05233_),
    .B2(net977),
    .A2(_05225_),
    .A1(net993));
 sg13g2_nand2_1 _25575_ (.Y(_06786_),
    .A(net993),
    .B(_05090_));
 sg13g2_mux4_1 _25576_ (.S0(net926),
    .A0(_06783_),
    .A1(_06784_),
    .A2(_06785_),
    .A3(_06786_),
    .S1(net992),
    .X(_06787_));
 sg13g2_nand2b_1 _25577_ (.Y(_06788_),
    .B(_06707_),
    .A_N(_05632_));
 sg13g2_nand3_1 _25578_ (.B(net863),
    .C(_05097_),
    .A(net977),
    .Y(_06789_));
 sg13g2_nand3_1 _25579_ (.B(_06788_),
    .C(_06789_),
    .A(_06787_),
    .Y(_06790_));
 sg13g2_mux2_1 _25580_ (.A0(net796),
    .A1(net638),
    .S(_08830_),
    .X(_06791_));
 sg13g2_o21ai_1 _25581_ (.B1(_06718_),
    .Y(_06792_),
    .A1(_00185_),
    .A2(_06791_));
 sg13g2_a21oi_1 _25582_ (.A1(_09673_),
    .A2(_06790_),
    .Y(_06793_),
    .B1(_06792_));
 sg13g2_nand2_1 _25583_ (.Y(_06794_),
    .A(_09416_),
    .B(net93));
 sg13g2_o21ai_1 _25584_ (.B1(_06794_),
    .Y(_06795_),
    .A1(_00231_),
    .A2(net94));
 sg13g2_nand2_1 _25585_ (.Y(_06796_),
    .A(net697),
    .B(_06795_));
 sg13g2_o21ai_1 _25586_ (.B1(_06796_),
    .Y(_06797_),
    .A1(net696),
    .A2(_00295_));
 sg13g2_mux2_1 _25587_ (.A0(net436),
    .A1(_09500_),
    .S(net93),
    .X(_06798_));
 sg13g2_nand2_1 _25588_ (.Y(_06799_),
    .A(net696),
    .B(_06798_));
 sg13g2_o21ai_1 _25589_ (.B1(_06799_),
    .Y(_06800_),
    .A1(net628),
    .A2(_08607_));
 sg13g2_a22oi_1 _25590_ (.Y(_06801_),
    .B1(_06800_),
    .B2(_11667_),
    .A2(_06797_),
    .A1(_11680_));
 sg13g2_nand2_1 _25591_ (.Y(_06802_),
    .A(_09408_),
    .B(_06757_));
 sg13g2_o21ai_1 _25592_ (.B1(_06802_),
    .Y(_06803_),
    .A1(_00239_),
    .A2(net94));
 sg13g2_nand2_1 _25593_ (.Y(_06804_),
    .A(_06683_),
    .B(_06803_));
 sg13g2_o21ai_1 _25594_ (.B1(_06804_),
    .Y(_06805_),
    .A1(net696),
    .A2(_10651_));
 sg13g2_inv_1 _25595_ (.Y(_06806_),
    .A(_09355_));
 sg13g2_mux2_1 _25596_ (.A0(net439),
    .A1(_06806_),
    .S(net93),
    .X(_06807_));
 sg13g2_nand2_1 _25597_ (.Y(_06808_),
    .A(net696),
    .B(_06807_));
 sg13g2_o21ai_1 _25598_ (.B1(_06808_),
    .Y(_06809_),
    .A1(net628),
    .A2(_08564_));
 sg13g2_a22oi_1 _25599_ (.Y(_06810_),
    .B1(_06809_),
    .B2(_11681_),
    .A2(_06805_),
    .A1(_11665_));
 sg13g2_nand3_1 _25600_ (.B(_06801_),
    .C(_06810_),
    .A(_06793_),
    .Y(_06811_));
 sg13g2_o21ai_1 _25601_ (.B1(_06717_),
    .Y(_06812_),
    .A1(_09680_),
    .A2(_09704_));
 sg13g2_nand3_1 _25602_ (.B(_06811_),
    .C(_06812_),
    .A(_06748_),
    .Y(_06813_));
 sg13g2_o21ai_1 _25603_ (.B1(_06813_),
    .Y(_02545_),
    .A1(_06782_),
    .A2(_06748_));
 sg13g2_inv_1 _25604_ (.Y(_06814_),
    .A(net14));
 sg13g2_mux2_1 _25605_ (.A0(_00241_),
    .A1(_09425_),
    .S(_06686_),
    .X(_06815_));
 sg13g2_nand2b_1 _25606_ (.Y(_06816_),
    .B(net927),
    .A_N(_10676_));
 sg13g2_o21ai_1 _25607_ (.B1(_06816_),
    .Y(_06817_),
    .A1(net927),
    .A2(_06815_));
 sg13g2_nand2_1 _25608_ (.Y(_06818_),
    .A(_09474_),
    .B(net93));
 sg13g2_o21ai_1 _25609_ (.B1(_06818_),
    .Y(_06819_),
    .A1(_02912_),
    .A2(net94));
 sg13g2_nor2_1 _25610_ (.A(net927),
    .B(_06819_),
    .Y(_06820_));
 sg13g2_a21oi_1 _25611_ (.A1(net927),
    .A2(_08450_),
    .Y(_06821_),
    .B1(_06820_));
 sg13g2_nand2_1 _25612_ (.Y(_06822_),
    .A(_09689_),
    .B(_11664_));
 sg13g2_nor2_1 _25613_ (.A(_09690_),
    .B(_06822_),
    .Y(_06823_));
 sg13g2_a22oi_1 _25614_ (.Y(_06824_),
    .B1(_06821_),
    .B2(_06823_),
    .A2(_06817_),
    .A1(_11665_));
 sg13g2_mux2_1 _25615_ (.A0(net438),
    .A1(_09451_),
    .S(net93),
    .X(_06825_));
 sg13g2_nand2_1 _25616_ (.Y(_06826_),
    .A(net697),
    .B(_06825_));
 sg13g2_o21ai_1 _25617_ (.B1(_06826_),
    .Y(_06827_),
    .A1(net628),
    .A2(_08522_));
 sg13g2_nand2_1 _25618_ (.Y(_06828_),
    .A(_11771_),
    .B(_05140_));
 sg13g2_o21ai_1 _25619_ (.B1(_06828_),
    .Y(_06829_),
    .A1(_06763_),
    .A2(_05052_));
 sg13g2_nand3_1 _25620_ (.B(net977),
    .C(_06829_),
    .A(net992),
    .Y(_06830_));
 sg13g2_o21ai_1 _25621_ (.B1(_06830_),
    .Y(_06831_),
    .A1(net977),
    .A2(net993));
 sg13g2_or2_1 _25622_ (.X(_06832_),
    .B(net1080),
    .A(_06763_));
 sg13g2_nand3_1 _25623_ (.B(_11768_),
    .C(_05453_),
    .A(net926),
    .Y(_06833_));
 sg13g2_a21oi_1 _25624_ (.A1(_06832_),
    .A2(_06833_),
    .Y(_06834_),
    .B1(net992));
 sg13g2_and2_1 _25625_ (.A(net992),
    .B(_11767_),
    .X(_06835_));
 sg13g2_a22oi_1 _25626_ (.Y(_06836_),
    .B1(_06835_),
    .B2(_05133_),
    .A2(_06766_),
    .A1(_05460_));
 sg13g2_a221oi_1 _25627_ (.B2(_05041_),
    .C1(net926),
    .B1(_06835_),
    .A1(_05072_),
    .Y(_06837_),
    .A2(_06766_));
 sg13g2_a21oi_1 _25628_ (.A1(net926),
    .A2(_06836_),
    .Y(_06838_),
    .B1(_06837_));
 sg13g2_nor3_1 _25629_ (.A(_06831_),
    .B(_06834_),
    .C(_06838_),
    .Y(_06839_));
 sg13g2_nand2b_1 _25630_ (.Y(_06840_),
    .B(_06707_),
    .A_N(_05061_));
 sg13g2_nand2_1 _25631_ (.Y(_06841_),
    .A(_09673_),
    .B(_06840_));
 sg13g2_nand2_1 _25632_ (.Y(_06842_),
    .A(net690),
    .B(net927));
 sg13g2_nand2_1 _25633_ (.Y(_06843_),
    .A(_08830_),
    .B(net496));
 sg13g2_a21oi_1 _25634_ (.A1(_06842_),
    .A2(_06843_),
    .Y(_06844_),
    .B1(_00185_));
 sg13g2_nor4_1 _25635_ (.A(_11666_),
    .B(_09683_),
    .C(_06717_),
    .D(_06844_),
    .Y(_06845_));
 sg13g2_o21ai_1 _25636_ (.B1(_06845_),
    .Y(_06846_),
    .A1(_06839_),
    .A2(_06841_));
 sg13g2_a21oi_1 _25637_ (.A1(_11667_),
    .A2(_06827_),
    .Y(_06847_),
    .B1(_06846_));
 sg13g2_inv_1 _25638_ (.Y(_06848_),
    .A(_09570_));
 sg13g2_mux2_1 _25639_ (.A0(_09562_),
    .A1(_06848_),
    .S(net93),
    .X(_06849_));
 sg13g2_nand2_1 _25640_ (.Y(_06850_),
    .A(net697),
    .B(_06849_));
 sg13g2_o21ai_1 _25641_ (.B1(_06850_),
    .Y(_06851_),
    .A1(_06685_),
    .A2(_08650_));
 sg13g2_nand2_1 _25642_ (.Y(_06852_),
    .A(_09386_),
    .B(net93));
 sg13g2_o21ai_1 _25643_ (.B1(_06852_),
    .Y(_06853_),
    .A1(_00233_),
    .A2(net94));
 sg13g2_nand2_1 _25644_ (.Y(_06854_),
    .A(_06685_),
    .B(_06853_));
 sg13g2_o21ai_1 _25645_ (.B1(_06854_),
    .Y(_06855_),
    .A1(net628),
    .A2(_10398_));
 sg13g2_a22oi_1 _25646_ (.Y(_06856_),
    .B1(_06855_),
    .B2(_11680_),
    .A2(_06851_),
    .A1(_11681_));
 sg13g2_nand3_1 _25647_ (.B(_06847_),
    .C(_06856_),
    .A(_06824_),
    .Y(_06857_));
 sg13g2_nand3_1 _25648_ (.B(_06812_),
    .C(_06857_),
    .A(_06748_),
    .Y(_06858_));
 sg13g2_o21ai_1 _25649_ (.B1(_06858_),
    .Y(_02546_),
    .A1(_06814_),
    .A2(_06748_));
 sg13g2_nor2_1 _25650_ (.A(_09111_),
    .B(net310),
    .Y(_06859_));
 sg13g2_buf_4 _25651_ (.X(_06860_),
    .A(_06859_));
 sg13g2_mux2_1 _25652_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(net861),
    .S(_06860_),
    .X(_02551_));
 sg13g2_mux2_1 _25653_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(net859),
    .S(_06860_),
    .X(_02552_));
 sg13g2_mux2_1 _25654_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(net858),
    .S(_06860_),
    .X(_02553_));
 sg13g2_mux2_1 _25655_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(net982),
    .S(_06860_),
    .X(_02554_));
 sg13g2_mux2_1 _25656_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(net981),
    .S(_06860_),
    .X(_02555_));
 sg13g2_mux2_1 _25657_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(net980),
    .S(_06860_),
    .X(_02556_));
 sg13g2_mux2_1 _25658_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(net979),
    .S(_06860_),
    .X(_02557_));
 sg13g2_mux2_1 _25659_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(net978),
    .S(_06860_),
    .X(_02558_));
 sg13g2_nor4_1 _25660_ (.A(net731),
    .B(net667),
    .C(_09111_),
    .D(net480),
    .Y(_06861_));
 sg13g2_buf_4 _25661_ (.X(_06862_),
    .A(_06861_));
 sg13g2_mux2_1 _25662_ (.A0(\cpu.spi.r_clk_count[1][0] ),
    .A1(net861),
    .S(_06862_),
    .X(_02559_));
 sg13g2_mux2_1 _25663_ (.A0(\cpu.spi.r_clk_count[1][1] ),
    .A1(net859),
    .S(_06862_),
    .X(_02560_));
 sg13g2_mux2_1 _25664_ (.A0(\cpu.spi.r_clk_count[1][2] ),
    .A1(net858),
    .S(_06862_),
    .X(_02561_));
 sg13g2_mux2_1 _25665_ (.A0(\cpu.spi.r_clk_count[1][3] ),
    .A1(net982),
    .S(_06862_),
    .X(_02562_));
 sg13g2_mux2_1 _25666_ (.A0(\cpu.spi.r_clk_count[1][4] ),
    .A1(net981),
    .S(_06862_),
    .X(_02563_));
 sg13g2_mux2_1 _25667_ (.A0(\cpu.spi.r_clk_count[1][5] ),
    .A1(net980),
    .S(_06862_),
    .X(_02564_));
 sg13g2_mux2_1 _25668_ (.A0(\cpu.spi.r_clk_count[1][6] ),
    .A1(net979),
    .S(_06862_),
    .X(_02565_));
 sg13g2_mux2_1 _25669_ (.A0(\cpu.spi.r_clk_count[1][7] ),
    .A1(net978),
    .S(_06862_),
    .X(_02566_));
 sg13g2_and4_1 _25670_ (.A(net609),
    .B(_09133_),
    .C(net894),
    .D(_11721_),
    .X(_06863_));
 sg13g2_buf_4 _25671_ (.X(_06864_),
    .A(_06863_));
 sg13g2_mux2_1 _25672_ (.A0(_04969_),
    .A1(net861),
    .S(_06864_),
    .X(_02567_));
 sg13g2_mux2_1 _25673_ (.A0(_05306_),
    .A1(net859),
    .S(_06864_),
    .X(_02568_));
 sg13g2_mux2_1 _25674_ (.A0(_05364_),
    .A1(net858),
    .S(_06864_),
    .X(_02569_));
 sg13g2_mux2_1 _25675_ (.A0(_05415_),
    .A1(net982),
    .S(_06864_),
    .X(_02570_));
 sg13g2_mux2_1 _25676_ (.A0(_05516_),
    .A1(net981),
    .S(_06864_),
    .X(_02571_));
 sg13g2_mux2_1 _25677_ (.A0(_05557_),
    .A1(net980),
    .S(_06864_),
    .X(_02572_));
 sg13g2_mux2_1 _25678_ (.A0(_05647_),
    .A1(net979),
    .S(_06864_),
    .X(_02573_));
 sg13g2_mux2_1 _25679_ (.A0(_05012_),
    .A1(net978),
    .S(_06864_),
    .X(_02574_));
 sg13g2_o21ai_1 _25680_ (.B1(_09114_),
    .Y(_06865_),
    .A1(net377),
    .A2(_09104_));
 sg13g2_buf_1 _25681_ (.A(_00225_),
    .X(_06866_));
 sg13g2_inv_1 _25682_ (.Y(_06867_),
    .A(_09116_));
 sg13g2_nor4_1 _25683_ (.A(\cpu.spi.r_state[3] ),
    .B(\cpu.spi.r_state[5] ),
    .C(net1104),
    .D(_11683_),
    .Y(_06868_));
 sg13g2_buf_1 _25684_ (.A(_06868_),
    .X(_06869_));
 sg13g2_and2_1 _25685_ (.A(_06867_),
    .B(_06869_),
    .X(_06870_));
 sg13g2_nor2_1 _25686_ (.A(_06866_),
    .B(net377),
    .Y(_06871_));
 sg13g2_a22oi_1 _25687_ (.Y(_06872_),
    .B1(_06871_),
    .B2(net80),
    .A2(_06870_),
    .A1(_06866_));
 sg13g2_nand3_1 _25688_ (.B(_06865_),
    .C(_06872_),
    .A(_09124_),
    .Y(_06873_));
 sg13g2_buf_2 _25689_ (.A(_06873_),
    .X(_06874_));
 sg13g2_buf_1 _25690_ (.A(_06874_),
    .X(_06875_));
 sg13g2_buf_1 _25691_ (.A(net489),
    .X(_06876_));
 sg13g2_nand2b_1 _25692_ (.Y(_06877_),
    .B(net424),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _25693_ (.B1(_06877_),
    .Y(_06878_),
    .A1(net389),
    .A2(_04969_));
 sg13g2_mux2_1 _25694_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net424),
    .X(_06879_));
 sg13g2_nor2_1 _25695_ (.A(net731),
    .B(_06879_),
    .Y(_06880_));
 sg13g2_a21oi_1 _25696_ (.A1(net644),
    .A2(_06878_),
    .Y(_06881_),
    .B1(_06880_));
 sg13g2_nand2_1 _25697_ (.Y(_06882_),
    .A(_06866_),
    .B(net627));
 sg13g2_buf_1 _25698_ (.A(_06882_),
    .X(_06883_));
 sg13g2_buf_1 _25699_ (.A(_06883_),
    .X(_06884_));
 sg13g2_nor2_1 _25700_ (.A(net996),
    .B(_04969_),
    .Y(_06885_));
 sg13g2_a21oi_1 _25701_ (.A1(net998),
    .A2(_00314_),
    .Y(_06886_),
    .B1(_06885_));
 sg13g2_mux2_1 _25702_ (.A0(_00314_),
    .A1(_00313_),
    .S(_11693_),
    .X(_06887_));
 sg13g2_nor2_1 _25703_ (.A(net997),
    .B(_06887_),
    .Y(_06888_));
 sg13g2_a21oi_1 _25704_ (.A1(net999),
    .A2(_06886_),
    .Y(_06889_),
    .B1(_06888_));
 sg13g2_nand2_1 _25705_ (.Y(_06890_),
    .A(net345),
    .B(_06889_));
 sg13g2_nor2_1 _25706_ (.A(_09001_),
    .B(_06869_),
    .Y(_06891_));
 sg13g2_and2_1 _25707_ (.A(_09191_),
    .B(_06889_),
    .X(_06892_));
 sg13g2_a21oi_1 _25708_ (.A1(_09001_),
    .A2(_09134_),
    .Y(_06893_),
    .B1(_06892_));
 sg13g2_buf_1 _25709_ (.A(_09105_),
    .X(_06894_));
 sg13g2_a22oi_1 _25710_ (.Y(_06895_),
    .B1(_06893_),
    .B2(_06894_),
    .A2(_06891_),
    .A1(_06890_));
 sg13g2_nand2_1 _25711_ (.Y(_06896_),
    .A(net453),
    .B(_06895_));
 sg13g2_o21ai_1 _25712_ (.B1(_06896_),
    .Y(_06897_),
    .A1(_06881_),
    .A2(net453));
 sg13g2_nand2_1 _25713_ (.Y(_06898_),
    .A(_09001_),
    .B(net30));
 sg13g2_o21ai_1 _25714_ (.B1(_06898_),
    .Y(_02575_),
    .A1(_06875_),
    .A2(_06897_));
 sg13g2_nand2b_1 _25715_ (.Y(_06899_),
    .B(net389),
    .A_N(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_o21ai_1 _25716_ (.B1(_06899_),
    .Y(_06900_),
    .A1(net366),
    .A2(_05306_));
 sg13g2_mux2_1 _25717_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(_11728_),
    .X(_06901_));
 sg13g2_nor2_1 _25718_ (.A(_11727_),
    .B(_06901_),
    .Y(_06902_));
 sg13g2_a21oi_1 _25719_ (.A1(net643),
    .A2(_06900_),
    .Y(_06903_),
    .B1(_06902_));
 sg13g2_nor2_1 _25720_ (.A(net998),
    .B(_05306_),
    .Y(_06904_));
 sg13g2_a21oi_1 _25721_ (.A1(net867),
    .A2(_00095_),
    .Y(_06905_),
    .B1(_06904_));
 sg13g2_mux2_1 _25722_ (.A0(_00095_),
    .A1(_00094_),
    .S(_11697_),
    .X(_06906_));
 sg13g2_nor2_1 _25723_ (.A(net997),
    .B(_06906_),
    .Y(_06907_));
 sg13g2_a21oi_1 _25724_ (.A1(net999),
    .A2(_06905_),
    .Y(_06908_),
    .B1(_06907_));
 sg13g2_nand2_1 _25725_ (.Y(_06909_),
    .A(net345),
    .B(_06908_));
 sg13g2_xor2_1 _25726_ (.B(\cpu.spi.r_count[1] ),
    .A(_09001_),
    .X(_06910_));
 sg13g2_nor2_1 _25727_ (.A(net627),
    .B(_06910_),
    .Y(_06911_));
 sg13g2_nand2b_1 _25728_ (.Y(_06912_),
    .B(net80),
    .A_N(_06908_));
 sg13g2_o21ai_1 _25729_ (.B1(_06912_),
    .Y(_06913_),
    .A1(net70),
    .A2(_06910_));
 sg13g2_a22oi_1 _25730_ (.Y(_06914_),
    .B1(_06913_),
    .B2(net925),
    .A2(_06911_),
    .A1(_06909_));
 sg13g2_nand2_1 _25731_ (.Y(_06915_),
    .A(net453),
    .B(_06914_));
 sg13g2_o21ai_1 _25732_ (.B1(_06915_),
    .Y(_06916_),
    .A1(net453),
    .A2(_06903_));
 sg13g2_nand2_1 _25733_ (.Y(_06917_),
    .A(\cpu.spi.r_count[1] ),
    .B(net30));
 sg13g2_o21ai_1 _25734_ (.B1(_06917_),
    .Y(_02576_),
    .A1(net30),
    .A2(_06916_));
 sg13g2_nand2b_1 _25735_ (.Y(_06918_),
    .B(net389),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _25736_ (.B1(_06918_),
    .Y(_06919_),
    .A1(net366),
    .A2(_05364_));
 sg13g2_mux2_1 _25737_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net424),
    .X(_06920_));
 sg13g2_nor2_1 _25738_ (.A(net644),
    .B(_06920_),
    .Y(_06921_));
 sg13g2_a21oi_1 _25739_ (.A1(net644),
    .A2(_06919_),
    .Y(_06922_),
    .B1(_06921_));
 sg13g2_nor2_1 _25740_ (.A(net998),
    .B(_05364_),
    .Y(_06923_));
 sg13g2_a21oi_1 _25741_ (.A1(net867),
    .A2(_00105_),
    .Y(_06924_),
    .B1(_06923_));
 sg13g2_mux2_1 _25742_ (.A0(_00105_),
    .A1(_00104_),
    .S(net996),
    .X(_06925_));
 sg13g2_nor2_1 _25743_ (.A(net997),
    .B(_06925_),
    .Y(_06926_));
 sg13g2_a21oi_1 _25744_ (.A1(net999),
    .A2(_06924_),
    .Y(_06927_),
    .B1(_06926_));
 sg13g2_nand2_1 _25745_ (.Y(_06928_),
    .A(net345),
    .B(_06927_));
 sg13g2_xnor2_1 _25746_ (.Y(_06929_),
    .A(\cpu.spi.r_count[2] ),
    .B(_09002_));
 sg13g2_nor2_1 _25747_ (.A(net627),
    .B(_06929_),
    .Y(_06930_));
 sg13g2_nand2b_1 _25748_ (.Y(_06931_),
    .B(net80),
    .A_N(_06927_));
 sg13g2_o21ai_1 _25749_ (.B1(_06931_),
    .Y(_06932_),
    .A1(net70),
    .A2(_06929_));
 sg13g2_a22oi_1 _25750_ (.Y(_06933_),
    .B1(_06932_),
    .B2(net925),
    .A2(_06930_),
    .A1(_06928_));
 sg13g2_nand2_1 _25751_ (.Y(_06934_),
    .A(_06884_),
    .B(_06933_));
 sg13g2_o21ai_1 _25752_ (.B1(_06934_),
    .Y(_06935_),
    .A1(net453),
    .A2(_06922_));
 sg13g2_nand2_1 _25753_ (.Y(_06936_),
    .A(\cpu.spi.r_count[2] ),
    .B(_06874_));
 sg13g2_o21ai_1 _25754_ (.B1(_06936_),
    .Y(_02577_),
    .A1(net30),
    .A2(_06935_));
 sg13g2_nand2b_1 _25755_ (.Y(_06937_),
    .B(net389),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _25756_ (.B1(_06937_),
    .Y(_06938_),
    .A1(net366),
    .A2(_05415_));
 sg13g2_mux2_1 _25757_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net424),
    .X(_06939_));
 sg13g2_nor2_1 _25758_ (.A(net644),
    .B(_06939_),
    .Y(_06940_));
 sg13g2_a21oi_1 _25759_ (.A1(net644),
    .A2(_06938_),
    .Y(_06941_),
    .B1(_06940_));
 sg13g2_xor2_1 _25760_ (.B(_09003_),
    .A(_09000_),
    .X(_06942_));
 sg13g2_nor2_1 _25761_ (.A(net627),
    .B(_06942_),
    .Y(_06943_));
 sg13g2_nor2_1 _25762_ (.A(net998),
    .B(_05415_),
    .Y(_06944_));
 sg13g2_a21oi_1 _25763_ (.A1(net867),
    .A2(_00115_),
    .Y(_06945_),
    .B1(_06944_));
 sg13g2_mux2_1 _25764_ (.A0(_00115_),
    .A1(_00114_),
    .S(net996),
    .X(_06946_));
 sg13g2_nor2_1 _25765_ (.A(net997),
    .B(_06946_),
    .Y(_06947_));
 sg13g2_a21oi_1 _25766_ (.A1(net999),
    .A2(_06945_),
    .Y(_06948_),
    .B1(_06947_));
 sg13g2_nand2_1 _25767_ (.Y(_06949_),
    .A(net377),
    .B(_06948_));
 sg13g2_nand2b_1 _25768_ (.Y(_06950_),
    .B(net80),
    .A_N(_06948_));
 sg13g2_o21ai_1 _25769_ (.B1(_06950_),
    .Y(_06951_),
    .A1(net70),
    .A2(_06942_));
 sg13g2_a22oi_1 _25770_ (.Y(_06952_),
    .B1(_06951_),
    .B2(net925),
    .A2(_06949_),
    .A1(_06943_));
 sg13g2_nand2_1 _25771_ (.Y(_06953_),
    .A(_06883_),
    .B(_06952_));
 sg13g2_o21ai_1 _25772_ (.B1(_06953_),
    .Y(_06954_),
    .A1(net453),
    .A2(_06941_));
 sg13g2_nand2_1 _25773_ (.Y(_06955_),
    .A(_09000_),
    .B(_06874_));
 sg13g2_o21ai_1 _25774_ (.B1(_06955_),
    .Y(_02578_),
    .A1(net30),
    .A2(_06954_));
 sg13g2_nand2b_1 _25775_ (.Y(_06956_),
    .B(net389),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _25776_ (.B1(_06956_),
    .Y(_06957_),
    .A1(net389),
    .A2(_05516_));
 sg13g2_mux2_1 _25777_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net424),
    .X(_06958_));
 sg13g2_nor2_1 _25778_ (.A(net731),
    .B(_06958_),
    .Y(_06959_));
 sg13g2_a21oi_1 _25779_ (.A1(net644),
    .A2(_06957_),
    .Y(_06960_),
    .B1(_06959_));
 sg13g2_nor2_1 _25780_ (.A(_09000_),
    .B(_09003_),
    .Y(_06961_));
 sg13g2_xnor2_1 _25781_ (.Y(_06962_),
    .A(\cpu.spi.r_count[4] ),
    .B(_06961_));
 sg13g2_nor2_1 _25782_ (.A(net627),
    .B(_06962_),
    .Y(_06963_));
 sg13g2_nor2_1 _25783_ (.A(net998),
    .B(_05516_),
    .Y(_06964_));
 sg13g2_a21oi_1 _25784_ (.A1(net867),
    .A2(_00126_),
    .Y(_06965_),
    .B1(_06964_));
 sg13g2_mux2_1 _25785_ (.A0(_00126_),
    .A1(_00125_),
    .S(net996),
    .X(_06966_));
 sg13g2_nor2_1 _25786_ (.A(net997),
    .B(_06966_),
    .Y(_06967_));
 sg13g2_a21oi_1 _25787_ (.A1(net999),
    .A2(_06965_),
    .Y(_06968_),
    .B1(_06967_));
 sg13g2_nand2_1 _25788_ (.Y(_06969_),
    .A(net377),
    .B(_06968_));
 sg13g2_nand2b_1 _25789_ (.Y(_06970_),
    .B(net80),
    .A_N(_06968_));
 sg13g2_o21ai_1 _25790_ (.B1(_06970_),
    .Y(_06971_),
    .A1(net70),
    .A2(_06962_));
 sg13g2_a22oi_1 _25791_ (.Y(_06972_),
    .B1(_06971_),
    .B2(net925),
    .A2(_06969_),
    .A1(_06963_));
 sg13g2_nand2_1 _25792_ (.Y(_06973_),
    .A(_06883_),
    .B(_06972_));
 sg13g2_o21ai_1 _25793_ (.B1(_06973_),
    .Y(_06974_),
    .A1(net453),
    .A2(_06960_));
 sg13g2_nand2_1 _25794_ (.Y(_06975_),
    .A(\cpu.spi.r_count[4] ),
    .B(_06874_));
 sg13g2_o21ai_1 _25795_ (.B1(_06975_),
    .Y(_02579_),
    .A1(net30),
    .A2(_06974_));
 sg13g2_nand2b_1 _25796_ (.Y(_06976_),
    .B(net389),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _25797_ (.B1(_06976_),
    .Y(_06977_),
    .A1(net389),
    .A2(_05557_));
 sg13g2_mux2_1 _25798_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net424),
    .X(_06978_));
 sg13g2_nor2_1 _25799_ (.A(net731),
    .B(_06978_),
    .Y(_06979_));
 sg13g2_a21oi_1 _25800_ (.A1(net644),
    .A2(_06977_),
    .Y(_06980_),
    .B1(_06979_));
 sg13g2_nor2_1 _25801_ (.A(net996),
    .B(_05557_),
    .Y(_06981_));
 sg13g2_a21oi_1 _25802_ (.A1(net998),
    .A2(_00133_),
    .Y(_06982_),
    .B1(_06981_));
 sg13g2_mux2_1 _25803_ (.A0(_00133_),
    .A1(_00132_),
    .S(net996),
    .X(_06983_));
 sg13g2_nor2_1 _25804_ (.A(net997),
    .B(_06983_),
    .Y(_06984_));
 sg13g2_a21oi_1 _25805_ (.A1(net999),
    .A2(_06982_),
    .Y(_06985_),
    .B1(_06984_));
 sg13g2_nand2_1 _25806_ (.Y(_06986_),
    .A(net345),
    .B(_06985_));
 sg13g2_xnor2_1 _25807_ (.Y(_06987_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09004_));
 sg13g2_nor2_1 _25808_ (.A(net627),
    .B(_06987_),
    .Y(_06988_));
 sg13g2_nand2b_1 _25809_ (.Y(_06989_),
    .B(net80),
    .A_N(_06985_));
 sg13g2_o21ai_1 _25810_ (.B1(_06989_),
    .Y(_06990_),
    .A1(net70),
    .A2(_06987_));
 sg13g2_a22oi_1 _25811_ (.Y(_06991_),
    .B1(_06990_),
    .B2(net925),
    .A2(_06988_),
    .A1(_06986_));
 sg13g2_nand2_1 _25812_ (.Y(_06992_),
    .A(_06883_),
    .B(_06991_));
 sg13g2_o21ai_1 _25813_ (.B1(_06992_),
    .Y(_06993_),
    .A1(net453),
    .A2(_06980_));
 sg13g2_nand2_1 _25814_ (.Y(_06994_),
    .A(\cpu.spi.r_count[5] ),
    .B(_06874_));
 sg13g2_o21ai_1 _25815_ (.B1(_06994_),
    .Y(_02580_),
    .A1(net30),
    .A2(_06993_));
 sg13g2_nand2b_1 _25816_ (.Y(_06995_),
    .B(_06876_),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _25817_ (.B1(_06995_),
    .Y(_06996_),
    .A1(_06876_),
    .A2(_05647_));
 sg13g2_mux2_1 _25818_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net424),
    .X(_06997_));
 sg13g2_nor2_1 _25819_ (.A(net731),
    .B(_06997_),
    .Y(_06998_));
 sg13g2_a21oi_1 _25820_ (.A1(net644),
    .A2(_06996_),
    .Y(_06999_),
    .B1(_06998_));
 sg13g2_nor2_1 _25821_ (.A(net996),
    .B(_05647_),
    .Y(_07000_));
 sg13g2_a21oi_1 _25822_ (.A1(net998),
    .A2(_00145_),
    .Y(_07001_),
    .B1(_07000_));
 sg13g2_mux2_1 _25823_ (.A0(_00145_),
    .A1(_00144_),
    .S(_11693_),
    .X(_07002_));
 sg13g2_nor2_1 _25824_ (.A(net997),
    .B(_07002_),
    .Y(_07003_));
 sg13g2_a21oi_1 _25825_ (.A1(net999),
    .A2(_07001_),
    .Y(_07004_),
    .B1(_07003_));
 sg13g2_nand2_1 _25826_ (.Y(_07005_),
    .A(net377),
    .B(_07004_));
 sg13g2_xnor2_1 _25827_ (.Y(_07006_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09005_));
 sg13g2_nor2_1 _25828_ (.A(net627),
    .B(_07006_),
    .Y(_07007_));
 sg13g2_nand2b_1 _25829_ (.Y(_07008_),
    .B(net80),
    .A_N(_07004_));
 sg13g2_o21ai_1 _25830_ (.B1(_07008_),
    .Y(_07009_),
    .A1(net70),
    .A2(_07006_));
 sg13g2_a22oi_1 _25831_ (.Y(_07010_),
    .B1(_07009_),
    .B2(net925),
    .A2(_07007_),
    .A1(_07005_));
 sg13g2_nand2_1 _25832_ (.Y(_07011_),
    .A(_06883_),
    .B(_07010_));
 sg13g2_o21ai_1 _25833_ (.B1(_07011_),
    .Y(_07012_),
    .A1(_06884_),
    .A2(_06999_));
 sg13g2_nand2_1 _25834_ (.Y(_07013_),
    .A(\cpu.spi.r_count[6] ),
    .B(_06874_));
 sg13g2_o21ai_1 _25835_ (.B1(_07013_),
    .Y(_02581_),
    .A1(net30),
    .A2(_07012_));
 sg13g2_nand2b_1 _25836_ (.Y(_07014_),
    .B(net489),
    .A_N(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_o21ai_1 _25837_ (.B1(_07014_),
    .Y(_07015_),
    .A1(net489),
    .A2(_05012_));
 sg13g2_mux2_1 _25838_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(net489),
    .X(_07016_));
 sg13g2_nor2_1 _25839_ (.A(net864),
    .B(_07016_),
    .Y(_07017_));
 sg13g2_a21oi_1 _25840_ (.A1(net731),
    .A2(_07015_),
    .Y(_07018_),
    .B1(_07017_));
 sg13g2_nor2_1 _25841_ (.A(_06883_),
    .B(_07018_),
    .Y(_07019_));
 sg13g2_nor2_1 _25842_ (.A(_11693_),
    .B(_05012_),
    .Y(_07020_));
 sg13g2_a21oi_1 _25843_ (.A1(_11694_),
    .A2(_00157_),
    .Y(_07021_),
    .B1(_07020_));
 sg13g2_mux2_1 _25844_ (.A0(_00157_),
    .A1(_00156_),
    .S(_11693_),
    .X(_07022_));
 sg13g2_nor2_1 _25845_ (.A(_11689_),
    .B(_07022_),
    .Y(_07023_));
 sg13g2_a21oi_1 _25846_ (.A1(net997),
    .A2(_07021_),
    .Y(_07024_),
    .B1(_07023_));
 sg13g2_nor2_1 _25847_ (.A(_09192_),
    .B(_09140_),
    .Y(_07025_));
 sg13g2_a21oi_1 _25848_ (.A1(_09192_),
    .A2(_07024_),
    .Y(_07026_),
    .B1(_07025_));
 sg13g2_nor2_1 _25849_ (.A(_08999_),
    .B(_07024_),
    .Y(_07027_));
 sg13g2_nor2b_1 _25850_ (.A(_09007_),
    .B_N(_08999_),
    .Y(_07028_));
 sg13g2_a21oi_1 _25851_ (.A1(_09007_),
    .A2(_07027_),
    .Y(_07029_),
    .B1(_07028_));
 sg13g2_o21ai_1 _25852_ (.B1(_06883_),
    .Y(_07030_),
    .A1(net627),
    .A2(_07029_));
 sg13g2_a21oi_1 _25853_ (.A1(_06894_),
    .A2(_07026_),
    .Y(_07031_),
    .B1(_07030_));
 sg13g2_or2_1 _25854_ (.X(_07032_),
    .B(_07031_),
    .A(_07019_));
 sg13g2_nor3_1 _25855_ (.A(_09007_),
    .B(_09135_),
    .C(_07019_),
    .Y(_07033_));
 sg13g2_o21ai_1 _25856_ (.B1(_08999_),
    .Y(_07034_),
    .A1(_06874_),
    .A2(_07033_));
 sg13g2_o21ai_1 _25857_ (.B1(_07034_),
    .Y(_02582_),
    .A1(_06875_),
    .A2(_07032_));
 sg13g2_inv_1 _25858_ (.Y(_07035_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_mux4_1 _25859_ (.S0(_05503_),
    .A0(_09051_),
    .A1(_09043_),
    .A2(_09065_),
    .A3(_09061_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07036_));
 sg13g2_nand2_1 _25860_ (.Y(_07037_),
    .A(_09057_),
    .B(_05503_));
 sg13g2_nand2b_1 _25861_ (.Y(_07038_),
    .B(_09052_),
    .A_N(_05503_));
 sg13g2_nand3_1 _25862_ (.B(_07037_),
    .C(_07038_),
    .A(_06247_),
    .Y(_07039_));
 sg13g2_o21ai_1 _25863_ (.B1(_07039_),
    .Y(_07040_),
    .A1(_06247_),
    .A2(_07036_));
 sg13g2_nand2b_1 _25864_ (.Y(_07041_),
    .B(_05503_),
    .A_N(_09048_));
 sg13g2_o21ai_1 _25865_ (.B1(_07041_),
    .Y(_07042_),
    .A1(_09047_),
    .A2(_05503_));
 sg13g2_a21o_1 _25866_ (.A2(_07042_),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B1(_00150_),
    .X(_07043_));
 sg13g2_mux4_1 _25867_ (.S0(_05503_),
    .A0(_09045_),
    .A1(_09055_),
    .A2(_09067_),
    .A3(_09063_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07044_));
 sg13g2_nor3_1 _25868_ (.A(_07035_),
    .B(_06247_),
    .C(_07044_),
    .Y(_07045_));
 sg13g2_a221oi_1 _25869_ (.B2(_06247_),
    .C1(_07045_),
    .B1(_07043_),
    .A1(_07035_),
    .Y(_07046_),
    .A2(_07040_));
 sg13g2_mux4_1 _25870_ (.S0(_04933_),
    .A0(_09045_),
    .A1(_09055_),
    .A2(_09067_),
    .A3(_09063_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07047_));
 sg13g2_nand2_1 _25871_ (.Y(_07048_),
    .A(_09048_),
    .B(_04933_));
 sg13g2_nand2b_1 _25872_ (.Y(_07049_),
    .B(_09047_),
    .A_N(_04933_));
 sg13g2_nand3_1 _25873_ (.B(_07048_),
    .C(_07049_),
    .A(_06246_),
    .Y(_07050_));
 sg13g2_o21ai_1 _25874_ (.B1(_07050_),
    .Y(_07051_),
    .A1(_06246_),
    .A2(_07047_));
 sg13g2_mux2_1 _25875_ (.A0(_09052_),
    .A1(_09057_),
    .S(_04933_),
    .X(_07052_));
 sg13g2_inv_1 _25876_ (.Y(_07053_),
    .A(_00110_));
 sg13g2_o21ai_1 _25877_ (.B1(_07053_),
    .Y(_07054_),
    .A1(_06245_),
    .A2(_07052_));
 sg13g2_mux4_1 _25878_ (.S0(_04933_),
    .A0(_09051_),
    .A1(_09043_),
    .A2(_09065_),
    .A3(_09061_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07055_));
 sg13g2_nor3_1 _25879_ (.A(_06245_),
    .B(_06246_),
    .C(_07055_),
    .Y(_07056_));
 sg13g2_a221oi_1 _25880_ (.B2(_06246_),
    .C1(_07056_),
    .B1(_07054_),
    .A1(_06245_),
    .Y(_07057_),
    .A2(_07051_));
 sg13g2_mux2_1 _25881_ (.A0(_07046_),
    .A1(_07057_),
    .S(_11701_),
    .X(_07058_));
 sg13g2_nor2_1 _25882_ (.A(net1105),
    .B(_11746_),
    .Y(_07059_));
 sg13g2_nor2b_1 _25883_ (.A(net1029),
    .B_N(net1105),
    .Y(_07060_));
 sg13g2_a22oi_1 _25884_ (.Y(_07061_),
    .B1(_07060_),
    .B2(net602),
    .A2(_07059_),
    .A1(_09137_));
 sg13g2_nand3b_1 _25885_ (.B(net345),
    .C(net897),
    .Y(_07062_),
    .A_N(_07061_));
 sg13g2_buf_4 _25886_ (.X(_07063_),
    .A(_07062_));
 sg13g2_mux2_1 _25887_ (.A0(_07058_),
    .A1(_09163_),
    .S(_07063_),
    .X(_02586_));
 sg13g2_mux2_1 _25888_ (.A0(_09163_),
    .A1(_09162_),
    .S(_07063_),
    .X(_02587_));
 sg13g2_mux2_1 _25889_ (.A0(_09162_),
    .A1(_09166_),
    .S(_07063_),
    .X(_02588_));
 sg13g2_mux2_1 _25890_ (.A0(_09166_),
    .A1(_09160_),
    .S(_07063_),
    .X(_02589_));
 sg13g2_mux2_1 _25891_ (.A0(_09160_),
    .A1(_09168_),
    .S(_07063_),
    .X(_02590_));
 sg13g2_mux2_1 _25892_ (.A0(_09168_),
    .A1(_09167_),
    .S(_07063_),
    .X(_02591_));
 sg13g2_mux2_1 _25893_ (.A0(_09167_),
    .A1(_09161_),
    .S(_07063_),
    .X(_02592_));
 sg13g2_mux2_1 _25894_ (.A0(_09161_),
    .A1(\cpu.spi.r_in[7] ),
    .S(_07063_),
    .X(_02593_));
 sg13g2_nor3_2 _25895_ (.A(_05098_),
    .B(net551),
    .C(_00228_),
    .Y(_07064_));
 sg13g2_and4_1 _25896_ (.A(net865),
    .B(net712),
    .C(_09133_),
    .D(_07064_),
    .X(_07065_));
 sg13g2_buf_1 _25897_ (.A(_07065_),
    .X(_07066_));
 sg13g2_mux2_1 _25898_ (.A0(\cpu.spi.r_mode[0][0] ),
    .A1(_11930_),
    .S(_07066_),
    .X(_02595_));
 sg13g2_mux2_1 _25899_ (.A0(_11705_),
    .A1(net859),
    .S(_07066_),
    .X(_02596_));
 sg13g2_nand4_1 _25900_ (.B(net366),
    .C(_09133_),
    .A(net865),
    .Y(_07067_),
    .D(_07064_));
 sg13g2_buf_1 _25901_ (.A(_07067_),
    .X(_07068_));
 sg13g2_mux2_1 _25902_ (.A0(net884),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_07068_),
    .X(_02597_));
 sg13g2_mux2_1 _25903_ (.A0(net883),
    .A1(_11706_),
    .S(_07068_),
    .X(_02598_));
 sg13g2_nand3_1 _25904_ (.B(_11721_),
    .C(_07064_),
    .A(_09133_),
    .Y(_07069_));
 sg13g2_buf_1 _25905_ (.A(_07069_),
    .X(_07070_));
 sg13g2_mux2_1 _25906_ (.A0(net884),
    .A1(\cpu.spi.r_mode[2][0] ),
    .S(_07070_),
    .X(_02599_));
 sg13g2_mux2_1 _25907_ (.A0(net883),
    .A1(_11710_),
    .S(_07070_),
    .X(_02600_));
 sg13g2_nor2b_1 _25908_ (.A(net602),
    .B_N(_00223_),
    .Y(_07071_));
 sg13g2_o21ai_1 _25909_ (.B1(net925),
    .Y(_07072_),
    .A1(_06866_),
    .A2(_07071_));
 sg13g2_o21ai_1 _25910_ (.B1(_07072_),
    .Y(_07073_),
    .A1(_09190_),
    .A2(_09895_));
 sg13g2_nand2_1 _25911_ (.Y(_07074_),
    .A(_11688_),
    .B(_07073_));
 sg13g2_nor2_1 _25912_ (.A(_09105_),
    .B(net866),
    .Y(_07075_));
 sg13g2_buf_2 _25913_ (.A(_07075_),
    .X(_07076_));
 sg13g2_a221oi_1 _25914_ (.B2(_06867_),
    .C1(_11752_),
    .B1(_07076_),
    .A1(_09177_),
    .Y(_07077_),
    .A2(_11747_));
 sg13g2_o21ai_1 _25915_ (.B1(_09121_),
    .Y(_07078_),
    .A1(_09116_),
    .A2(_09114_));
 sg13g2_and2_1 _25916_ (.A(_07077_),
    .B(_07078_),
    .X(_07079_));
 sg13g2_buf_4 _25917_ (.X(_07080_),
    .A(_07079_));
 sg13g2_mux2_1 _25918_ (.A0(\cpu.spi.r_out[0] ),
    .A1(_07074_),
    .S(_07080_),
    .X(_02601_));
 sg13g2_buf_1 _25919_ (.A(_09106_),
    .X(_07081_));
 sg13g2_mux2_1 _25920_ (.A0(_00178_),
    .A1(_00223_),
    .S(net602),
    .X(_07082_));
 sg13g2_a22oi_1 _25921_ (.Y(_07083_),
    .B1(_07076_),
    .B2(_09904_),
    .A2(net866),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _25922_ (.B1(_07083_),
    .Y(_07084_),
    .A1(net801),
    .A2(_07082_));
 sg13g2_mux2_1 _25923_ (.A0(\cpu.spi.r_out[1] ),
    .A1(_07084_),
    .S(_07080_),
    .X(_02602_));
 sg13g2_mux2_1 _25924_ (.A0(_00179_),
    .A1(_00178_),
    .S(net602),
    .X(_07085_));
 sg13g2_a22oi_1 _25925_ (.Y(_07086_),
    .B1(_07076_),
    .B2(net1018),
    .A2(net866),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _25926_ (.B1(_07086_),
    .Y(_07087_),
    .A1(net801),
    .A2(_07085_));
 sg13g2_mux2_1 _25927_ (.A0(\cpu.spi.r_out[2] ),
    .A1(_07087_),
    .S(_07080_),
    .X(_02603_));
 sg13g2_mux2_1 _25928_ (.A0(_00287_),
    .A1(_00179_),
    .S(net602),
    .X(_07088_));
 sg13g2_a22oi_1 _25929_ (.Y(_07089_),
    .B1(_07076_),
    .B2(net1098),
    .A2(net866),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _25930_ (.B1(_07089_),
    .Y(_07090_),
    .A1(net801),
    .A2(_07088_));
 sg13g2_mux2_1 _25931_ (.A0(\cpu.spi.r_out[3] ),
    .A1(_07090_),
    .S(_07080_),
    .X(_02604_));
 sg13g2_mux2_1 _25932_ (.A0(_00180_),
    .A1(_00287_),
    .S(net602),
    .X(_07091_));
 sg13g2_a22oi_1 _25933_ (.Y(_07092_),
    .B1(_07076_),
    .B2(_09921_),
    .A2(net866),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _25934_ (.B1(_07092_),
    .Y(_07093_),
    .A1(net801),
    .A2(_07091_));
 sg13g2_mux2_1 _25935_ (.A0(\cpu.spi.r_out[4] ),
    .A1(_07093_),
    .S(_07080_),
    .X(_02605_));
 sg13g2_mux2_1 _25936_ (.A0(_00181_),
    .A1(_00180_),
    .S(_11753_),
    .X(_07094_));
 sg13g2_a22oi_1 _25937_ (.Y(_07095_),
    .B1(_07076_),
    .B2(_09927_),
    .A2(net866),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _25938_ (.B1(_07095_),
    .Y(_07096_),
    .A1(net801),
    .A2(_07094_));
 sg13g2_mux2_1 _25939_ (.A0(\cpu.spi.r_out[5] ),
    .A1(_07096_),
    .S(_07080_),
    .X(_02606_));
 sg13g2_buf_1 _25940_ (.A(_00182_),
    .X(_07097_));
 sg13g2_mux2_1 _25941_ (.A0(_07097_),
    .A1(_00181_),
    .S(_11753_),
    .X(_07098_));
 sg13g2_a22oi_1 _25942_ (.Y(_07099_),
    .B1(_07076_),
    .B2(_09933_),
    .A2(net866),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _25943_ (.B1(_07099_),
    .Y(_07100_),
    .A1(_07081_),
    .A2(_07098_));
 sg13g2_mux2_1 _25944_ (.A0(\cpu.spi.r_out[6] ),
    .A1(_07100_),
    .S(_07080_),
    .X(_02607_));
 sg13g2_buf_1 _25945_ (.A(_00281_),
    .X(_07101_));
 sg13g2_mux2_1 _25946_ (.A0(_07101_),
    .A1(_07097_),
    .S(net602),
    .X(_07102_));
 sg13g2_a22oi_1 _25947_ (.Y(_07103_),
    .B1(_07076_),
    .B2(_09940_),
    .A2(_11714_),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _25948_ (.B1(_07103_),
    .Y(_07104_),
    .A1(_07081_),
    .A2(_07102_));
 sg13g2_mux2_1 _25949_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_07104_),
    .S(_07080_),
    .X(_02608_));
 sg13g2_nand3_1 _25950_ (.B(net897),
    .C(_09188_),
    .A(_09116_),
    .Y(_07105_));
 sg13g2_buf_1 _25951_ (.A(_07105_),
    .X(_07106_));
 sg13g2_nand2_1 _25952_ (.Y(_07107_),
    .A(net867),
    .B(_07106_));
 sg13g2_o21ai_1 _25953_ (.B1(_07107_),
    .Y(_02611_),
    .A1(_03703_),
    .A2(_07106_));
 sg13g2_nand2_1 _25954_ (.Y(_07108_),
    .A(_11690_),
    .B(_07106_));
 sg13g2_o21ai_1 _25955_ (.B1(_07108_),
    .Y(_02612_),
    .A1(_06178_),
    .A2(_07106_));
 sg13g2_mux2_1 _25956_ (.A0(\cpu.spi.r_src[0] ),
    .A1(net858),
    .S(_07066_),
    .X(_02613_));
 sg13g2_mux2_1 _25957_ (.A0(net862),
    .A1(\cpu.spi.r_src[1] ),
    .S(_07068_),
    .X(_02614_));
 sg13g2_mux2_1 _25958_ (.A0(net862),
    .A1(_11691_),
    .S(_07070_),
    .X(_02615_));
 sg13g2_and2_1 _25959_ (.A(_09133_),
    .B(_05014_),
    .X(_07109_));
 sg13g2_buf_4 _25960_ (.X(_07110_),
    .A(_07109_));
 sg13g2_mux2_1 _25961_ (.A0(\cpu.spi.r_timeout[0] ),
    .A1(net861),
    .S(_07110_),
    .X(_02616_));
 sg13g2_mux2_1 _25962_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(net859),
    .S(_07110_),
    .X(_02617_));
 sg13g2_mux2_1 _25963_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(net858),
    .S(_07110_),
    .X(_02618_));
 sg13g2_mux2_1 _25964_ (.A0(\cpu.spi.r_timeout[3] ),
    .A1(net982),
    .S(_07110_),
    .X(_02619_));
 sg13g2_mux2_1 _25965_ (.A0(\cpu.spi.r_timeout[4] ),
    .A1(net981),
    .S(_07110_),
    .X(_02620_));
 sg13g2_mux2_1 _25966_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(net980),
    .S(_07110_),
    .X(_02621_));
 sg13g2_mux2_1 _25967_ (.A0(\cpu.spi.r_timeout[6] ),
    .A1(net979),
    .S(_07110_),
    .X(_02622_));
 sg13g2_mux2_1 _25968_ (.A0(\cpu.spi.r_timeout[7] ),
    .A1(net978),
    .S(_07110_),
    .X(_02623_));
 sg13g2_nand2_1 _25969_ (.Y(_07111_),
    .A(_09136_),
    .B(_09172_));
 sg13g2_or3_1 _25970_ (.A(_00226_),
    .B(_09144_),
    .C(_09172_),
    .X(_07112_));
 sg13g2_nand3_1 _25971_ (.B(_07111_),
    .C(_07112_),
    .A(_09139_),
    .Y(_07113_));
 sg13g2_nand2_1 _25972_ (.Y(_07114_),
    .A(_09106_),
    .B(_09136_));
 sg13g2_o21ai_1 _25973_ (.B1(_07113_),
    .Y(_07115_),
    .A1(_09136_),
    .A2(_09139_));
 sg13g2_nand3_1 _25974_ (.B(_09113_),
    .C(_07115_),
    .A(_09105_),
    .Y(_07116_));
 sg13g2_o21ai_1 _25975_ (.B1(_07116_),
    .Y(_07117_),
    .A1(_07113_),
    .A2(_07114_));
 sg13g2_nand2_1 _25976_ (.Y(_07118_),
    .A(net897),
    .B(_07117_));
 sg13g2_buf_2 _25977_ (.A(_07118_),
    .X(_07119_));
 sg13g2_buf_1 _25978_ (.A(_07119_),
    .X(_07120_));
 sg13g2_and2_1 _25979_ (.A(net925),
    .B(\cpu.spi.r_timeout[0] ),
    .X(_07121_));
 sg13g2_a21oi_1 _25980_ (.A1(net801),
    .A2(_00284_),
    .Y(_07122_),
    .B1(_07121_));
 sg13g2_nand2_1 _25981_ (.Y(_07123_),
    .A(_09146_),
    .B(net29));
 sg13g2_o21ai_1 _25982_ (.B1(_07123_),
    .Y(_02624_),
    .A1(net29),
    .A2(_07122_));
 sg13g2_nor3_1 _25983_ (.A(_09146_),
    .B(_09147_),
    .C(_07119_),
    .Y(_07124_));
 sg13g2_a21oi_1 _25984_ (.A1(_09146_),
    .A2(_09147_),
    .Y(_07125_),
    .B1(_07124_));
 sg13g2_nor2_1 _25985_ (.A(_09106_),
    .B(_07119_),
    .Y(_07126_));
 sg13g2_buf_2 _25986_ (.A(_07126_),
    .X(_07127_));
 sg13g2_a22oi_1 _25987_ (.Y(_07128_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[1] ),
    .A2(net29),
    .A1(_09147_));
 sg13g2_o21ai_1 _25988_ (.B1(_07128_),
    .Y(_02625_),
    .A1(net1028),
    .A2(_07125_));
 sg13g2_o21ai_1 _25989_ (.B1(\cpu.spi.r_timeout_count[2] ),
    .Y(_07129_),
    .A1(_09146_),
    .A2(_09147_));
 sg13g2_o21ai_1 _25990_ (.B1(_07129_),
    .Y(_07130_),
    .A1(_09149_),
    .A2(_07120_));
 sg13g2_nand2_1 _25991_ (.Y(_07131_),
    .A(net801),
    .B(_07130_));
 sg13g2_a22oi_1 _25992_ (.Y(_07132_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[2] ),
    .A2(_07120_),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_nand2_1 _25993_ (.Y(_02626_),
    .A(_07131_),
    .B(_07132_));
 sg13g2_nor2_1 _25994_ (.A(_09151_),
    .B(_07119_),
    .Y(_07133_));
 sg13g2_a21oi_1 _25995_ (.A1(\cpu.spi.r_timeout_count[3] ),
    .A2(_09149_),
    .Y(_07134_),
    .B1(_07133_));
 sg13g2_a22oi_1 _25996_ (.Y(_07135_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[3] ),
    .A2(net29),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_o21ai_1 _25997_ (.B1(_07135_),
    .Y(_02627_),
    .A1(net1028),
    .A2(_07134_));
 sg13g2_nor2_1 _25998_ (.A(_09153_),
    .B(_07119_),
    .Y(_07136_));
 sg13g2_a21oi_1 _25999_ (.A1(\cpu.spi.r_timeout_count[4] ),
    .A2(_09151_),
    .Y(_07137_),
    .B1(_07136_));
 sg13g2_a22oi_1 _26000_ (.Y(_07138_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[4] ),
    .A2(net29),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_o21ai_1 _26001_ (.B1(_07138_),
    .Y(_02628_),
    .A1(net1028),
    .A2(_07137_));
 sg13g2_nor2_1 _26002_ (.A(_09155_),
    .B(_07119_),
    .Y(_07139_));
 sg13g2_a21oi_1 _26003_ (.A1(\cpu.spi.r_timeout_count[5] ),
    .A2(_09153_),
    .Y(_07140_),
    .B1(_07139_));
 sg13g2_a22oi_1 _26004_ (.Y(_07141_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[5] ),
    .A2(net29),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_o21ai_1 _26005_ (.B1(_07141_),
    .Y(_02629_),
    .A1(net1028),
    .A2(_07140_));
 sg13g2_nor2_1 _26006_ (.A(_09157_),
    .B(_07119_),
    .Y(_07142_));
 sg13g2_a21oi_1 _26007_ (.A1(\cpu.spi.r_timeout_count[6] ),
    .A2(_09155_),
    .Y(_07143_),
    .B1(_07142_));
 sg13g2_a22oi_1 _26008_ (.Y(_07144_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[6] ),
    .A2(net29),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_o21ai_1 _26009_ (.B1(_07144_),
    .Y(_02630_),
    .A1(net1028),
    .A2(_07143_));
 sg13g2_nor3_1 _26010_ (.A(_09145_),
    .B(_09157_),
    .C(_07119_),
    .Y(_07145_));
 sg13g2_a21oi_1 _26011_ (.A1(_09145_),
    .A2(_09157_),
    .Y(_07146_),
    .B1(_07145_));
 sg13g2_a22oi_1 _26012_ (.Y(_07147_),
    .B1(_07127_),
    .B2(\cpu.spi.r_timeout[7] ),
    .A2(net29),
    .A1(_09145_));
 sg13g2_o21ai_1 _26013_ (.B1(_07147_),
    .Y(_02631_),
    .A1(net1028),
    .A2(_07146_));
 sg13g2_buf_1 _26014_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07148_));
 sg13g2_nor2_1 _26015_ (.A(_07148_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07149_));
 sg13g2_nand2_1 _26016_ (.Y(_07150_),
    .A(net342),
    .B(_07149_));
 sg13g2_nor2_1 _26017_ (.A(net896),
    .B(_07150_),
    .Y(_07151_));
 sg13g2_buf_1 _26018_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07152_));
 sg13g2_buf_1 _26019_ (.A(_07152_),
    .X(_07153_));
 sg13g2_buf_1 _26020_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07154_));
 sg13g2_buf_1 _26021_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07155_));
 sg13g2_buf_1 _26022_ (.A(_07155_),
    .X(_07156_));
 sg13g2_nor2_2 _26023_ (.A(net1066),
    .B(net923),
    .Y(_07157_));
 sg13g2_buf_2 _26024_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07158_));
 sg13g2_inv_1 _26025_ (.Y(_07159_),
    .A(_07158_));
 sg13g2_nand3_1 _26026_ (.B(net924),
    .C(_07157_),
    .A(_07159_),
    .Y(_07160_));
 sg13g2_o21ai_1 _26027_ (.B1(_07160_),
    .Y(_07161_),
    .A1(net924),
    .A2(_07157_));
 sg13g2_and2_1 _26028_ (.A(_07151_),
    .B(_07161_),
    .X(_07162_));
 sg13g2_buf_2 _26029_ (.A(_07162_),
    .X(_07163_));
 sg13g2_mux2_1 _26030_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07163_),
    .X(_02644_));
 sg13g2_mux2_1 _26031_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07163_),
    .X(_02645_));
 sg13g2_mux2_1 _26032_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07163_),
    .X(_02646_));
 sg13g2_mux2_1 _26033_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07163_),
    .X(_02647_));
 sg13g2_mux2_1 _26034_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07163_),
    .X(_02648_));
 sg13g2_mux2_1 _26035_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07163_),
    .X(_02649_));
 sg13g2_xor2_1 _26036_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07164_));
 sg13g2_mux2_1 _26037_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07164_),
    .S(_07163_),
    .X(_02650_));
 sg13g2_and4_1 _26038_ (.A(_07158_),
    .B(net924),
    .C(_07151_),
    .D(_07157_),
    .X(_07165_));
 sg13g2_buf_1 _26039_ (.A(_07165_),
    .X(_07166_));
 sg13g2_mux2_1 _26040_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net173),
    .X(_02651_));
 sg13g2_mux2_1 _26041_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net173),
    .X(_02652_));
 sg13g2_mux2_1 _26042_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net173),
    .X(_02653_));
 sg13g2_mux2_1 _26043_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net173),
    .X(_02654_));
 sg13g2_mux2_1 _26044_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net173),
    .X(_02655_));
 sg13g2_mux2_1 _26045_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net173),
    .X(_02656_));
 sg13g2_mux2_1 _26046_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net173),
    .X(_02657_));
 sg13g2_mux2_1 _26047_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07164_),
    .S(net173),
    .X(_02658_));
 sg13g2_nor2_1 _26048_ (.A(net1038),
    .B(net1037),
    .Y(_07167_));
 sg13g2_nand3_1 _26049_ (.B(_07167_),
    .C(_06234_),
    .A(net995),
    .Y(_07168_));
 sg13g2_nor2_2 _26050_ (.A(_05489_),
    .B(_07168_),
    .Y(_07169_));
 sg13g2_buf_1 _26051_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07170_));
 sg13g2_buf_1 _26052_ (.A(_07170_),
    .X(_07171_));
 sg13g2_buf_2 _26053_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07172_));
 sg13g2_inv_1 _26054_ (.Y(_07173_),
    .A(_07172_));
 sg13g2_buf_1 _26055_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07174_));
 sg13g2_inv_1 _26056_ (.Y(_07175_),
    .A(_07174_));
 sg13g2_buf_1 _26057_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07176_));
 sg13g2_nor3_2 _26058_ (.A(_07173_),
    .B(_07175_),
    .C(_07176_),
    .Y(_07177_));
 sg13g2_buf_1 _26059_ (.A(_07174_),
    .X(_07178_));
 sg13g2_or2_1 _26060_ (.X(_07179_),
    .B(_07170_),
    .A(_07172_));
 sg13g2_buf_1 _26061_ (.A(_07179_),
    .X(_07180_));
 sg13g2_nor3_1 _26062_ (.A(net921),
    .B(_07176_),
    .C(_07180_),
    .Y(_07181_));
 sg13g2_a21oi_1 _26063_ (.A1(_07171_),
    .A2(_07177_),
    .Y(_07182_),
    .B1(_07181_));
 sg13g2_nor2_1 _26064_ (.A(_07172_),
    .B(_07176_),
    .Y(_07183_));
 sg13g2_xnor2_1 _26065_ (.Y(_07184_),
    .A(net921),
    .B(_07183_));
 sg13g2_buf_1 _26066_ (.A(_07184_),
    .X(_07185_));
 sg13g2_inv_2 _26067_ (.Y(_07186_),
    .A(net695));
 sg13g2_buf_1 _26068_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07187_));
 sg13g2_nor2_2 _26069_ (.A(_07187_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07188_));
 sg13g2_nand2_1 _26070_ (.Y(_07189_),
    .A(_09780_),
    .B(_07188_));
 sg13g2_buf_1 _26071_ (.A(_07189_),
    .X(_07190_));
 sg13g2_o21ai_1 _26072_ (.B1(_07182_),
    .Y(_07191_),
    .A1(_07186_),
    .A2(_07190_));
 sg13g2_and2_1 _26073_ (.A(net897),
    .B(_07191_),
    .X(_07192_));
 sg13g2_o21ai_1 _26074_ (.B1(_07192_),
    .Y(_07193_),
    .A1(_07169_),
    .A2(_07182_));
 sg13g2_buf_2 _26075_ (.A(_07193_),
    .X(_07194_));
 sg13g2_buf_1 _26076_ (.A(_07194_),
    .X(_07195_));
 sg13g2_and2_1 _26077_ (.A(\cpu.uart.r_out[1] ),
    .B(net695),
    .X(_07196_));
 sg13g2_a21oi_1 _26078_ (.A1(net1020),
    .A2(_07186_),
    .Y(_07197_),
    .B1(_07196_));
 sg13g2_nand2_1 _26079_ (.Y(_07198_),
    .A(\cpu.uart.r_out[0] ),
    .B(net62));
 sg13g2_o21ai_1 _26080_ (.B1(_07198_),
    .Y(_02659_),
    .A1(net62),
    .A2(_07197_));
 sg13g2_and2_1 _26081_ (.A(\cpu.uart.r_out[2] ),
    .B(_07185_),
    .X(_07199_));
 sg13g2_a21oi_1 _26082_ (.A1(net1019),
    .A2(_07186_),
    .Y(_07200_),
    .B1(_07199_));
 sg13g2_nand2_1 _26083_ (.Y(_07201_),
    .A(\cpu.uart.r_out[1] ),
    .B(net62));
 sg13g2_o21ai_1 _26084_ (.B1(_07201_),
    .Y(_02660_),
    .A1(net62),
    .A2(_07200_));
 sg13g2_and2_1 _26085_ (.A(\cpu.uart.r_out[3] ),
    .B(net695),
    .X(_07202_));
 sg13g2_a21oi_1 _26086_ (.A1(net1018),
    .A2(_07186_),
    .Y(_07203_),
    .B1(_07202_));
 sg13g2_nand2_1 _26087_ (.Y(_07204_),
    .A(\cpu.uart.r_out[2] ),
    .B(_07194_));
 sg13g2_o21ai_1 _26088_ (.B1(_07204_),
    .Y(_02661_),
    .A1(_07195_),
    .A2(_07203_));
 sg13g2_and2_1 _26089_ (.A(\cpu.uart.r_out[4] ),
    .B(net695),
    .X(_07205_));
 sg13g2_a21oi_1 _26090_ (.A1(net1098),
    .A2(_07186_),
    .Y(_07206_),
    .B1(_07205_));
 sg13g2_nand2_1 _26091_ (.Y(_07207_),
    .A(\cpu.uart.r_out[3] ),
    .B(_07194_));
 sg13g2_o21ai_1 _26092_ (.B1(_07207_),
    .Y(_02662_),
    .A1(net62),
    .A2(_07206_));
 sg13g2_and2_1 _26093_ (.A(\cpu.uart.r_out[5] ),
    .B(net695),
    .X(_07208_));
 sg13g2_a21oi_1 _26094_ (.A1(net1016),
    .A2(_07186_),
    .Y(_07209_),
    .B1(_07208_));
 sg13g2_nand2_1 _26095_ (.Y(_07210_),
    .A(\cpu.uart.r_out[4] ),
    .B(_07194_));
 sg13g2_o21ai_1 _26096_ (.B1(_07210_),
    .Y(_02663_),
    .A1(net62),
    .A2(_07209_));
 sg13g2_and2_1 _26097_ (.A(\cpu.uart.r_out[6] ),
    .B(net695),
    .X(_07211_));
 sg13g2_a21oi_1 _26098_ (.A1(net1015),
    .A2(_07186_),
    .Y(_07212_),
    .B1(_07211_));
 sg13g2_nand2_1 _26099_ (.Y(_07213_),
    .A(\cpu.uart.r_out[5] ),
    .B(_07194_));
 sg13g2_o21ai_1 _26100_ (.B1(_07213_),
    .Y(_02664_),
    .A1(_07195_),
    .A2(_07212_));
 sg13g2_and2_1 _26101_ (.A(\cpu.uart.r_out[7] ),
    .B(net695),
    .X(_07214_));
 sg13g2_a21oi_1 _26102_ (.A1(net1014),
    .A2(_07186_),
    .Y(_07215_),
    .B1(_07214_));
 sg13g2_nand2_1 _26103_ (.Y(_07216_),
    .A(\cpu.uart.r_out[6] ),
    .B(_07194_));
 sg13g2_o21ai_1 _26104_ (.B1(_07216_),
    .Y(_02665_),
    .A1(net62),
    .A2(_07215_));
 sg13g2_nor3_1 _26105_ (.A(_07101_),
    .B(net695),
    .C(_07194_),
    .Y(_07217_));
 sg13g2_a21o_1 _26106_ (.A2(net62),
    .A1(\cpu.uart.r_out[7] ),
    .B1(_07217_),
    .X(_02666_));
 sg13g2_nand2b_1 _26107_ (.Y(_07218_),
    .B(_09808_),
    .A_N(_09769_));
 sg13g2_buf_1 _26108_ (.A(_07218_),
    .X(_07219_));
 sg13g2_nor3_1 _26109_ (.A(_07154_),
    .B(_07155_),
    .C(net1067),
    .Y(_07220_));
 sg13g2_a22oi_1 _26110_ (.Y(_07221_),
    .B1(_07219_),
    .B2(_07220_),
    .A2(net1067),
    .A1(net1066));
 sg13g2_nor4_1 _26111_ (.A(_07158_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_07155_),
    .D(net1067),
    .Y(_07222_));
 sg13g2_a21o_1 _26112_ (.A2(_07219_),
    .A1(_07154_),
    .B1(_07155_),
    .X(_07223_));
 sg13g2_a22oi_1 _26113_ (.Y(_07224_),
    .B1(_07223_),
    .B2(net1067),
    .A2(_07222_),
    .A1(_07164_));
 sg13g2_o21ai_1 _26114_ (.B1(_07224_),
    .Y(_07225_),
    .A1(_07159_),
    .A2(_07221_));
 sg13g2_nor2_1 _26115_ (.A(_07159_),
    .B(net1066),
    .Y(_07226_));
 sg13g2_nor2b_1 _26116_ (.A(net1067),
    .B_N(_07164_),
    .Y(_07227_));
 sg13g2_nand2_1 _26117_ (.Y(_07228_),
    .A(net1066),
    .B(net1067));
 sg13g2_nor2_1 _26118_ (.A(_07158_),
    .B(_07228_),
    .Y(_07229_));
 sg13g2_a21oi_1 _26119_ (.A1(_07226_),
    .A2(_07227_),
    .Y(_07230_),
    .B1(_07229_));
 sg13g2_nor3_1 _26120_ (.A(_07156_),
    .B(_07150_),
    .C(_07230_),
    .Y(_07231_));
 sg13g2_nor2b_1 _26121_ (.A(_07157_),
    .B_N(net924),
    .Y(_07232_));
 sg13g2_nor3_1 _26122_ (.A(net342),
    .B(_07220_),
    .C(_07232_),
    .Y(_07233_));
 sg13g2_nor4_2 _26123_ (.A(net896),
    .B(_07225_),
    .C(_07231_),
    .Y(_07234_),
    .D(_07233_));
 sg13g2_and2_1 _26124_ (.A(_07158_),
    .B(net1066),
    .X(_07235_));
 sg13g2_buf_1 _26125_ (.A(_07235_),
    .X(_07236_));
 sg13g2_o21ai_1 _26126_ (.B1(net924),
    .Y(_07237_),
    .A1(net923),
    .A2(_07236_));
 sg13g2_nor2b_1 _26127_ (.A(_07222_),
    .B_N(_07237_),
    .Y(_07238_));
 sg13g2_and2_1 _26128_ (.A(_07234_),
    .B(_07238_),
    .X(_07239_));
 sg13g2_nor2_1 _26129_ (.A(_07148_),
    .B(_07234_),
    .Y(_07240_));
 sg13g2_a21oi_1 _26130_ (.A1(_07148_),
    .A2(_07239_),
    .Y(_02669_),
    .B1(_07240_));
 sg13g2_nand2_1 _26131_ (.Y(_07241_),
    .A(_07148_),
    .B(_07238_));
 sg13g2_inv_1 _26132_ (.Y(_07242_),
    .A(\cpu.uart.r_rcnt[1] ));
 sg13g2_a21oi_1 _26133_ (.A1(_07234_),
    .A2(_07241_),
    .Y(_07243_),
    .B1(_07242_));
 sg13g2_a21o_1 _26134_ (.A2(_07239_),
    .A1(_07149_),
    .B1(_07243_),
    .X(_02670_));
 sg13g2_nand2_1 _26135_ (.Y(_07244_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07185_));
 sg13g2_xnor2_1 _26136_ (.Y(_07245_),
    .A(\cpu.uart.r_x_invert ),
    .B(_07244_));
 sg13g2_buf_1 _26137_ (.A(_07176_),
    .X(_07246_));
 sg13g2_nor2_1 _26138_ (.A(_07175_),
    .B(net920),
    .Y(_07247_));
 sg13g2_nand2_1 _26139_ (.Y(_07248_),
    .A(_07175_),
    .B(net920));
 sg13g2_nor2_1 _26140_ (.A(_07180_),
    .B(_07247_),
    .Y(_07249_));
 sg13g2_a221oi_1 _26141_ (.B2(_07249_),
    .C1(net896),
    .B1(_07248_),
    .A1(_07172_),
    .Y(_07250_),
    .A2(_07247_));
 sg13g2_mux2_1 _26142_ (.A0(_00280_),
    .A1(_07245_),
    .S(_07250_),
    .X(_07251_));
 sg13g2_buf_1 _26143_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07252_));
 sg13g2_a21oi_1 _26144_ (.A1(_07170_),
    .A2(_07178_),
    .Y(_07253_),
    .B1(_07173_));
 sg13g2_nor2_1 _26145_ (.A(_07172_),
    .B(_07170_),
    .Y(_07254_));
 sg13g2_nor2_1 _26146_ (.A(net921),
    .B(_07190_),
    .Y(_07255_));
 sg13g2_a21oi_1 _26147_ (.A1(net921),
    .A2(_07254_),
    .Y(_07256_),
    .B1(_07255_));
 sg13g2_nor2b_1 _26148_ (.A(net921),
    .B_N(_07170_),
    .Y(_07257_));
 sg13g2_a21oi_1 _26149_ (.A1(net342),
    .A2(_07188_),
    .Y(_07258_),
    .B1(_07175_));
 sg13g2_a21oi_1 _26150_ (.A1(_07219_),
    .A2(_07257_),
    .Y(_07259_),
    .B1(_07258_));
 sg13g2_nor2b_1 _26151_ (.A(_07259_),
    .B_N(_07183_),
    .Y(_07260_));
 sg13g2_a221oi_1 _26152_ (.B2(_07176_),
    .C1(_07260_),
    .B1(_07256_),
    .A1(_07190_),
    .Y(_07261_),
    .A2(_07253_));
 sg13g2_nand3_1 _26153_ (.B(_07169_),
    .C(_07177_),
    .A(_07171_),
    .Y(_07262_));
 sg13g2_buf_1 _26154_ (.A(_07262_),
    .X(_07263_));
 sg13g2_a21oi_1 _26155_ (.A1(_07261_),
    .A2(_07263_),
    .Y(_07264_),
    .B1(net779));
 sg13g2_mux2_1 _26156_ (.A0(_07251_),
    .A1(net1065),
    .S(_07264_),
    .X(_02675_));
 sg13g2_inv_1 _26157_ (.Y(_07265_),
    .A(_07263_));
 sg13g2_inv_1 _26158_ (.Y(_07266_),
    .A(_07181_));
 sg13g2_a21oi_1 _26159_ (.A1(net922),
    .A2(_07188_),
    .Y(_07267_),
    .B1(_07176_));
 sg13g2_o21ai_1 _26160_ (.B1(_07246_),
    .Y(_07268_),
    .A1(net922),
    .A2(_07188_));
 sg13g2_o21ai_1 _26161_ (.B1(_07268_),
    .Y(_07269_),
    .A1(_07173_),
    .A2(_07267_));
 sg13g2_nand2_1 _26162_ (.Y(_07270_),
    .A(_07178_),
    .B(_07269_));
 sg13g2_nand3_1 _26163_ (.B(_07266_),
    .C(_07270_),
    .A(net897),
    .Y(_07271_));
 sg13g2_nor3_1 _26164_ (.A(_07219_),
    .B(_07265_),
    .C(_07271_),
    .Y(_07272_));
 sg13g2_and2_1 _26165_ (.A(net921),
    .B(net920),
    .X(_07273_));
 sg13g2_buf_1 _26166_ (.A(_07273_),
    .X(_07274_));
 sg13g2_a22oi_1 _26167_ (.Y(_07275_),
    .B1(_07274_),
    .B2(_07180_),
    .A2(_07183_),
    .A1(_07175_));
 sg13g2_nand2_1 _26168_ (.Y(_07276_),
    .A(_07272_),
    .B(_07275_));
 sg13g2_nor2b_1 _26169_ (.A(_07187_),
    .B_N(_07272_),
    .Y(_07277_));
 sg13g2_a21oi_1 _26170_ (.A1(_07187_),
    .A2(_07276_),
    .Y(_07278_),
    .B1(_07277_));
 sg13g2_inv_1 _26171_ (.Y(_02678_),
    .A(_07278_));
 sg13g2_nand2_1 _26172_ (.Y(_07279_),
    .A(_07187_),
    .B(_07275_));
 sg13g2_nand2_1 _26173_ (.Y(_07280_),
    .A(_07272_),
    .B(_07279_));
 sg13g2_o21ai_1 _26174_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07281_),
    .A1(_07187_),
    .A2(_07276_));
 sg13g2_o21ai_1 _26175_ (.B1(_07281_),
    .Y(_02679_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07280_));
 sg13g2_nand2_1 _26176_ (.Y(_07282_),
    .A(net667),
    .B(net124));
 sg13g2_buf_1 _26177_ (.A(_07282_),
    .X(_07283_));
 sg13g2_buf_1 _26178_ (.A(_07283_),
    .X(_07284_));
 sg13g2_nand2_1 _26179_ (.Y(_07285_),
    .A(net123),
    .B(net375));
 sg13g2_buf_1 _26180_ (.A(_07285_),
    .X(_07286_));
 sg13g2_buf_1 _26181_ (.A(_07286_),
    .X(_07287_));
 sg13g2_buf_1 _26182_ (.A(_07286_),
    .X(_07288_));
 sg13g2_and4_1 _26183_ (.A(_10032_),
    .B(_10038_),
    .C(_10045_),
    .D(_10040_),
    .X(_07289_));
 sg13g2_and2_1 _26184_ (.A(_04862_),
    .B(_07289_),
    .X(_07290_));
 sg13g2_buf_1 _26185_ (.A(_07290_),
    .X(_07291_));
 sg13g2_nand2_1 _26186_ (.Y(_07292_),
    .A(net71),
    .B(_07291_));
 sg13g2_o21ai_1 _26187_ (.B1(_07292_),
    .Y(_07293_),
    .A1(_09896_),
    .A2(net72));
 sg13g2_o21ai_1 _26188_ (.B1(net82),
    .Y(_07294_),
    .A1(net78),
    .A2(_07289_));
 sg13g2_inv_1 _26189_ (.Y(_07295_),
    .A(_04862_));
 sg13g2_a22oi_1 _26190_ (.Y(_02465_),
    .B1(_07294_),
    .B2(_07295_),
    .A2(_07293_),
    .A1(net73));
 sg13g2_and2_1 _26191_ (.A(_05299_),
    .B(_07291_),
    .X(_07296_));
 sg13g2_buf_1 _26192_ (.A(_07296_),
    .X(_07297_));
 sg13g2_nand2_1 _26193_ (.Y(_07298_),
    .A(net71),
    .B(_07297_));
 sg13g2_o21ai_1 _26194_ (.B1(_07298_),
    .Y(_07299_),
    .A1(_09905_),
    .A2(net72));
 sg13g2_o21ai_1 _26195_ (.B1(net82),
    .Y(_07300_),
    .A1(net78),
    .A2(_07291_));
 sg13g2_inv_1 _26196_ (.Y(_07301_),
    .A(_05299_));
 sg13g2_a22oi_1 _26197_ (.Y(_02466_),
    .B1(_07300_),
    .B2(_07301_),
    .A2(_07299_),
    .A1(net73));
 sg13g2_and2_1 _26198_ (.A(_05380_),
    .B(_07297_),
    .X(_07302_));
 sg13g2_buf_1 _26199_ (.A(_07302_),
    .X(_07303_));
 sg13g2_nand2_1 _26200_ (.Y(_07304_),
    .A(net71),
    .B(_07303_));
 sg13g2_o21ai_1 _26201_ (.B1(_07304_),
    .Y(_07305_),
    .A1(_09910_),
    .A2(net72));
 sg13g2_o21ai_1 _26202_ (.B1(net82),
    .Y(_07306_),
    .A1(net78),
    .A2(_07297_));
 sg13g2_inv_1 _26203_ (.Y(_07307_),
    .A(_05380_));
 sg13g2_a22oi_1 _26204_ (.Y(_02467_),
    .B1(_07306_),
    .B2(_07307_),
    .A2(_07305_),
    .A1(net73));
 sg13g2_nand3_1 _26205_ (.B(_10038_),
    .C(_10045_),
    .A(_10032_),
    .Y(_07308_));
 sg13g2_nor4_1 _26206_ (.A(_07295_),
    .B(_07301_),
    .C(_07307_),
    .D(_07308_),
    .Y(_07309_));
 sg13g2_and2_1 _26207_ (.A(_10034_),
    .B(_07309_),
    .X(_07310_));
 sg13g2_buf_2 _26208_ (.A(_07310_),
    .X(_07311_));
 sg13g2_nand3_1 _26209_ (.B(_07286_),
    .C(_07311_),
    .A(_05436_),
    .Y(_07312_));
 sg13g2_o21ai_1 _26210_ (.B1(_07312_),
    .Y(_07313_),
    .A1(net1098),
    .A2(net72));
 sg13g2_o21ai_1 _26211_ (.B1(net82),
    .Y(_07314_),
    .A1(net78),
    .A2(_07311_));
 sg13g2_inv_1 _26212_ (.Y(_07315_),
    .A(_05436_));
 sg13g2_a22oi_1 _26213_ (.Y(_02468_),
    .B1(_07314_),
    .B2(_07315_),
    .A2(_07313_),
    .A1(net73));
 sg13g2_nand4_1 _26214_ (.B(_05484_),
    .C(_07286_),
    .A(_05436_),
    .Y(_07316_),
    .D(_07303_));
 sg13g2_o21ai_1 _26215_ (.B1(_07316_),
    .Y(_07317_),
    .A1(_09921_),
    .A2(net72));
 sg13g2_and2_1 _26216_ (.A(_05436_),
    .B(_07303_),
    .X(_07318_));
 sg13g2_o21ai_1 _26217_ (.B1(net82),
    .Y(_07319_),
    .A1(net78),
    .A2(_07318_));
 sg13g2_inv_1 _26218_ (.Y(_07320_),
    .A(_05484_));
 sg13g2_a22oi_1 _26219_ (.Y(_02469_),
    .B1(_07319_),
    .B2(_07320_),
    .A2(_07317_),
    .A1(net73));
 sg13g2_and3_1 _26220_ (.X(_07321_),
    .A(_05436_),
    .B(_05484_),
    .C(_05583_));
 sg13g2_buf_1 _26221_ (.A(_07321_),
    .X(_07322_));
 sg13g2_nand3_1 _26222_ (.B(_07311_),
    .C(_07322_),
    .A(net71),
    .Y(_07323_));
 sg13g2_o21ai_1 _26223_ (.B1(_07323_),
    .Y(_07324_),
    .A1(_09927_),
    .A2(net72));
 sg13g2_nand3_1 _26224_ (.B(_05484_),
    .C(_07311_),
    .A(_05436_),
    .Y(_07325_));
 sg13g2_a21oi_1 _26225_ (.A1(net71),
    .A2(_07325_),
    .Y(_07326_),
    .B1(net79));
 sg13g2_nor2_1 _26226_ (.A(_05583_),
    .B(_07326_),
    .Y(_07327_));
 sg13g2_a21oi_1 _26227_ (.A1(net73),
    .A2(_07324_),
    .Y(_02470_),
    .B1(_07327_));
 sg13g2_and2_1 _26228_ (.A(_07303_),
    .B(_07322_),
    .X(_07328_));
 sg13g2_buf_1 _26229_ (.A(_07328_),
    .X(_07329_));
 sg13g2_nand3_1 _26230_ (.B(_07286_),
    .C(_07329_),
    .A(_05673_),
    .Y(_07330_));
 sg13g2_o21ai_1 _26231_ (.B1(_07330_),
    .Y(_07331_),
    .A1(_09933_),
    .A2(net72));
 sg13g2_o21ai_1 _26232_ (.B1(net82),
    .Y(_07332_),
    .A1(net78),
    .A2(_07329_));
 sg13g2_inv_1 _26233_ (.Y(_07333_),
    .A(_05673_));
 sg13g2_a22oi_1 _26234_ (.Y(_02471_),
    .B1(_07332_),
    .B2(_07333_),
    .A2(_07331_),
    .A1(net73));
 sg13g2_nand4_1 _26235_ (.B(_05025_),
    .C(_07311_),
    .A(_05673_),
    .Y(_07334_),
    .D(_07322_));
 sg13g2_nand2b_1 _26236_ (.Y(_07335_),
    .B(net71),
    .A_N(_07334_));
 sg13g2_o21ai_1 _26237_ (.B1(_07335_),
    .Y(_07336_),
    .A1(_09940_),
    .A2(net72));
 sg13g2_nand3_1 _26238_ (.B(_07311_),
    .C(_07322_),
    .A(_05673_),
    .Y(_07337_));
 sg13g2_a21oi_1 _26239_ (.A1(net71),
    .A2(_07337_),
    .Y(_07338_),
    .B1(_09954_));
 sg13g2_nor2_1 _26240_ (.A(_05025_),
    .B(_07338_),
    .Y(_07339_));
 sg13g2_a21oi_1 _26241_ (.A1(net73),
    .A2(_07336_),
    .Y(_02472_),
    .B1(_07339_));
 sg13g2_and3_1 _26242_ (.X(_07340_),
    .A(_05673_),
    .B(_05025_),
    .C(_07322_));
 sg13g2_buf_1 _26243_ (.A(_07340_),
    .X(_07341_));
 sg13g2_nand2_1 _26244_ (.Y(_07342_),
    .A(_07303_),
    .B(_07341_));
 sg13g2_nor3_1 _26245_ (.A(_05692_),
    .B(net90),
    .C(_07342_),
    .Y(_07343_));
 sg13g2_a21oi_1 _26246_ (.A1(_10008_),
    .A2(net78),
    .Y(_07344_),
    .B1(_07343_));
 sg13g2_a21oi_1 _26247_ (.A1(_07288_),
    .A2(_07342_),
    .Y(_07345_),
    .B1(_09954_));
 sg13g2_nand2b_1 _26248_ (.Y(_07346_),
    .B(_05692_),
    .A_N(_07345_));
 sg13g2_o21ai_1 _26249_ (.B1(_07346_),
    .Y(_02473_),
    .A1(net79),
    .A2(_07344_));
 sg13g2_nand4_1 _26250_ (.B(_10040_),
    .C(_07309_),
    .A(_05692_),
    .Y(_07347_),
    .D(_07341_));
 sg13g2_nor3_1 _26251_ (.A(_05702_),
    .B(net90),
    .C(_07347_),
    .Y(_07348_));
 sg13g2_a21oi_1 _26252_ (.A1(_10013_),
    .A2(net90),
    .Y(_07349_),
    .B1(_07348_));
 sg13g2_a21oi_1 _26253_ (.A1(_07288_),
    .A2(_07347_),
    .Y(_07350_),
    .B1(_09954_));
 sg13g2_nand2b_1 _26254_ (.Y(_07351_),
    .B(_05702_),
    .A_N(_07350_));
 sg13g2_o21ai_1 _26255_ (.B1(_07351_),
    .Y(_02474_),
    .A1(net79),
    .A2(_07349_));
 sg13g2_nand2_1 _26256_ (.Y(_07352_),
    .A(_05692_),
    .B(_05702_));
 sg13g2_nand3_1 _26257_ (.B(_05025_),
    .C(_07329_),
    .A(_05673_),
    .Y(_07353_));
 sg13g2_buf_1 _26258_ (.A(_07353_),
    .X(_07354_));
 sg13g2_nor4_1 _26259_ (.A(_05109_),
    .B(net90),
    .C(_07352_),
    .D(_07354_),
    .Y(_07355_));
 sg13g2_a21oi_1 _26260_ (.A1(_10018_),
    .A2(net90),
    .Y(_07356_),
    .B1(_07355_));
 sg13g2_nor2_1 _26261_ (.A(_07352_),
    .B(_07354_),
    .Y(_07357_));
 sg13g2_nor2_1 _26262_ (.A(net124),
    .B(_07357_),
    .Y(_07358_));
 sg13g2_o21ai_1 _26263_ (.B1(_05109_),
    .Y(_07359_),
    .A1(net79),
    .A2(_07358_));
 sg13g2_o21ai_1 _26264_ (.B1(_07359_),
    .Y(_02475_),
    .A1(net79),
    .A2(_07356_));
 sg13g2_nand3_1 _26265_ (.B(_05702_),
    .C(_05109_),
    .A(_05692_),
    .Y(_07360_));
 sg13g2_or2_1 _26266_ (.X(_07361_),
    .B(_07360_),
    .A(_07334_));
 sg13g2_buf_1 _26267_ (.A(_07361_),
    .X(_07362_));
 sg13g2_nor3_1 _26268_ (.A(_05124_),
    .B(net90),
    .C(_07362_),
    .Y(_07363_));
 sg13g2_a21oi_1 _26269_ (.A1(_10025_),
    .A2(net90),
    .Y(_07364_),
    .B1(_07363_));
 sg13g2_nor2b_1 _26270_ (.A(net124),
    .B_N(_07362_),
    .Y(_07365_));
 sg13g2_o21ai_1 _26271_ (.B1(_05124_),
    .Y(_07366_),
    .A1(net79),
    .A2(_07365_));
 sg13g2_o21ai_1 _26272_ (.B1(_07366_),
    .Y(_02476_),
    .A1(_09955_),
    .A2(_07364_));
 sg13g2_inv_1 _26273_ (.Y(_07367_),
    .A(_05124_));
 sg13g2_nor2_1 _26274_ (.A(_07367_),
    .B(_07360_),
    .Y(_07368_));
 sg13g2_nor2b_1 _26275_ (.A(_07342_),
    .B_N(_07368_),
    .Y(_07369_));
 sg13g2_nand3_1 _26276_ (.B(_07286_),
    .C(_07369_),
    .A(_05150_),
    .Y(_07370_));
 sg13g2_o21ai_1 _26277_ (.B1(_07370_),
    .Y(_07371_),
    .A1(_10030_),
    .A2(_07287_));
 sg13g2_o21ai_1 _26278_ (.B1(net82),
    .Y(_07372_),
    .A1(net101),
    .A2(_07369_));
 sg13g2_inv_1 _26279_ (.Y(_07373_),
    .A(_05150_));
 sg13g2_a22oi_1 _26280_ (.Y(_02477_),
    .B1(_07372_),
    .B2(_07373_),
    .A2(_07371_),
    .A1(_07284_));
 sg13g2_and4_1 _26281_ (.A(_05150_),
    .B(_07311_),
    .C(_07341_),
    .D(_07368_),
    .X(_07374_));
 sg13g2_nand3_1 _26282_ (.B(_07286_),
    .C(_07374_),
    .A(_05183_),
    .Y(_07375_));
 sg13g2_o21ai_1 _26283_ (.B1(_07375_),
    .Y(_07376_),
    .A1(_10036_),
    .A2(net71));
 sg13g2_o21ai_1 _26284_ (.B1(net82),
    .Y(_07377_),
    .A1(_09966_),
    .A2(_07374_));
 sg13g2_inv_1 _26285_ (.Y(_07378_),
    .A(_05183_));
 sg13g2_a22oi_1 _26286_ (.Y(_02478_),
    .B1(_07377_),
    .B2(_07378_),
    .A2(_07376_),
    .A1(_07284_));
 sg13g2_nand2_1 _26287_ (.Y(_07379_),
    .A(_05150_),
    .B(_07368_));
 sg13g2_nor3_1 _26288_ (.A(_07378_),
    .B(_07354_),
    .C(_07379_),
    .Y(_07380_));
 sg13g2_o21ai_1 _26289_ (.B1(_07282_),
    .Y(_07381_),
    .A1(net124),
    .A2(_07380_));
 sg13g2_inv_1 _26290_ (.Y(_07382_),
    .A(_07380_));
 sg13g2_nor3_1 _26291_ (.A(_05216_),
    .B(net124),
    .C(_07382_),
    .Y(_07383_));
 sg13g2_a221oi_1 _26292_ (.B2(_05216_),
    .C1(_07383_),
    .B1(_07381_),
    .A1(_10043_),
    .Y(_07384_),
    .A2(_09966_));
 sg13g2_inv_1 _26293_ (.Y(_02479_),
    .A(_07384_));
 sg13g2_nand4_1 _26294_ (.B(_05150_),
    .C(_05183_),
    .A(_05124_),
    .Y(_07385_),
    .D(_05216_));
 sg13g2_nor3_1 _26295_ (.A(_05244_),
    .B(_07362_),
    .C(_07385_),
    .Y(_07386_));
 sg13g2_a22oi_1 _26296_ (.Y(_07387_),
    .B1(_07287_),
    .B2(_07386_),
    .A2(net124),
    .A1(_10048_));
 sg13g2_nor2_1 _26297_ (.A(_07362_),
    .B(_07385_),
    .Y(_07388_));
 sg13g2_o21ai_1 _26298_ (.B1(_07283_),
    .Y(_07389_),
    .A1(_09965_),
    .A2(_07388_));
 sg13g2_nand2_1 _26299_ (.Y(_07390_),
    .A(_05244_),
    .B(_07389_));
 sg13g2_o21ai_1 _26300_ (.B1(_07390_),
    .Y(_02480_),
    .A1(_09955_),
    .A2(_07387_));
 sg13g2_buf_1 _26301_ (.A(net779),
    .X(_07391_));
 sg13g2_nor2_1 _26302_ (.A(\cpu.r_clk_invert ),
    .B(net679),
    .Y(_07392_));
 sg13g2_a21oi_1 _26303_ (.A1(_09063_),
    .A2(_07391_),
    .Y(_02547_),
    .B1(_07392_));
 sg13g2_nand2b_1 _26304_ (.Y(_07393_),
    .B(net897),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26305_ (.A(_07393_),
    .X(_07394_));
 sg13g2_nor2b_1 _26306_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(_11873_),
    .Y(_07395_));
 sg13g2_nand4_1 _26307_ (.B(_02879_),
    .C(_12013_),
    .A(_09223_),
    .Y(_07396_),
    .D(net863));
 sg13g2_buf_2 _26308_ (.A(_07396_),
    .X(_07397_));
 sg13g2_nor2_1 _26309_ (.A(net488),
    .B(_07397_),
    .Y(_07398_));
 sg13g2_nor3_1 _26310_ (.A(_07394_),
    .B(_07395_),
    .C(_07398_),
    .Y(_00741_));
 sg13g2_nor2_1 _26311_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net411),
    .Y(_07399_));
 sg13g2_nor2_1 _26312_ (.A(net536),
    .B(_07397_),
    .Y(_07400_));
 sg13g2_nor3_1 _26313_ (.A(_07394_),
    .B(_07399_),
    .C(_07400_),
    .Y(_00742_));
 sg13g2_nor2_1 _26314_ (.A(\cpu.dcache.r_valid[2] ),
    .B(net472),
    .Y(_07401_));
 sg13g2_nor2_1 _26315_ (.A(net600),
    .B(_07397_),
    .Y(_07402_));
 sg13g2_nor3_1 _26316_ (.A(_07394_),
    .B(_07401_),
    .C(_07402_),
    .Y(_00743_));
 sg13g2_nor2_1 _26317_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net370),
    .Y(_07403_));
 sg13g2_nor2_1 _26318_ (.A(net482),
    .B(_07397_),
    .Y(_07404_));
 sg13g2_nor3_1 _26319_ (.A(_07394_),
    .B(_07403_),
    .C(_07404_),
    .Y(_00744_));
 sg13g2_a21oi_1 _26320_ (.A1(_12378_),
    .A2(_11782_),
    .Y(_07405_),
    .B1(\cpu.dcache.r_valid[4] ));
 sg13g2_nor2_1 _26321_ (.A(net599),
    .B(_07397_),
    .Y(_07406_));
 sg13g2_nor3_1 _26322_ (.A(_07394_),
    .B(_07405_),
    .C(_07406_),
    .Y(_00745_));
 sg13g2_nor2_1 _26323_ (.A(\cpu.dcache.r_valid[5] ),
    .B(_12492_),
    .Y(_07407_));
 sg13g2_nor2_1 _26324_ (.A(net534),
    .B(_07397_),
    .Y(_07408_));
 sg13g2_nor3_1 _26325_ (.A(_07394_),
    .B(_07407_),
    .C(_07408_),
    .Y(_00746_));
 sg13g2_nor2_1 _26326_ (.A(\cpu.dcache.r_valid[6] ),
    .B(net418),
    .Y(_07409_));
 sg13g2_nor2_1 _26327_ (.A(_12545_),
    .B(_07397_),
    .Y(_07410_));
 sg13g2_nor3_1 _26328_ (.A(_07394_),
    .B(_07409_),
    .C(_07410_),
    .Y(_00747_));
 sg13g2_nor2_1 _26329_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net367),
    .Y(_07411_));
 sg13g2_nor2_1 _26330_ (.A(net479),
    .B(_07397_),
    .Y(_07412_));
 sg13g2_nor3_1 _26331_ (.A(_07394_),
    .B(_07411_),
    .C(_07412_),
    .Y(_00748_));
 sg13g2_nor2_1 _26332_ (.A(net1011),
    .B(net1010),
    .Y(_07413_));
 sg13g2_nand3_1 _26333_ (.B(_07413_),
    .C(_04731_),
    .A(_10059_),
    .Y(_07414_));
 sg13g2_buf_1 _26334_ (.A(_07414_),
    .X(_07415_));
 sg13g2_nor2_1 _26335_ (.A(_03702_),
    .B(net572),
    .Y(_07416_));
 sg13g2_a21oi_1 _26336_ (.A1(_08735_),
    .A2(net572),
    .Y(_07417_),
    .B1(_07416_));
 sg13g2_nor3_1 _26337_ (.A(net311),
    .B(_09185_),
    .C(_07417_),
    .Y(_00797_));
 sg13g2_and4_1 _26338_ (.A(_03217_),
    .B(_10921_),
    .C(\cpu.dec.do_flush_all ),
    .D(net737),
    .X(_00930_));
 sg13g2_and4_1 _26339_ (.A(_03217_),
    .B(_10888_),
    .C(\cpu.dec.do_flush_all ),
    .D(_10723_),
    .X(_00948_));
 sg13g2_o21ai_1 _26340_ (.B1(net347),
    .Y(_07418_),
    .A1(net1027),
    .A2(_10181_));
 sg13g2_nand2_1 _26341_ (.Y(_07419_),
    .A(_06684_),
    .B(net1027));
 sg13g2_nor2_1 _26342_ (.A(_11345_),
    .B(_10376_),
    .Y(_07420_));
 sg13g2_nand4_1 _26343_ (.B(net737),
    .C(_10244_),
    .A(net719),
    .Y(_07421_),
    .D(_07420_));
 sg13g2_mux2_1 _26344_ (.A0(_10288_),
    .A1(_09073_),
    .S(_07421_),
    .X(_07422_));
 sg13g2_nand2_1 _26345_ (.Y(_07423_),
    .A(net572),
    .B(_07422_));
 sg13g2_o21ai_1 _26346_ (.B1(_07423_),
    .Y(_07424_),
    .A1(_03747_),
    .A2(net572));
 sg13g2_nand2_1 _26347_ (.Y(_07425_),
    .A(_09128_),
    .B(_07424_));
 sg13g2_a21oi_1 _26348_ (.A1(_07418_),
    .A2(_07419_),
    .Y(_00949_),
    .B1(_07425_));
 sg13g2_nand2_1 _26349_ (.Y(_07426_),
    .A(_08764_),
    .B(net737));
 sg13g2_nor2_1 _26350_ (.A(_00310_),
    .B(_07426_),
    .Y(_07427_));
 sg13g2_inv_1 _26351_ (.Y(_07428_),
    .A(_09650_));
 sg13g2_nor2_1 _26352_ (.A(net1031),
    .B(net1030),
    .Y(_07429_));
 sg13g2_a22oi_1 _26353_ (.Y(_07430_),
    .B1(_11782_),
    .B2(_07429_),
    .A2(_07428_),
    .A1(_09223_));
 sg13g2_nand3_1 _26354_ (.B(_11362_),
    .C(_07430_),
    .A(_11361_),
    .Y(_07431_));
 sg13g2_a21oi_1 _26355_ (.A1(_09021_),
    .A2(_07431_),
    .Y(_07432_),
    .B1(_09181_));
 sg13g2_o21ai_1 _26356_ (.B1(_07432_),
    .Y(_07433_),
    .A1(_09019_),
    .A2(_07427_));
 sg13g2_nor3_1 _26357_ (.A(_09019_),
    .B(_00298_),
    .C(_04790_),
    .Y(_07434_));
 sg13g2_o21ai_1 _26358_ (.B1(_07434_),
    .Y(_07435_),
    .A1(_11336_),
    .A2(_04768_));
 sg13g2_nor2b_1 _26359_ (.A(_07433_),
    .B_N(_07435_),
    .Y(_01068_));
 sg13g2_nand3b_1 _26360_ (.B(_07432_),
    .C(_07427_),
    .Y(_07436_),
    .A_N(_04790_));
 sg13g2_a22oi_1 _26361_ (.Y(_07437_),
    .B1(_07427_),
    .B2(net1033),
    .A2(_07432_),
    .A1(_08762_));
 sg13g2_o21ai_1 _26362_ (.B1(_07437_),
    .Y(_01069_),
    .A1(_04769_),
    .A2(_07436_));
 sg13g2_inv_1 _26363_ (.Y(_07438_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26364_ (.Y(_07439_),
    .B(net897),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26365_ (.A(_07439_),
    .X(_07440_));
 sg13g2_a21oi_1 _26366_ (.A1(_07438_),
    .A2(_06413_),
    .Y(_02424_),
    .B1(_07440_));
 sg13g2_nor2_1 _26367_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06324_),
    .Y(_07441_));
 sg13g2_nor2_1 _26368_ (.A(_07440_),
    .B(_07441_),
    .Y(_02425_));
 sg13g2_nor2_1 _26369_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06340_),
    .Y(_07442_));
 sg13g2_nor2_1 _26370_ (.A(_07440_),
    .B(_07442_),
    .Y(_02426_));
 sg13g2_inv_1 _26371_ (.Y(_07443_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26372_ (.A1(_07443_),
    .A2(net216),
    .Y(_02427_),
    .B1(_07440_));
 sg13g2_nor2_1 _26373_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06372_),
    .Y(_07444_));
 sg13g2_nor2_1 _26374_ (.A(_07440_),
    .B(_07444_),
    .Y(_02428_));
 sg13g2_inv_1 _26375_ (.Y(_07445_),
    .A(\cpu.icache.r_valid[5] ));
 sg13g2_a21oi_1 _26376_ (.A1(_07445_),
    .A2(_06385_),
    .Y(_02429_),
    .B1(_07440_));
 sg13g2_inv_1 _26377_ (.Y(_07446_),
    .A(\cpu.icache.r_valid[6] ));
 sg13g2_a21oi_1 _26378_ (.A1(_07446_),
    .A2(_06394_),
    .Y(_02430_),
    .B1(_07440_));
 sg13g2_nor2_1 _26379_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06408_),
    .Y(_07447_));
 sg13g2_nor2_1 _26380_ (.A(_07440_),
    .B(_07447_),
    .Y(_02431_));
 sg13g2_nand3_1 _26381_ (.B(_09957_),
    .C(net399),
    .A(_09915_),
    .Y(_07448_));
 sg13g2_and2_1 _26382_ (.A(net123),
    .B(net363),
    .X(_07449_));
 sg13g2_buf_1 _26383_ (.A(_07449_),
    .X(_07450_));
 sg13g2_a22oi_1 _26384_ (.Y(_07451_),
    .B1(_07450_),
    .B2(net964),
    .A2(_07448_),
    .A1(_09031_));
 sg13g2_nor2_1 _26385_ (.A(net617),
    .B(_07451_),
    .Y(_00317_));
 sg13g2_nor2_1 _26386_ (.A(_02879_),
    .B(net994),
    .Y(_07452_));
 sg13g2_nor2b_1 _26387_ (.A(_07452_),
    .B_N(_00315_),
    .Y(_00586_));
 sg13g2_a21oi_1 _26388_ (.A1(_06698_),
    .A2(_06701_),
    .Y(_00587_),
    .B1(_07452_));
 sg13g2_xnor2_1 _26389_ (.Y(_07453_),
    .A(_06705_),
    .B(_11780_));
 sg13g2_nor2_1 _26390_ (.A(_07452_),
    .B(_07453_),
    .Y(_00588_));
 sg13g2_nor2_1 _26391_ (.A(_09131_),
    .B(net572),
    .Y(_07454_));
 sg13g2_a21oi_1 _26392_ (.A1(net1053),
    .A2(net572),
    .Y(_07455_),
    .B1(_07454_));
 sg13g2_nor2_1 _26393_ (.A(_09187_),
    .B(_07455_),
    .Y(_00798_));
 sg13g2_nor2_1 _26394_ (.A(_10343_),
    .B(net1027),
    .Y(_07456_));
 sg13g2_nand3_1 _26395_ (.B(_07420_),
    .C(_07456_),
    .A(_10244_),
    .Y(_07457_));
 sg13g2_a21oi_1 _26396_ (.A1(net719),
    .A2(_07457_),
    .Y(_07458_),
    .B1(_09123_));
 sg13g2_nor2_1 _26397_ (.A(_03686_),
    .B(_07458_),
    .Y(_07459_));
 sg13g2_nor2_1 _26398_ (.A(_10343_),
    .B(_07459_),
    .Y(_07460_));
 sg13g2_a21oi_1 _26399_ (.A1(_03747_),
    .A2(_07459_),
    .Y(_07461_),
    .B1(_07460_));
 sg13g2_a22oi_1 _26400_ (.Y(_07462_),
    .B1(net737),
    .B2(net1110),
    .A2(net311),
    .A1(_06720_));
 sg13g2_or2_1 _26401_ (.X(_07463_),
    .B(_07462_),
    .A(_04125_));
 sg13g2_buf_1 _26402_ (.A(_07463_),
    .X(_07464_));
 sg13g2_mux2_1 _26403_ (.A0(net719),
    .A1(_07461_),
    .S(_07464_),
    .X(_07465_));
 sg13g2_nand2b_1 _26404_ (.Y(_00799_),
    .B(_06655_),
    .A_N(_07465_));
 sg13g2_mux2_1 _26405_ (.A0(net1037),
    .A1(_10416_),
    .S(net572),
    .X(_07466_));
 sg13g2_and2_1 _26406_ (.A(_11663_),
    .B(_07466_),
    .X(_00800_));
 sg13g2_nand2_1 _26407_ (.Y(_07467_),
    .A(_09021_),
    .B(_07431_));
 sg13g2_nor4_1 _26408_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11337_),
    .C(_03337_),
    .D(_07426_),
    .Y(_07468_));
 sg13g2_nor2_1 _26409_ (.A(_10068_),
    .B(_07468_),
    .Y(_07469_));
 sg13g2_nand2_1 _26410_ (.Y(_07470_),
    .A(net1110),
    .B(_11339_));
 sg13g2_a21oi_1 _26411_ (.A1(_07467_),
    .A2(_07469_),
    .Y(_07471_),
    .B1(_07470_));
 sg13g2_nor3_1 _26412_ (.A(_06720_),
    .B(_04992_),
    .C(_07471_),
    .Y(_07472_));
 sg13g2_nor2_1 _26413_ (.A(_06684_),
    .B(net98),
    .Y(_07473_));
 sg13g2_o21ai_1 _26414_ (.B1(_06655_),
    .Y(_00946_),
    .A1(_07472_),
    .A2(_07473_));
 sg13g2_nand2_1 _26415_ (.Y(_07474_),
    .A(_09223_),
    .B(net1027));
 sg13g2_nand3_1 _26416_ (.B(\cpu.dec.do_flush_write ),
    .C(_11342_),
    .A(net719),
    .Y(_07475_));
 sg13g2_buf_1 _26417_ (.A(_09183_),
    .X(_07476_));
 sg13g2_a21oi_1 _26418_ (.A1(_07474_),
    .A2(_07475_),
    .Y(_00947_),
    .B1(net571));
 sg13g2_nand2_1 _26419_ (.Y(_07477_),
    .A(\cpu.dec.io ),
    .B(_11342_));
 sg13g2_nand2_1 _26420_ (.Y(_07478_),
    .A(_02878_),
    .B(net1027));
 sg13g2_a21oi_1 _26421_ (.A1(_07477_),
    .A2(_07478_),
    .Y(_00950_),
    .B1(_07476_));
 sg13g2_nor2_1 _26422_ (.A(_09073_),
    .B(_07464_),
    .Y(_07479_));
 sg13g2_nand2_1 _26423_ (.Y(_07480_),
    .A(_10288_),
    .B(_07415_));
 sg13g2_o21ai_1 _26424_ (.B1(_07480_),
    .Y(_07481_),
    .A1(net608),
    .A2(net572));
 sg13g2_nor2b_1 _26425_ (.A(_07481_),
    .B_N(_07464_),
    .Y(_07482_));
 sg13g2_nor3_1 _26426_ (.A(_09185_),
    .B(_07479_),
    .C(_07482_),
    .Y(_00997_));
 sg13g2_a22oi_1 _26427_ (.Y(_07483_),
    .B1(_03444_),
    .B2(net1111),
    .A2(_11342_),
    .A1(_11337_));
 sg13g2_nor2_1 _26428_ (.A(_09187_),
    .B(_07483_),
    .Y(_00998_));
 sg13g2_nor2_2 _26429_ (.A(net841),
    .B(_05774_),
    .Y(_07484_));
 sg13g2_mux2_1 _26430_ (.A0(_10242_),
    .A1(_09094_),
    .S(_07484_),
    .X(_07485_));
 sg13g2_nand2_1 _26431_ (.Y(_07486_),
    .A(net347),
    .B(_07485_));
 sg13g2_a21oi_1 _26432_ (.A1(_11338_),
    .A2(_07486_),
    .Y(_01074_),
    .B1(_07476_));
 sg13g2_buf_1 _26433_ (.A(_09186_),
    .X(_07487_));
 sg13g2_nand2_1 _26434_ (.Y(_07488_),
    .A(_09119_),
    .B(_07484_));
 sg13g2_o21ai_1 _26435_ (.B1(_07488_),
    .Y(_07489_),
    .A1(_05835_),
    .A2(_07484_));
 sg13g2_nor2_1 _26436_ (.A(net674),
    .B(_08838_),
    .Y(_07490_));
 sg13g2_a21oi_1 _26437_ (.A1(net347),
    .A2(_07489_),
    .Y(_07491_),
    .B1(_07490_));
 sg13g2_nor2_1 _26438_ (.A(net570),
    .B(_07491_),
    .Y(_01075_));
 sg13g2_mux2_1 _26439_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_09943_),
    .S(_07484_),
    .X(_07492_));
 sg13g2_a21oi_1 _26440_ (.A1(_09023_),
    .A2(_07492_),
    .Y(_07493_),
    .B1(_10460_));
 sg13g2_nor2_1 _26441_ (.A(net570),
    .B(_07493_),
    .Y(_01076_));
 sg13g2_nand2_1 _26442_ (.Y(_07494_),
    .A(net1068),
    .B(_05868_));
 sg13g2_nor4_2 _26443_ (.A(net1090),
    .B(net942),
    .C(net939),
    .Y(_07495_),
    .D(_07494_));
 sg13g2_nor2b_1 _26444_ (.A(_00257_),
    .B_N(_05766_),
    .Y(_07496_));
 sg13g2_and2_1 _26445_ (.A(_05764_),
    .B(_07496_),
    .X(_07497_));
 sg13g2_buf_1 _26446_ (.A(_07497_),
    .X(_07498_));
 sg13g2_o21ai_1 _26447_ (.B1(_07498_),
    .Y(_07499_),
    .A1(_03747_),
    .A2(_00255_));
 sg13g2_or2_1 _26448_ (.X(_07500_),
    .B(_07499_),
    .A(_04501_));
 sg13g2_buf_1 _26449_ (.A(_07500_),
    .X(_07501_));
 sg13g2_buf_1 _26450_ (.A(_07501_),
    .X(_07502_));
 sg13g2_nand2_1 _26451_ (.Y(_07503_),
    .A(_03219_),
    .B(_10921_));
 sg13g2_a21oi_1 _26452_ (.A1(_07499_),
    .A2(_07503_),
    .Y(_07504_),
    .B1(net311));
 sg13g2_buf_2 _26453_ (.A(_07504_),
    .X(_07505_));
 sg13g2_o21ai_1 _26454_ (.B1(_07505_),
    .Y(_07506_),
    .A1(_07495_),
    .A2(_07502_));
 sg13g2_nor2_1 _26455_ (.A(_09952_),
    .B(_07501_),
    .Y(_07507_));
 sg13g2_buf_2 _26456_ (.A(_07507_),
    .X(_07508_));
 sg13g2_buf_1 _26457_ (.A(_07508_),
    .X(_07509_));
 sg13g2_a22oi_1 _26458_ (.Y(_07510_),
    .B1(net126),
    .B2(_07495_),
    .A2(_07506_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26459_ (.A(net570),
    .B(_07510_),
    .Y(_01077_));
 sg13g2_nor3_1 _26460_ (.A(net940),
    .B(_04798_),
    .C(net709),
    .Y(_07511_));
 sg13g2_buf_2 _26461_ (.A(_07511_),
    .X(_07512_));
 sg13g2_nor2_1 _26462_ (.A(_10614_),
    .B(_07494_),
    .Y(_07513_));
 sg13g2_and2_1 _26463_ (.A(net939),
    .B(_07494_),
    .X(_07514_));
 sg13g2_a21oi_1 _26464_ (.A1(net942),
    .A2(_07513_),
    .Y(_07515_),
    .B1(_07514_));
 sg13g2_nor2_1 _26465_ (.A(_05835_),
    .B(net942),
    .Y(_07516_));
 sg13g2_nand2_1 _26466_ (.Y(_07517_),
    .A(_07516_),
    .B(_07513_));
 sg13g2_o21ai_1 _26467_ (.B1(_07517_),
    .Y(_07518_),
    .A1(net938),
    .A2(_07515_));
 sg13g2_buf_2 _26468_ (.A(_07518_),
    .X(_07519_));
 sg13g2_nor2b_2 _26469_ (.A(net172),
    .B_N(_07519_),
    .Y(_07520_));
 sg13g2_buf_1 _26470_ (.A(net172),
    .X(_07521_));
 sg13g2_buf_1 _26471_ (.A(_07505_),
    .X(_07522_));
 sg13g2_o21ai_1 _26472_ (.B1(net171),
    .Y(_07523_),
    .A1(_05829_),
    .A2(net150));
 sg13g2_a22oi_1 _26473_ (.Y(_07524_),
    .B1(_07523_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07520_),
    .A1(_07512_));
 sg13g2_nor2_1 _26474_ (.A(net570),
    .B(_07524_),
    .Y(_01078_));
 sg13g2_o21ai_1 _26475_ (.B1(_07522_),
    .Y(_07525_),
    .A1(_05838_),
    .A2(_07521_));
 sg13g2_a22oi_1 _26476_ (.Y(_07526_),
    .B1(_07525_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07508_),
    .A1(_05838_));
 sg13g2_nor2_1 _26477_ (.A(net570),
    .B(_07526_),
    .Y(_01079_));
 sg13g2_nand2_1 _26478_ (.Y(_07527_),
    .A(net940),
    .B(net991));
 sg13g2_nor3_1 _26479_ (.A(net835),
    .B(net941),
    .C(_07527_),
    .Y(_07528_));
 sg13g2_buf_2 _26480_ (.A(_07528_),
    .X(_07529_));
 sg13g2_buf_1 _26481_ (.A(net172),
    .X(_07530_));
 sg13g2_nand2b_1 _26482_ (.Y(_07531_),
    .B(net940),
    .A_N(net941));
 sg13g2_o21ai_1 _26483_ (.B1(_05793_),
    .Y(_07532_),
    .A1(net835),
    .A2(_07531_));
 sg13g2_and2_1 _26484_ (.A(net1068),
    .B(_07532_),
    .X(_07533_));
 sg13g2_buf_1 _26485_ (.A(_07533_),
    .X(_07534_));
 sg13g2_and2_1 _26486_ (.A(_07519_),
    .B(_07534_),
    .X(_07535_));
 sg13g2_o21ai_1 _26487_ (.B1(net171),
    .Y(_07536_),
    .A1(net149),
    .A2(_07535_));
 sg13g2_a22oi_1 _26488_ (.Y(_07537_),
    .B1(_07536_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07529_),
    .A1(_07520_));
 sg13g2_nor2_1 _26489_ (.A(net570),
    .B(_07537_),
    .Y(_01080_));
 sg13g2_nor2_1 _26490_ (.A(_05792_),
    .B(_05781_),
    .Y(_07538_));
 sg13g2_and2_1 _26491_ (.A(_07519_),
    .B(_07538_),
    .X(_07539_));
 sg13g2_buf_1 _26492_ (.A(_07539_),
    .X(_07540_));
 sg13g2_o21ai_1 _26493_ (.B1(net171),
    .Y(_07541_),
    .A1(net149),
    .A2(_07540_));
 sg13g2_a22oi_1 _26494_ (.Y(_07542_),
    .B1(_07541_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07540_),
    .A1(net126));
 sg13g2_nor2_1 _26495_ (.A(net570),
    .B(_07542_),
    .Y(_01081_));
 sg13g2_nor2_1 _26496_ (.A(net709),
    .B(_07527_),
    .Y(_07543_));
 sg13g2_buf_2 _26497_ (.A(_07543_),
    .X(_07544_));
 sg13g2_nor2_1 _26498_ (.A(_05792_),
    .B(net709),
    .Y(_07545_));
 sg13g2_and2_1 _26499_ (.A(_07519_),
    .B(_07545_),
    .X(_07546_));
 sg13g2_o21ai_1 _26500_ (.B1(net171),
    .Y(_07547_),
    .A1(net149),
    .A2(_07546_));
 sg13g2_a22oi_1 _26501_ (.Y(_07548_),
    .B1(_07547_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07544_),
    .A1(_07520_));
 sg13g2_nor2_1 _26502_ (.A(net570),
    .B(_07548_),
    .Y(_01082_));
 sg13g2_and2_1 _26503_ (.A(_05808_),
    .B(_07519_),
    .X(_07549_));
 sg13g2_buf_1 _26504_ (.A(_07549_),
    .X(_07550_));
 sg13g2_o21ai_1 _26505_ (.B1(net171),
    .Y(_07551_),
    .A1(_07530_),
    .A2(_07550_));
 sg13g2_a22oi_1 _26506_ (.Y(_07552_),
    .B1(_07551_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07550_),
    .A1(net126));
 sg13g2_nor2_1 _26507_ (.A(_07487_),
    .B(_07552_),
    .Y(_01083_));
 sg13g2_a21oi_1 _26508_ (.A1(net1068),
    .A2(_05817_),
    .Y(_07553_),
    .B1(_04798_));
 sg13g2_and2_1 _26509_ (.A(_06062_),
    .B(_07553_),
    .X(_07554_));
 sg13g2_buf_2 _26510_ (.A(_07554_),
    .X(_07555_));
 sg13g2_nor2_1 _26511_ (.A(_05817_),
    .B(_05870_),
    .Y(_07556_));
 sg13g2_o21ai_1 _26512_ (.B1(net1068),
    .Y(_07557_),
    .A1(_05808_),
    .A2(_07556_));
 sg13g2_nor2b_1 _26513_ (.A(_07557_),
    .B_N(_07519_),
    .Y(_07558_));
 sg13g2_nand2_1 _26514_ (.Y(_07559_),
    .A(_03219_),
    .B(_10811_));
 sg13g2_a21oi_1 _26515_ (.A1(_07499_),
    .A2(_07559_),
    .Y(_07560_),
    .B1(net311));
 sg13g2_buf_2 _26516_ (.A(_07560_),
    .X(_07561_));
 sg13g2_buf_1 _26517_ (.A(_07561_),
    .X(_07562_));
 sg13g2_o21ai_1 _26518_ (.B1(net170),
    .Y(_07563_),
    .A1(net149),
    .A2(_07558_));
 sg13g2_a22oi_1 _26519_ (.Y(_07564_),
    .B1(_07563_),
    .B2(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A2(_07555_),
    .A1(_07520_));
 sg13g2_nor2_1 _26520_ (.A(_07487_),
    .B(_07564_),
    .Y(_01084_));
 sg13g2_buf_1 _26521_ (.A(_09186_),
    .X(_07565_));
 sg13g2_nor4_1 _26522_ (.A(net1090),
    .B(net942),
    .C(net939),
    .D(net1068),
    .Y(_07566_));
 sg13g2_nand3_1 _26523_ (.B(net939),
    .C(net1068),
    .A(net1090),
    .Y(_07567_));
 sg13g2_nand2b_1 _26524_ (.Y(_07568_),
    .B(_07567_),
    .A_N(_07566_));
 sg13g2_nand2b_1 _26525_ (.Y(_07569_),
    .B(net942),
    .A_N(net1068));
 sg13g2_a21oi_1 _26526_ (.A1(_05868_),
    .A2(_07569_),
    .Y(_07570_),
    .B1(net834));
 sg13g2_a22oi_1 _26527_ (.Y(_07571_),
    .B1(_07570_),
    .B2(net938),
    .A2(_07568_),
    .A1(_05868_));
 sg13g2_buf_2 _26528_ (.A(_07571_),
    .X(_07572_));
 sg13g2_nor2_1 _26529_ (.A(net940),
    .B(_05781_),
    .Y(_07573_));
 sg13g2_nor2b_1 _26530_ (.A(_07572_),
    .B_N(_07573_),
    .Y(_07574_));
 sg13g2_o21ai_1 _26531_ (.B1(net170),
    .Y(_07575_),
    .A1(net149),
    .A2(_07574_));
 sg13g2_a22oi_1 _26532_ (.Y(_07576_),
    .B1(_07575_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07574_),
    .A1(net126));
 sg13g2_nor2_1 _26533_ (.A(net569),
    .B(_07576_),
    .Y(_01085_));
 sg13g2_nor2_1 _26534_ (.A(net172),
    .B(_07572_),
    .Y(_07577_));
 sg13g2_o21ai_1 _26535_ (.B1(net170),
    .Y(_07578_),
    .A1(_05888_),
    .A2(net150));
 sg13g2_a22oi_1 _26536_ (.Y(_07579_),
    .B1(_07578_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07577_),
    .A1(_07512_));
 sg13g2_nor2_1 _26537_ (.A(net569),
    .B(_07579_),
    .Y(_01086_));
 sg13g2_o21ai_1 _26538_ (.B1(_07562_),
    .Y(_07580_),
    .A1(_05894_),
    .A2(net150));
 sg13g2_a22oi_1 _26539_ (.Y(_07581_),
    .B1(_07580_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07508_),
    .A1(_05894_));
 sg13g2_nor2_1 _26540_ (.A(_07565_),
    .B(_07581_),
    .Y(_01087_));
 sg13g2_nor2_1 _26541_ (.A(net939),
    .B(_05767_),
    .Y(_07582_));
 sg13g2_a22oi_1 _26542_ (.Y(_07583_),
    .B1(_07516_),
    .B2(_07582_),
    .A2(_05843_),
    .A1(_05767_));
 sg13g2_inv_1 _26543_ (.Y(_07584_),
    .A(_07583_));
 sg13g2_a22oi_1 _26544_ (.Y(_07585_),
    .B1(_07584_),
    .B2(_05868_),
    .A2(_07570_),
    .A1(_05835_));
 sg13g2_buf_2 _26545_ (.A(_07585_),
    .X(_07586_));
 sg13g2_nor2b_2 _26546_ (.A(_07586_),
    .B_N(_07573_),
    .Y(_07587_));
 sg13g2_o21ai_1 _26547_ (.B1(net171),
    .Y(_07588_),
    .A1(net149),
    .A2(_07587_));
 sg13g2_a22oi_1 _26548_ (.Y(_07589_),
    .B1(_07588_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07587_),
    .A1(net126));
 sg13g2_nor2_1 _26549_ (.A(net569),
    .B(_07589_),
    .Y(_01088_));
 sg13g2_nor2b_1 _26550_ (.A(_07572_),
    .B_N(_07534_),
    .Y(_07590_));
 sg13g2_o21ai_1 _26551_ (.B1(net170),
    .Y(_07591_),
    .A1(net149),
    .A2(_07590_));
 sg13g2_a22oi_1 _26552_ (.Y(_07592_),
    .B1(_07591_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07577_),
    .A1(_07529_));
 sg13g2_nor2_1 _26553_ (.A(net569),
    .B(_07592_),
    .Y(_01089_));
 sg13g2_nor2b_1 _26554_ (.A(_07572_),
    .B_N(_07538_),
    .Y(_07593_));
 sg13g2_o21ai_1 _26555_ (.B1(net170),
    .Y(_07594_),
    .A1(net149),
    .A2(_07593_));
 sg13g2_a22oi_1 _26556_ (.Y(_07595_),
    .B1(_07594_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07593_),
    .A1(net126));
 sg13g2_nor2_1 _26557_ (.A(net569),
    .B(_07595_),
    .Y(_01090_));
 sg13g2_nor2b_1 _26558_ (.A(_07572_),
    .B_N(_07545_),
    .Y(_07596_));
 sg13g2_o21ai_1 _26559_ (.B1(net170),
    .Y(_07597_),
    .A1(_07530_),
    .A2(_07596_));
 sg13g2_a22oi_1 _26560_ (.Y(_07598_),
    .B1(_07597_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07577_),
    .A1(_07544_));
 sg13g2_nor2_1 _26561_ (.A(net569),
    .B(_07598_),
    .Y(_01091_));
 sg13g2_nor2_2 _26562_ (.A(_05892_),
    .B(_05976_),
    .Y(_07599_));
 sg13g2_buf_1 _26563_ (.A(net172),
    .X(_07600_));
 sg13g2_o21ai_1 _26564_ (.B1(_07562_),
    .Y(_07601_),
    .A1(net148),
    .A2(_07599_));
 sg13g2_a22oi_1 _26565_ (.Y(_07602_),
    .B1(_07601_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07599_),
    .A1(net126));
 sg13g2_nor2_1 _26566_ (.A(_07565_),
    .B(_07602_),
    .Y(_01092_));
 sg13g2_nor2_1 _26567_ (.A(_07557_),
    .B(_07572_),
    .Y(_07603_));
 sg13g2_o21ai_1 _26568_ (.B1(net170),
    .Y(_07604_),
    .A1(net148),
    .A2(_07603_));
 sg13g2_a22oi_1 _26569_ (.Y(_07605_),
    .B1(_07604_),
    .B2(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07577_),
    .A1(_07555_));
 sg13g2_nor2_1 _26570_ (.A(net569),
    .B(_07605_),
    .Y(_01093_));
 sg13g2_nor2_1 _26571_ (.A(_05835_),
    .B(_07515_),
    .Y(_07606_));
 sg13g2_or2_1 _26572_ (.X(_07607_),
    .B(_07606_),
    .A(_07495_));
 sg13g2_buf_1 _26573_ (.A(_07607_),
    .X(_07608_));
 sg13g2_and2_1 _26574_ (.A(_07573_),
    .B(_07608_),
    .X(_07609_));
 sg13g2_buf_1 _26575_ (.A(_07609_),
    .X(_07610_));
 sg13g2_o21ai_1 _26576_ (.B1(net170),
    .Y(_07611_),
    .A1(net148),
    .A2(_07610_));
 sg13g2_a22oi_1 _26577_ (.Y(_07612_),
    .B1(_07611_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07610_),
    .A1(net126));
 sg13g2_nor2_1 _26578_ (.A(net569),
    .B(_07612_),
    .Y(_01094_));
 sg13g2_buf_1 _26579_ (.A(_09186_),
    .X(_07613_));
 sg13g2_nor2b_1 _26580_ (.A(net172),
    .B_N(_07608_),
    .Y(_07614_));
 sg13g2_o21ai_1 _26581_ (.B1(_07561_),
    .Y(_07615_),
    .A1(_05930_),
    .A2(net150));
 sg13g2_a22oi_1 _26582_ (.Y(_07616_),
    .B1(_07615_),
    .B2(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A2(_07614_),
    .A1(_07512_));
 sg13g2_nor2_1 _26583_ (.A(net568),
    .B(_07616_),
    .Y(_01095_));
 sg13g2_o21ai_1 _26584_ (.B1(_07561_),
    .Y(_07617_),
    .A1(_05938_),
    .A2(net150));
 sg13g2_a22oi_1 _26585_ (.Y(_07618_),
    .B1(_07617_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07508_),
    .A1(_05938_));
 sg13g2_nor2_1 _26586_ (.A(net568),
    .B(_07618_),
    .Y(_01096_));
 sg13g2_and2_1 _26587_ (.A(_07534_),
    .B(_07608_),
    .X(_07619_));
 sg13g2_o21ai_1 _26588_ (.B1(_07561_),
    .Y(_07620_),
    .A1(net148),
    .A2(_07619_));
 sg13g2_a22oi_1 _26589_ (.Y(_07621_),
    .B1(_07620_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07614_),
    .A1(_07529_));
 sg13g2_nor2_1 _26590_ (.A(net568),
    .B(_07621_),
    .Y(_01097_));
 sg13g2_and2_1 _26591_ (.A(_07538_),
    .B(_07608_),
    .X(_07622_));
 sg13g2_buf_1 _26592_ (.A(_07622_),
    .X(_07623_));
 sg13g2_o21ai_1 _26593_ (.B1(_07561_),
    .Y(_07624_),
    .A1(net148),
    .A2(_07623_));
 sg13g2_a22oi_1 _26594_ (.Y(_07625_),
    .B1(_07624_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07623_),
    .A1(_07509_));
 sg13g2_nor2_1 _26595_ (.A(net568),
    .B(_07625_),
    .Y(_01098_));
 sg13g2_nor3_1 _26596_ (.A(_05794_),
    .B(net709),
    .C(_07586_),
    .Y(_07626_));
 sg13g2_o21ai_1 _26597_ (.B1(_07505_),
    .Y(_07627_),
    .A1(net172),
    .A2(_07626_));
 sg13g2_and2_1 _26598_ (.A(_11807_),
    .B(_07626_),
    .X(_07628_));
 sg13g2_inv_1 _26599_ (.Y(_07629_),
    .A(net150));
 sg13g2_a22oi_1 _26600_ (.Y(_07630_),
    .B1(_07628_),
    .B2(_07629_),
    .A2(_07627_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26601_ (.A(net568),
    .B(_07630_),
    .Y(_01099_));
 sg13g2_and2_1 _26602_ (.A(_07545_),
    .B(_07608_),
    .X(_07631_));
 sg13g2_o21ai_1 _26603_ (.B1(_07561_),
    .Y(_07632_),
    .A1(net148),
    .A2(_07631_));
 sg13g2_a22oi_1 _26604_ (.Y(_07633_),
    .B1(_07632_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07614_),
    .A1(_07544_));
 sg13g2_nor2_1 _26605_ (.A(net568),
    .B(_07633_),
    .Y(_01100_));
 sg13g2_and2_1 _26606_ (.A(_05808_),
    .B(_07608_),
    .X(_07634_));
 sg13g2_buf_1 _26607_ (.A(_07634_),
    .X(_07635_));
 sg13g2_o21ai_1 _26608_ (.B1(_07561_),
    .Y(_07636_),
    .A1(net148),
    .A2(_07635_));
 sg13g2_a22oi_1 _26609_ (.Y(_07637_),
    .B1(_07636_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07635_),
    .A1(_07509_));
 sg13g2_nor2_1 _26610_ (.A(net568),
    .B(_07637_),
    .Y(_01101_));
 sg13g2_nor2_2 _26611_ (.A(_05793_),
    .B(_07586_),
    .Y(_07638_));
 sg13g2_o21ai_1 _26612_ (.B1(net171),
    .Y(_07639_),
    .A1(net148),
    .A2(_07638_));
 sg13g2_a22oi_1 _26613_ (.Y(_07640_),
    .B1(_07639_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07638_),
    .A1(_07508_));
 sg13g2_nor2_1 _26614_ (.A(_07613_),
    .B(_07640_),
    .Y(_01102_));
 sg13g2_nor2_1 _26615_ (.A(_07502_),
    .B(_07586_),
    .Y(_07641_));
 sg13g2_nor2b_1 _26616_ (.A(_07586_),
    .B_N(_07534_),
    .Y(_07642_));
 sg13g2_o21ai_1 _26617_ (.B1(net171),
    .Y(_07643_),
    .A1(_07600_),
    .A2(_07642_));
 sg13g2_a22oi_1 _26618_ (.Y(_07644_),
    .B1(_07643_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07641_),
    .A1(_07529_));
 sg13g2_nor2_1 _26619_ (.A(net568),
    .B(_07644_),
    .Y(_01103_));
 sg13g2_o21ai_1 _26620_ (.B1(_07522_),
    .Y(_07645_),
    .A1(_05971_),
    .A2(_07521_));
 sg13g2_a22oi_1 _26621_ (.Y(_07646_),
    .B1(_07645_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07508_),
    .A1(_05971_));
 sg13g2_nor2_1 _26622_ (.A(_07613_),
    .B(_07646_),
    .Y(_01104_));
 sg13g2_buf_1 _26623_ (.A(_09186_),
    .X(_07647_));
 sg13g2_o21ai_1 _26624_ (.B1(_07505_),
    .Y(_07648_),
    .A1(_05977_),
    .A2(net150));
 sg13g2_a22oi_1 _26625_ (.Y(_07649_),
    .B1(_07648_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07641_),
    .A1(_07544_));
 sg13g2_nor2_1 _26626_ (.A(net567),
    .B(_07649_),
    .Y(_01105_));
 sg13g2_o21ai_1 _26627_ (.B1(_07505_),
    .Y(_07650_),
    .A1(_05982_),
    .A2(net150));
 sg13g2_a22oi_1 _26628_ (.Y(_07651_),
    .B1(_07650_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07508_),
    .A1(_05982_));
 sg13g2_nor2_1 _26629_ (.A(net567),
    .B(_07651_),
    .Y(_01106_));
 sg13g2_nor2_1 _26630_ (.A(_07557_),
    .B(_07586_),
    .Y(_07652_));
 sg13g2_o21ai_1 _26631_ (.B1(_07505_),
    .Y(_07653_),
    .A1(_07600_),
    .A2(_07652_));
 sg13g2_a22oi_1 _26632_ (.Y(_07654_),
    .B1(_07653_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07641_),
    .A1(_07555_));
 sg13g2_nor2_1 _26633_ (.A(_07647_),
    .B(_07654_),
    .Y(_01107_));
 sg13g2_and2_1 _26634_ (.A(_07519_),
    .B(_07573_),
    .X(_07655_));
 sg13g2_buf_1 _26635_ (.A(_07655_),
    .X(_07656_));
 sg13g2_o21ai_1 _26636_ (.B1(_07505_),
    .Y(_07657_),
    .A1(net172),
    .A2(_07656_));
 sg13g2_a22oi_1 _26637_ (.Y(_07658_),
    .B1(_07657_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07656_),
    .A1(_07508_));
 sg13g2_nor2_1 _26638_ (.A(_07647_),
    .B(_07658_),
    .Y(_01108_));
 sg13g2_nand2_1 _26639_ (.Y(_07659_),
    .A(net1032),
    .B(_00255_));
 sg13g2_nand3_1 _26640_ (.B(_07498_),
    .C(_07659_),
    .A(net379),
    .Y(_07660_));
 sg13g2_buf_1 _26641_ (.A(_07660_),
    .X(_07661_));
 sg13g2_buf_1 _26642_ (.A(_07661_),
    .X(_07662_));
 sg13g2_a22oi_1 _26643_ (.Y(_07663_),
    .B1(_05762_),
    .B2(_03219_),
    .A2(_00255_),
    .A1(_09098_));
 sg13g2_a22oi_1 _26644_ (.Y(_07664_),
    .B1(_07496_),
    .B2(_07663_),
    .A2(_10888_),
    .A1(_03219_));
 sg13g2_nor2_1 _26645_ (.A(_04501_),
    .B(_07664_),
    .Y(_07665_));
 sg13g2_buf_2 _26646_ (.A(_07665_),
    .X(_07666_));
 sg13g2_o21ai_1 _26647_ (.B1(_07666_),
    .Y(_07667_),
    .A1(_07495_),
    .A2(_07662_));
 sg13g2_nor2_1 _26648_ (.A(_09952_),
    .B(_07661_),
    .Y(_07668_));
 sg13g2_buf_2 _26649_ (.A(_07668_),
    .X(_07669_));
 sg13g2_buf_1 _26650_ (.A(_07669_),
    .X(_07670_));
 sg13g2_a22oi_1 _26651_ (.Y(_07671_),
    .B1(_07670_),
    .B2(_07495_),
    .A2(_07667_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26652_ (.A(net567),
    .B(_07671_),
    .Y(_01109_));
 sg13g2_nor2b_1 _26653_ (.A(net214),
    .B_N(_07519_),
    .Y(_07672_));
 sg13g2_buf_1 _26654_ (.A(net214),
    .X(_07673_));
 sg13g2_buf_1 _26655_ (.A(_07666_),
    .X(_07674_));
 sg13g2_o21ai_1 _26656_ (.B1(net168),
    .Y(_07675_),
    .A1(_05829_),
    .A2(net194));
 sg13g2_a22oi_1 _26657_ (.Y(_07676_),
    .B1(_07675_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07672_),
    .A1(_07512_));
 sg13g2_nor2_1 _26658_ (.A(net567),
    .B(_07676_),
    .Y(_01110_));
 sg13g2_o21ai_1 _26659_ (.B1(net168),
    .Y(_07677_),
    .A1(_05838_),
    .A2(_07673_));
 sg13g2_a22oi_1 _26660_ (.Y(_07678_),
    .B1(_07677_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(_07670_),
    .A1(_05838_));
 sg13g2_nor2_1 _26661_ (.A(net567),
    .B(_07678_),
    .Y(_01111_));
 sg13g2_o21ai_1 _26662_ (.B1(net168),
    .Y(_07679_),
    .A1(_07535_),
    .A2(net194));
 sg13g2_a22oi_1 _26663_ (.Y(_07680_),
    .B1(_07679_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07672_),
    .A1(_07529_));
 sg13g2_nor2_1 _26664_ (.A(net567),
    .B(_07680_),
    .Y(_01112_));
 sg13g2_o21ai_1 _26665_ (.B1(net168),
    .Y(_07681_),
    .A1(_07540_),
    .A2(net194));
 sg13g2_a22oi_1 _26666_ (.Y(_07682_),
    .B1(_07681_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(net169),
    .A1(_07540_));
 sg13g2_nor2_1 _26667_ (.A(net567),
    .B(_07682_),
    .Y(_01113_));
 sg13g2_o21ai_1 _26668_ (.B1(net168),
    .Y(_07683_),
    .A1(_07546_),
    .A2(net194));
 sg13g2_a22oi_1 _26669_ (.Y(_07684_),
    .B1(_07683_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07672_),
    .A1(_07544_));
 sg13g2_nor2_1 _26670_ (.A(net567),
    .B(_07684_),
    .Y(_01114_));
 sg13g2_buf_1 _26671_ (.A(_09186_),
    .X(_07685_));
 sg13g2_o21ai_1 _26672_ (.B1(net168),
    .Y(_07686_),
    .A1(_07550_),
    .A2(net194));
 sg13g2_a22oi_1 _26673_ (.Y(_07687_),
    .B1(_07686_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(net169),
    .A1(_07550_));
 sg13g2_nor2_1 _26674_ (.A(net566),
    .B(_07687_),
    .Y(_01115_));
 sg13g2_nand2_1 _26675_ (.Y(_07688_),
    .A(_07498_),
    .B(_07659_));
 sg13g2_nand2_1 _26676_ (.Y(_07689_),
    .A(_03219_),
    .B(_10852_));
 sg13g2_a21oi_1 _26677_ (.A1(_07688_),
    .A2(_07689_),
    .Y(_07690_),
    .B1(net311));
 sg13g2_buf_2 _26678_ (.A(_07690_),
    .X(_07691_));
 sg13g2_buf_1 _26679_ (.A(_07691_),
    .X(_07692_));
 sg13g2_o21ai_1 _26680_ (.B1(net167),
    .Y(_07693_),
    .A1(_07558_),
    .A2(net194));
 sg13g2_a22oi_1 _26681_ (.Y(_07694_),
    .B1(_07693_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07672_),
    .A1(_07555_));
 sg13g2_nor2_1 _26682_ (.A(net566),
    .B(_07694_),
    .Y(_01116_));
 sg13g2_o21ai_1 _26683_ (.B1(net167),
    .Y(_07695_),
    .A1(_07574_),
    .A2(net194));
 sg13g2_a22oi_1 _26684_ (.Y(_07696_),
    .B1(_07695_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net169),
    .A1(_07574_));
 sg13g2_nor2_1 _26685_ (.A(_07685_),
    .B(_07696_),
    .Y(_01117_));
 sg13g2_nor2_1 _26686_ (.A(_07572_),
    .B(net214),
    .Y(_07697_));
 sg13g2_o21ai_1 _26687_ (.B1(net167),
    .Y(_07698_),
    .A1(_05888_),
    .A2(net194));
 sg13g2_a22oi_1 _26688_ (.Y(_07699_),
    .B1(_07698_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07697_),
    .A1(_07512_));
 sg13g2_nor2_1 _26689_ (.A(net566),
    .B(_07699_),
    .Y(_01118_));
 sg13g2_buf_1 _26690_ (.A(net214),
    .X(_07700_));
 sg13g2_o21ai_1 _26691_ (.B1(net167),
    .Y(_07701_),
    .A1(_05894_),
    .A2(net193));
 sg13g2_a22oi_1 _26692_ (.Y(_07702_),
    .B1(_07701_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net169),
    .A1(_05894_));
 sg13g2_nor2_1 _26693_ (.A(net566),
    .B(_07702_),
    .Y(_01119_));
 sg13g2_o21ai_1 _26694_ (.B1(net168),
    .Y(_07703_),
    .A1(_07587_),
    .A2(net193));
 sg13g2_a22oi_1 _26695_ (.Y(_07704_),
    .B1(_07703_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net169),
    .A1(_07587_));
 sg13g2_nor2_1 _26696_ (.A(net566),
    .B(_07704_),
    .Y(_01120_));
 sg13g2_o21ai_1 _26697_ (.B1(net167),
    .Y(_07705_),
    .A1(_07590_),
    .A2(net193));
 sg13g2_a22oi_1 _26698_ (.Y(_07706_),
    .B1(_07705_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07697_),
    .A1(_07529_));
 sg13g2_nor2_1 _26699_ (.A(net566),
    .B(_07706_),
    .Y(_01121_));
 sg13g2_o21ai_1 _26700_ (.B1(_07692_),
    .Y(_07707_),
    .A1(_07593_),
    .A2(net193));
 sg13g2_a22oi_1 _26701_ (.Y(_07708_),
    .B1(_07707_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net169),
    .A1(_07593_));
 sg13g2_nor2_1 _26702_ (.A(_07685_),
    .B(_07708_),
    .Y(_01122_));
 sg13g2_o21ai_1 _26703_ (.B1(_07692_),
    .Y(_07709_),
    .A1(_07596_),
    .A2(net193));
 sg13g2_a22oi_1 _26704_ (.Y(_07710_),
    .B1(_07709_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07697_),
    .A1(_07544_));
 sg13g2_nor2_1 _26705_ (.A(net566),
    .B(_07710_),
    .Y(_01123_));
 sg13g2_o21ai_1 _26706_ (.B1(net167),
    .Y(_07711_),
    .A1(_07599_),
    .A2(net193));
 sg13g2_a22oi_1 _26707_ (.Y(_07712_),
    .B1(_07711_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(net169),
    .A1(_07599_));
 sg13g2_nor2_1 _26708_ (.A(net566),
    .B(_07712_),
    .Y(_01124_));
 sg13g2_buf_1 _26709_ (.A(_09186_),
    .X(_07713_));
 sg13g2_o21ai_1 _26710_ (.B1(net167),
    .Y(_07714_),
    .A1(_07603_),
    .A2(net193));
 sg13g2_a22oi_1 _26711_ (.Y(_07715_),
    .B1(_07714_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07697_),
    .A1(_07555_));
 sg13g2_nor2_1 _26712_ (.A(net565),
    .B(_07715_),
    .Y(_01125_));
 sg13g2_o21ai_1 _26713_ (.B1(net167),
    .Y(_07716_),
    .A1(_07610_),
    .A2(net193));
 sg13g2_a22oi_1 _26714_ (.Y(_07717_),
    .B1(_07716_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(net169),
    .A1(_07610_));
 sg13g2_nor2_1 _26715_ (.A(net565),
    .B(_07717_),
    .Y(_01126_));
 sg13g2_nor2b_1 _26716_ (.A(net214),
    .B_N(_07608_),
    .Y(_07718_));
 sg13g2_o21ai_1 _26717_ (.B1(_07691_),
    .Y(_07719_),
    .A1(_05930_),
    .A2(_07700_));
 sg13g2_a22oi_1 _26718_ (.Y(_07720_),
    .B1(_07719_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07718_),
    .A1(_07512_));
 sg13g2_nor2_1 _26719_ (.A(net565),
    .B(_07720_),
    .Y(_01127_));
 sg13g2_o21ai_1 _26720_ (.B1(_07691_),
    .Y(_07721_),
    .A1(_05938_),
    .A2(_07700_));
 sg13g2_a22oi_1 _26721_ (.Y(_07722_),
    .B1(_07721_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07669_),
    .A1(_05938_));
 sg13g2_nor2_1 _26722_ (.A(net565),
    .B(_07722_),
    .Y(_01128_));
 sg13g2_buf_1 _26723_ (.A(net214),
    .X(_07723_));
 sg13g2_o21ai_1 _26724_ (.B1(_07691_),
    .Y(_07724_),
    .A1(_07619_),
    .A2(net192));
 sg13g2_a22oi_1 _26725_ (.Y(_07725_),
    .B1(_07724_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07718_),
    .A1(_07529_));
 sg13g2_nor2_1 _26726_ (.A(net565),
    .B(_07725_),
    .Y(_01129_));
 sg13g2_o21ai_1 _26727_ (.B1(_07691_),
    .Y(_07726_),
    .A1(_07623_),
    .A2(net192));
 sg13g2_a22oi_1 _26728_ (.Y(_07727_),
    .B1(_07726_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07669_),
    .A1(_07623_));
 sg13g2_nor2_1 _26729_ (.A(net565),
    .B(_07727_),
    .Y(_01130_));
 sg13g2_inv_1 _26730_ (.Y(_07728_),
    .A(_07673_));
 sg13g2_o21ai_1 _26731_ (.B1(_07674_),
    .Y(_07729_),
    .A1(_07626_),
    .A2(net192));
 sg13g2_a22oi_1 _26732_ (.Y(_07730_),
    .B1(_07729_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07728_),
    .A1(_07628_));
 sg13g2_nor2_1 _26733_ (.A(_07713_),
    .B(_07730_),
    .Y(_01131_));
 sg13g2_o21ai_1 _26734_ (.B1(_07691_),
    .Y(_07731_),
    .A1(_07631_),
    .A2(net192));
 sg13g2_a22oi_1 _26735_ (.Y(_07732_),
    .B1(_07731_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07718_),
    .A1(_07544_));
 sg13g2_nor2_1 _26736_ (.A(net565),
    .B(_07732_),
    .Y(_01132_));
 sg13g2_o21ai_1 _26737_ (.B1(_07691_),
    .Y(_07733_),
    .A1(_07635_),
    .A2(net192));
 sg13g2_a22oi_1 _26738_ (.Y(_07734_),
    .B1(_07733_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07669_),
    .A1(_07635_));
 sg13g2_nor2_1 _26739_ (.A(net565),
    .B(_07734_),
    .Y(_01133_));
 sg13g2_o21ai_1 _26740_ (.B1(_07674_),
    .Y(_07735_),
    .A1(_07638_),
    .A2(_07723_));
 sg13g2_a22oi_1 _26741_ (.Y(_07736_),
    .B1(_07735_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07669_),
    .A1(_07638_));
 sg13g2_nor2_1 _26742_ (.A(_07713_),
    .B(_07736_),
    .Y(_01134_));
 sg13g2_buf_1 _26743_ (.A(_09183_),
    .X(_07737_));
 sg13g2_nor2_1 _26744_ (.A(_07586_),
    .B(net214),
    .Y(_07738_));
 sg13g2_o21ai_1 _26745_ (.B1(net168),
    .Y(_07739_),
    .A1(_07642_),
    .A2(net192));
 sg13g2_a22oi_1 _26746_ (.Y(_07740_),
    .B1(_07739_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07738_),
    .A1(_07529_));
 sg13g2_nor2_1 _26747_ (.A(net564),
    .B(_07740_),
    .Y(_01135_));
 sg13g2_o21ai_1 _26748_ (.B1(_07666_),
    .Y(_07741_),
    .A1(_05971_),
    .A2(net192));
 sg13g2_a22oi_1 _26749_ (.Y(_07742_),
    .B1(_07741_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07669_),
    .A1(_05971_));
 sg13g2_nor2_1 _26750_ (.A(net564),
    .B(_07742_),
    .Y(_01136_));
 sg13g2_o21ai_1 _26751_ (.B1(_07666_),
    .Y(_07743_),
    .A1(_05977_),
    .A2(net192));
 sg13g2_a22oi_1 _26752_ (.Y(_07744_),
    .B1(_07743_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07738_),
    .A1(_07544_));
 sg13g2_nor2_1 _26753_ (.A(net564),
    .B(_07744_),
    .Y(_01137_));
 sg13g2_o21ai_1 _26754_ (.B1(_07666_),
    .Y(_07745_),
    .A1(_05982_),
    .A2(_07723_));
 sg13g2_a22oi_1 _26755_ (.Y(_07746_),
    .B1(_07745_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07669_),
    .A1(_05982_));
 sg13g2_nor2_1 _26756_ (.A(net564),
    .B(_07746_),
    .Y(_01138_));
 sg13g2_o21ai_1 _26757_ (.B1(_07666_),
    .Y(_07747_),
    .A1(_07652_),
    .A2(_07662_));
 sg13g2_a22oi_1 _26758_ (.Y(_07748_),
    .B1(_07747_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07738_),
    .A1(_07555_));
 sg13g2_nor2_1 _26759_ (.A(_07737_),
    .B(_07748_),
    .Y(_01139_));
 sg13g2_o21ai_1 _26760_ (.B1(_07666_),
    .Y(_07749_),
    .A1(_07656_),
    .A2(net214));
 sg13g2_a22oi_1 _26761_ (.Y(_07750_),
    .B1(_07749_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07669_),
    .A1(_07656_));
 sg13g2_nor2_1 _26762_ (.A(_07737_),
    .B(_07750_),
    .Y(_01140_));
 sg13g2_inv_1 _26763_ (.Y(_07751_),
    .A(_04923_));
 sg13g2_nor2_1 _26764_ (.A(_07751_),
    .B(_06236_),
    .Y(_07752_));
 sg13g2_buf_2 _26765_ (.A(_07752_),
    .X(_07753_));
 sg13g2_nand2_1 _26766_ (.Y(_07754_),
    .A(net959),
    .B(_07753_));
 sg13g2_or2_1 _26767_ (.X(_07755_),
    .B(_06236_),
    .A(_07751_));
 sg13g2_buf_2 _26768_ (.A(_07755_),
    .X(_07756_));
 sg13g2_nand2_1 _26769_ (.Y(_07757_),
    .A(_09050_),
    .B(_07756_));
 sg13g2_a21oi_1 _26770_ (.A1(_07754_),
    .A2(_07757_),
    .Y(_01941_),
    .B1(net571));
 sg13g2_nand2_1 _26771_ (.Y(_07758_),
    .A(net954),
    .B(_07753_));
 sg13g2_nand2_1 _26772_ (.Y(_07759_),
    .A(_09042_),
    .B(_07756_));
 sg13g2_a21oi_1 _26773_ (.A1(_07758_),
    .A2(_07759_),
    .Y(_01942_),
    .B1(net571));
 sg13g2_nand2_1 _26774_ (.Y(_07760_),
    .A(net855),
    .B(_07753_));
 sg13g2_nand2_1 _26775_ (.Y(_07761_),
    .A(_09044_),
    .B(_07756_));
 sg13g2_a21oi_1 _26776_ (.A1(_07760_),
    .A2(_07761_),
    .Y(_01943_),
    .B1(net571));
 sg13g2_nand2_1 _26777_ (.Y(_07762_),
    .A(net1017),
    .B(_07753_));
 sg13g2_nand2_1 _26778_ (.Y(_07763_),
    .A(_09054_),
    .B(_07756_));
 sg13g2_a21oi_1 _26779_ (.A1(_07762_),
    .A2(_07763_),
    .Y(_01944_),
    .B1(net571));
 sg13g2_nand2_1 _26780_ (.Y(_07764_),
    .A(net1016),
    .B(_07753_));
 sg13g2_nand2_1 _26781_ (.Y(_07765_),
    .A(\cpu.gpio.r_enable_in[4] ),
    .B(_07756_));
 sg13g2_a21oi_1 _26782_ (.A1(_07764_),
    .A2(_07765_),
    .Y(_01945_),
    .B1(net571));
 sg13g2_nand2_1 _26783_ (.Y(_07766_),
    .A(net1015),
    .B(_07753_));
 sg13g2_nand2_1 _26784_ (.Y(_07767_),
    .A(\cpu.gpio.r_enable_in[5] ),
    .B(_07756_));
 sg13g2_a21oi_1 _26785_ (.A1(_07766_),
    .A2(_07767_),
    .Y(_01946_),
    .B1(net571));
 sg13g2_nand2_1 _26786_ (.Y(_07768_),
    .A(net1014),
    .B(_07753_));
 sg13g2_nand2_1 _26787_ (.Y(_07769_),
    .A(\cpu.gpio.r_enable_in[6] ),
    .B(_07756_));
 sg13g2_a21oi_1 _26788_ (.A1(_07768_),
    .A2(_07769_),
    .Y(_01947_),
    .B1(net571));
 sg13g2_nand2_1 _26789_ (.Y(_07770_),
    .A(net1012),
    .B(_07753_));
 sg13g2_nand2_1 _26790_ (.Y(_07771_),
    .A(\cpu.gpio.r_enable_in[7] ),
    .B(_07756_));
 sg13g2_buf_1 _26791_ (.A(_09183_),
    .X(_07772_));
 sg13g2_a21oi_1 _26792_ (.A1(_07770_),
    .A2(_07771_),
    .Y(_01948_),
    .B1(net563));
 sg13g2_buf_1 _26793_ (.A(_06236_),
    .X(_07773_));
 sg13g2_nor2_1 _26794_ (.A(net310),
    .B(net81),
    .Y(_07774_));
 sg13g2_nand2_1 _26795_ (.Y(_07775_),
    .A(_09922_),
    .B(_07774_));
 sg13g2_o21ai_1 _26796_ (.B1(\cpu.gpio.r_enable_io[4] ),
    .Y(_07776_),
    .A1(net310),
    .A2(net81));
 sg13g2_a21oi_1 _26797_ (.A1(_07775_),
    .A2(_07776_),
    .Y(_01949_),
    .B1(net563));
 sg13g2_nand2_1 _26798_ (.Y(_07777_),
    .A(net1015),
    .B(_07774_));
 sg13g2_o21ai_1 _26799_ (.B1(_09056_),
    .Y(_07778_),
    .A1(net310),
    .A2(net81));
 sg13g2_a21oi_1 _26800_ (.A1(_07777_),
    .A2(_07778_),
    .Y(_01950_),
    .B1(net563));
 sg13g2_nand2_1 _26801_ (.Y(_07779_),
    .A(net1014),
    .B(_07774_));
 sg13g2_o21ai_1 _26802_ (.B1(\cpu.gpio.r_enable_io[6] ),
    .Y(_07780_),
    .A1(_05307_),
    .A2(net81));
 sg13g2_a21oi_1 _26803_ (.A1(_07779_),
    .A2(_07780_),
    .Y(_01951_),
    .B1(net563));
 sg13g2_nand2_1 _26804_ (.Y(_07781_),
    .A(net1012),
    .B(_07774_));
 sg13g2_o21ai_1 _26805_ (.B1(\cpu.gpio.r_enable_io[7] ),
    .Y(_07782_),
    .A1(_05307_),
    .A2(net81));
 sg13g2_a21oi_1 _26806_ (.A1(_07781_),
    .A2(_07782_),
    .Y(_01952_),
    .B1(_07772_));
 sg13g2_nor4_1 _26807_ (.A(net609),
    .B(_04907_),
    .C(net597),
    .D(_06236_),
    .Y(_07783_));
 sg13g2_buf_2 _26808_ (.A(_07783_),
    .X(_07784_));
 sg13g2_nand2_1 _26809_ (.Y(_07785_),
    .A(_09922_),
    .B(_07784_));
 sg13g2_nand2b_1 _26810_ (.Y(_07786_),
    .B(net7),
    .A_N(_07784_));
 sg13g2_a21oi_1 _26811_ (.A1(_07785_),
    .A2(_07786_),
    .Y(_01953_),
    .B1(net563));
 sg13g2_nand2_1 _26812_ (.Y(_07787_),
    .A(net1015),
    .B(_07784_));
 sg13g2_nand2b_1 _26813_ (.Y(_07788_),
    .B(net8),
    .A_N(_07784_));
 sg13g2_a21oi_1 _26814_ (.A1(_07787_),
    .A2(_07788_),
    .Y(_01954_),
    .B1(net563));
 sg13g2_nand2_1 _26815_ (.Y(_07789_),
    .A(net1014),
    .B(_07784_));
 sg13g2_nand2b_1 _26816_ (.Y(_07790_),
    .B(net9),
    .A_N(_07784_));
 sg13g2_a21oi_1 _26817_ (.A1(_07789_),
    .A2(_07790_),
    .Y(_01955_),
    .B1(net563));
 sg13g2_nand2_1 _26818_ (.Y(_07791_),
    .A(net1012),
    .B(_07784_));
 sg13g2_nand2b_1 _26819_ (.Y(_07792_),
    .B(net10),
    .A_N(_07784_));
 sg13g2_a21oi_1 _26820_ (.A1(_07791_),
    .A2(_07792_),
    .Y(_01956_),
    .B1(net563));
 sg13g2_nor2_1 _26821_ (.A(_04939_),
    .B(net81),
    .Y(_07793_));
 sg13g2_nand2_1 _26822_ (.Y(_07794_),
    .A(net959),
    .B(_07793_));
 sg13g2_o21ai_1 _26823_ (.B1(_04937_),
    .Y(_07795_),
    .A1(_04939_),
    .A2(net81));
 sg13g2_nand3_1 _26824_ (.B(_07794_),
    .C(_07795_),
    .A(net680),
    .Y(_02002_));
 sg13g2_nand2_1 _26825_ (.Y(_07796_),
    .A(net954),
    .B(_07793_));
 sg13g2_buf_1 _26826_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07797_));
 sg13g2_o21ai_1 _26827_ (.B1(_07797_),
    .Y(_07798_),
    .A1(_04939_),
    .A2(_07773_));
 sg13g2_a21oi_1 _26828_ (.A1(_07796_),
    .A2(_07798_),
    .Y(_02003_),
    .B1(_07772_));
 sg13g2_nand2_1 _26829_ (.Y(_07799_),
    .A(net855),
    .B(_07793_));
 sg13g2_o21ai_1 _26830_ (.B1(\cpu.gpio.r_src_o[6][2] ),
    .Y(_07800_),
    .A1(_04939_),
    .A2(_07773_));
 sg13g2_buf_1 _26831_ (.A(_09183_),
    .X(_07801_));
 sg13g2_a21oi_1 _26832_ (.A1(_07799_),
    .A2(_07800_),
    .Y(_02004_),
    .B1(net562));
 sg13g2_nand2_1 _26833_ (.Y(_07802_),
    .A(net1017),
    .B(_07793_));
 sg13g2_o21ai_1 _26834_ (.B1(\cpu.gpio.r_src_o[6][3] ),
    .Y(_07803_),
    .A1(_04939_),
    .A2(net81));
 sg13g2_a21oi_1 _26835_ (.A1(_07802_),
    .A2(_07803_),
    .Y(_02005_),
    .B1(net562));
 sg13g2_nor4_1 _26836_ (.A(_11726_),
    .B(net609),
    .C(net480),
    .D(_06236_),
    .Y(_07804_));
 sg13g2_buf_1 _26837_ (.A(_07804_),
    .X(_07805_));
 sg13g2_nand2_1 _26838_ (.Y(_07806_),
    .A(_09896_),
    .B(_07805_));
 sg13g2_nand2b_1 _26839_ (.Y(_07807_),
    .B(_04916_),
    .A_N(_07805_));
 sg13g2_a21oi_1 _26840_ (.A1(_07806_),
    .A2(_07807_),
    .Y(_02010_),
    .B1(_07801_));
 sg13g2_nand2_1 _26841_ (.Y(_07808_),
    .A(net954),
    .B(_07805_));
 sg13g2_nand2b_1 _26842_ (.Y(_07809_),
    .B(\cpu.gpio.r_uart_rx_src[1] ),
    .A_N(_07805_));
 sg13g2_a21oi_1 _26843_ (.A1(_07808_),
    .A2(_07809_),
    .Y(_02011_),
    .B1(net562));
 sg13g2_nand2_1 _26844_ (.Y(_07810_),
    .A(net855),
    .B(_07805_));
 sg13g2_nand2b_1 _26845_ (.Y(_07811_),
    .B(\cpu.gpio.r_uart_rx_src[2] ),
    .A_N(_07805_));
 sg13g2_a21oi_1 _26846_ (.A1(_07810_),
    .A2(_07811_),
    .Y(_02012_),
    .B1(_07801_));
 sg13g2_and2_1 _26847_ (.A(\cpu.i_wstrobe_d ),
    .B(_00316_),
    .X(_02269_));
 sg13g2_a21oi_1 _26848_ (.A1(_06269_),
    .A2(_06281_),
    .Y(_02270_),
    .B1(_06292_));
 sg13g2_xor2_1 _26849_ (.B(_06276_),
    .A(_06265_),
    .X(_07812_));
 sg13g2_nor2_1 _26850_ (.A(_06292_),
    .B(_07812_),
    .Y(_02271_));
 sg13g2_xnor2_1 _26851_ (.Y(_07813_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05025_));
 sg13g2_xnor2_1 _26852_ (.Y(_07814_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10015_));
 sg13g2_xnor2_1 _26853_ (.Y(_07815_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10038_));
 sg13g2_xnor2_1 _26854_ (.Y(_07816_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10020_));
 sg13g2_nand4_1 _26855_ (.B(_07814_),
    .C(_07815_),
    .A(_07813_),
    .Y(_07817_),
    .D(_07816_));
 sg13g2_xnor2_1 _26856_ (.Y(_07818_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05702_));
 sg13g2_xnor2_1 _26857_ (.Y(_07819_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05583_));
 sg13g2_xnor2_1 _26858_ (.Y(_07820_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05692_));
 sg13g2_xnor2_1 _26859_ (.Y(_07821_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_09983_));
 sg13g2_nand4_1 _26860_ (.B(_07819_),
    .C(_07820_),
    .A(_07818_),
    .Y(_07822_),
    .D(_07821_));
 sg13g2_xnor2_1 _26861_ (.Y(_07823_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_09972_));
 sg13g2_xnor2_1 _26862_ (.Y(_07824_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05109_));
 sg13g2_xnor2_1 _26863_ (.Y(_07825_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10010_));
 sg13g2_xnor2_1 _26864_ (.Y(_07826_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05244_));
 sg13g2_nand4_1 _26865_ (.B(_07824_),
    .C(_07825_),
    .A(_07823_),
    .Y(_07827_),
    .D(_07826_));
 sg13g2_xnor2_1 _26866_ (.Y(_07828_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_09967_));
 sg13g2_xnor2_1 _26867_ (.Y(_07829_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05436_));
 sg13g2_xnor2_1 _26868_ (.Y(_07830_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04862_));
 sg13g2_xnor2_1 _26869_ (.Y(_07831_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_09978_));
 sg13g2_nand4_1 _26870_ (.B(_07829_),
    .C(_07830_),
    .A(_07828_),
    .Y(_07832_),
    .D(_07831_));
 sg13g2_nor4_1 _26871_ (.A(_07817_),
    .B(_07822_),
    .C(_07827_),
    .D(_07832_),
    .Y(_07833_));
 sg13g2_xnor2_1 _26872_ (.Y(_07834_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05484_));
 sg13g2_xnor2_1 _26873_ (.Y(_07835_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05124_));
 sg13g2_xnor2_1 _26874_ (.Y(_07836_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10003_));
 sg13g2_xnor2_1 _26875_ (.Y(_07837_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_09991_));
 sg13g2_nand4_1 _26876_ (.B(_07835_),
    .C(_07836_),
    .A(_07834_),
    .Y(_07838_),
    .D(_07837_));
 sg13g2_xnor2_1 _26877_ (.Y(_07839_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_09968_));
 sg13g2_xnor2_1 _26878_ (.Y(_07840_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_09987_));
 sg13g2_xnor2_1 _26879_ (.Y(_07841_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05183_));
 sg13g2_xnor2_1 _26880_ (.Y(_07842_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05380_));
 sg13g2_nand4_1 _26881_ (.B(_07840_),
    .C(_07841_),
    .A(_07839_),
    .Y(_07843_),
    .D(_07842_));
 sg13g2_xnor2_1 _26882_ (.Y(_07844_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05150_));
 sg13g2_xnor2_1 _26883_ (.Y(_07845_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05673_));
 sg13g2_xnor2_1 _26884_ (.Y(_07846_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05299_));
 sg13g2_xnor2_1 _26885_ (.Y(_07847_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10027_));
 sg13g2_nand4_1 _26886_ (.B(_07845_),
    .C(_07846_),
    .A(_07844_),
    .Y(_07848_),
    .D(_07847_));
 sg13g2_xnor2_1 _26887_ (.Y(_07849_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10032_));
 sg13g2_xnor2_1 _26888_ (.Y(_07850_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_09996_));
 sg13g2_xnor2_1 _26889_ (.Y(_07851_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10045_));
 sg13g2_xnor2_1 _26890_ (.Y(_07852_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05216_));
 sg13g2_nand4_1 _26891_ (.B(_07850_),
    .C(_07851_),
    .A(_07849_),
    .Y(_07853_),
    .D(_07852_));
 sg13g2_nor4_1 _26892_ (.A(_07838_),
    .B(_07843_),
    .C(_07848_),
    .D(_07853_),
    .Y(_07854_));
 sg13g2_a22oi_1 _26893_ (.Y(_07855_),
    .B1(_07833_),
    .B2(_07854_),
    .A2(_07450_),
    .A1(net1019));
 sg13g2_nand3_1 _26894_ (.B(net123),
    .C(net399),
    .A(_09904_),
    .Y(_07856_));
 sg13g2_nand2_1 _26895_ (.Y(_07857_),
    .A(_09036_),
    .B(_07856_));
 sg13g2_a21oi_1 _26896_ (.A1(_07855_),
    .A2(_07857_),
    .Y(_02432_),
    .B1(net562));
 sg13g2_and2_1 _26897_ (.A(net123),
    .B(net401),
    .X(_07858_));
 sg13g2_buf_1 _26898_ (.A(_07858_),
    .X(_07859_));
 sg13g2_nand2_1 _26899_ (.Y(_07860_),
    .A(net1020),
    .B(_07859_));
 sg13g2_nand2_1 _26900_ (.Y(_07861_),
    .A(net123),
    .B(net401));
 sg13g2_buf_1 _26901_ (.A(_07861_),
    .X(_07862_));
 sg13g2_nand2_1 _26902_ (.Y(_07863_),
    .A(\cpu.intr.r_enable[0] ),
    .B(_07862_));
 sg13g2_a21oi_1 _26903_ (.A1(_07860_),
    .A2(_07863_),
    .Y(_02481_),
    .B1(net562));
 sg13g2_nand2_1 _26904_ (.Y(_07864_),
    .A(net954),
    .B(_07859_));
 sg13g2_nand2_1 _26905_ (.Y(_07865_),
    .A(_09037_),
    .B(_07862_));
 sg13g2_a21oi_1 _26906_ (.A1(_07864_),
    .A2(_07865_),
    .Y(_02482_),
    .B1(net562));
 sg13g2_nand2_1 _26907_ (.Y(_07866_),
    .A(net855),
    .B(_07859_));
 sg13g2_nand2_1 _26908_ (.Y(_07867_),
    .A(\cpu.intr.r_enable[2] ),
    .B(_07862_));
 sg13g2_a21oi_1 _26909_ (.A1(_07866_),
    .A2(_07867_),
    .Y(_02483_),
    .B1(net562));
 sg13g2_nand2_1 _26910_ (.Y(_07868_),
    .A(net1017),
    .B(_07859_));
 sg13g2_nand2_1 _26911_ (.Y(_07869_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_07862_));
 sg13g2_a21oi_1 _26912_ (.A1(_07868_),
    .A2(_07869_),
    .Y(_02484_),
    .B1(net562));
 sg13g2_nand2_1 _26913_ (.Y(_07870_),
    .A(net1016),
    .B(_07859_));
 sg13g2_nand2_1 _26914_ (.Y(_07871_),
    .A(_09071_),
    .B(_07862_));
 sg13g2_buf_1 _26915_ (.A(_09183_),
    .X(_07872_));
 sg13g2_a21oi_1 _26916_ (.A1(_07870_),
    .A2(_07871_),
    .Y(_02485_),
    .B1(net561));
 sg13g2_nand2_1 _26917_ (.Y(_07873_),
    .A(_09928_),
    .B(_07859_));
 sg13g2_nand2_1 _26918_ (.Y(_07874_),
    .A(\cpu.intr.r_enable[5] ),
    .B(_07862_));
 sg13g2_a21oi_1 _26919_ (.A1(_07873_),
    .A2(_07874_),
    .Y(_02486_),
    .B1(net561));
 sg13g2_nand3_1 _26920_ (.B(net123),
    .C(net399),
    .A(_09909_),
    .Y(_07875_));
 sg13g2_a221oi_1 _26921_ (.B2(_09030_),
    .C1(_09854_),
    .B1(_07875_),
    .A1(_09910_),
    .Y(_07876_),
    .A2(_07450_));
 sg13g2_nor2_1 _26922_ (.A(net564),
    .B(_07876_),
    .Y(_02487_));
 sg13g2_and2_1 _26923_ (.A(_06745_),
    .B(_06714_),
    .X(_07877_));
 sg13g2_nand4_1 _26924_ (.B(_09707_),
    .C(_06715_),
    .A(_09661_),
    .Y(_07878_),
    .D(_07877_));
 sg13g2_buf_1 _26925_ (.A(_07878_),
    .X(_07879_));
 sg13g2_o21ai_1 _26926_ (.B1(net781),
    .Y(_07880_),
    .A1(_06744_),
    .A2(_07879_));
 sg13g2_and2_1 _26927_ (.A(_09685_),
    .B(_09700_),
    .X(_07881_));
 sg13g2_o21ai_1 _26928_ (.B1(net19),
    .Y(_07882_),
    .A1(_07879_),
    .A2(_07881_));
 sg13g2_nand2b_1 _26929_ (.Y(_02517_),
    .B(_07882_),
    .A_N(_07880_));
 sg13g2_nand3b_1 _26930_ (.B(_06719_),
    .C(_09663_),
    .Y(_07883_),
    .A_N(_09685_));
 sg13g2_a21o_1 _26931_ (.A2(_07883_),
    .A1(_06744_),
    .B1(_07879_),
    .X(_07884_));
 sg13g2_nand2_1 _26932_ (.Y(_07885_),
    .A(_09685_),
    .B(_06744_));
 sg13g2_nor2_1 _26933_ (.A(net69),
    .B(_07885_),
    .Y(_07886_));
 sg13g2_o21ai_1 _26934_ (.B1(net20),
    .Y(_07887_),
    .A1(_07879_),
    .A2(_07886_));
 sg13g2_nand3_1 _26935_ (.B(_07884_),
    .C(_07887_),
    .A(net680),
    .Y(_02518_));
 sg13g2_nor2b_1 _26936_ (.A(net324),
    .B_N(_09685_),
    .Y(_07888_));
 sg13g2_buf_1 _26937_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07889_));
 sg13g2_o21ai_1 _26938_ (.B1(_07889_),
    .Y(_07890_),
    .A1(_07879_),
    .A2(_07888_));
 sg13g2_nand2b_1 _26939_ (.Y(_02519_),
    .B(_07890_),
    .A_N(_07880_));
 sg13g2_inv_1 _26940_ (.Y(_07891_),
    .A(_06719_));
 sg13g2_nor4_1 _26941_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09671_),
    .C(_09686_),
    .D(\cpu.qspi.r_state[1] ),
    .Y(_07892_));
 sg13g2_nand4_1 _26942_ (.B(_06601_),
    .C(_07877_),
    .A(_07891_),
    .Y(_07893_),
    .D(_07892_));
 sg13g2_a21oi_1 _26943_ (.A1(_09711_),
    .A2(_07893_),
    .Y(_02520_),
    .B1(_07872_));
 sg13g2_nand2_1 _26944_ (.Y(_07894_),
    .A(net1012),
    .B(_06648_));
 sg13g2_nand2_1 _26945_ (.Y(_07895_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06651_));
 sg13g2_a21oi_1 _26946_ (.A1(_07894_),
    .A2(_07895_),
    .Y(_02521_),
    .B1(_07872_));
 sg13g2_nor4_1 _26947_ (.A(net945),
    .B(_07101_),
    .C(_04872_),
    .D(_06646_),
    .Y(_07896_));
 sg13g2_a21oi_1 _26948_ (.A1(\cpu.qspi.r_mask[1] ),
    .A2(_06663_),
    .Y(_07897_),
    .B1(_07896_));
 sg13g2_nand2_1 _26949_ (.Y(_02522_),
    .A(net629),
    .B(_07897_));
 sg13g2_nor2_1 _26950_ (.A(_07101_),
    .B(_06675_),
    .Y(_07898_));
 sg13g2_a21oi_1 _26951_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06675_),
    .Y(_07899_),
    .B1(_07898_));
 sg13g2_nor2_1 _26952_ (.A(net564),
    .B(_07899_),
    .Y(_02523_));
 sg13g2_nand2_1 _26953_ (.Y(_07900_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06651_));
 sg13g2_nand2_1 _26954_ (.Y(_07901_),
    .A(net1014),
    .B(_06648_));
 sg13g2_nand3_1 _26955_ (.B(_07900_),
    .C(_07901_),
    .A(net680),
    .Y(_02524_));
 sg13g2_nor4_1 _26956_ (.A(net945),
    .B(_07097_),
    .C(_04872_),
    .D(_06646_),
    .Y(_07902_));
 sg13g2_a21oi_1 _26957_ (.A1(\cpu.qspi.r_quad[1] ),
    .A2(_06663_),
    .Y(_07903_),
    .B1(_07902_));
 sg13g2_nor2_1 _26958_ (.A(net564),
    .B(_07903_),
    .Y(_02525_));
 sg13g2_nand2_1 _26959_ (.Y(_07904_),
    .A(_07097_),
    .B(_06672_));
 sg13g2_o21ai_1 _26960_ (.B1(_07904_),
    .Y(_07905_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06672_));
 sg13g2_nand2_1 _26961_ (.Y(_02526_),
    .A(net629),
    .B(_07905_));
 sg13g2_nor2_1 _26962_ (.A(_04885_),
    .B(net95),
    .Y(_07906_));
 sg13g2_nand2_1 _26963_ (.Y(_07907_),
    .A(net959),
    .B(_07906_));
 sg13g2_o21ai_1 _26964_ (.B1(_09689_),
    .Y(_07908_),
    .A1(_04885_),
    .A2(net95));
 sg13g2_nand3_1 _26965_ (.B(_07907_),
    .C(_07908_),
    .A(net680),
    .Y(_02539_));
 sg13g2_nand2_1 _26966_ (.Y(_07909_),
    .A(net954),
    .B(_07906_));
 sg13g2_o21ai_1 _26967_ (.B1(_09690_),
    .Y(_07910_),
    .A1(_04885_),
    .A2(net95));
 sg13g2_nand3_1 _26968_ (.B(_07909_),
    .C(_07910_),
    .A(net680),
    .Y(_02540_));
 sg13g2_nor4_1 _26969_ (.A(_11666_),
    .B(net1101),
    .C(_11664_),
    .D(_06719_),
    .Y(_07911_));
 sg13g2_nor2b_1 _26970_ (.A(_06603_),
    .B_N(_07911_),
    .Y(_07912_));
 sg13g2_or3_1 _26971_ (.A(_11664_),
    .B(_06719_),
    .C(_07912_),
    .X(_07913_));
 sg13g2_inv_1 _26972_ (.Y(_07914_),
    .A(_06743_));
 sg13g2_nor3_1 _26973_ (.A(_11665_),
    .B(_09738_),
    .C(_09683_),
    .Y(_07915_));
 sg13g2_nand4_1 _26974_ (.B(_06612_),
    .C(_06714_),
    .A(_09661_),
    .Y(_07916_),
    .D(_07915_));
 sg13g2_a21oi_1 _26975_ (.A1(_11666_),
    .A2(_07914_),
    .Y(_07917_),
    .B1(_07916_));
 sg13g2_mux2_1 _26976_ (.A0(net3),
    .A1(_07913_),
    .S(_07917_),
    .X(_07918_));
 sg13g2_and2_1 _26977_ (.A(net645),
    .B(_07918_),
    .X(_02541_));
 sg13g2_nor2_1 _26978_ (.A(net6),
    .B(_07917_),
    .Y(_07919_));
 sg13g2_a21oi_1 _26979_ (.A1(_09703_),
    .A2(_07912_),
    .Y(_07920_),
    .B1(_11664_));
 sg13g2_and2_1 _26980_ (.A(_07917_),
    .B(_07920_),
    .X(_07921_));
 sg13g2_nor3_1 _26981_ (.A(net679),
    .B(_07919_),
    .C(_07921_),
    .Y(_02542_));
 sg13g2_nor3_1 _26982_ (.A(_09116_),
    .B(_09105_),
    .C(_09136_),
    .Y(_07922_));
 sg13g2_nor3_1 _26983_ (.A(_09114_),
    .B(_09194_),
    .C(_07922_),
    .Y(_07923_));
 sg13g2_buf_1 _26984_ (.A(_07923_),
    .X(_07924_));
 sg13g2_nand3_1 _26985_ (.B(net1029),
    .C(_07924_),
    .A(_09142_),
    .Y(_07925_));
 sg13g2_o21ai_1 _26986_ (.B1(_07925_),
    .Y(_07926_),
    .A1(_09142_),
    .A2(_07924_));
 sg13g2_nand2_1 _26987_ (.Y(_02548_),
    .A(net629),
    .B(_07926_));
 sg13g2_nand2_1 _26988_ (.Y(_07927_),
    .A(_09142_),
    .B(_11687_));
 sg13g2_a21oi_1 _26989_ (.A1(_07924_),
    .A2(_07927_),
    .Y(_07928_),
    .B1(_09143_));
 sg13g2_inv_1 _26990_ (.Y(_07929_),
    .A(_09142_));
 sg13g2_and4_1 _26991_ (.A(_07929_),
    .B(_09143_),
    .C(_11687_),
    .D(_07924_),
    .X(_07930_));
 sg13g2_o21ai_1 _26992_ (.B1(net629),
    .Y(_02549_),
    .A1(_07928_),
    .A2(_07930_));
 sg13g2_nor2_1 _26993_ (.A(_09142_),
    .B(_09143_),
    .Y(_07931_));
 sg13g2_or2_1 _26994_ (.X(_07932_),
    .B(_07931_),
    .A(_00226_));
 sg13g2_a21oi_1 _26995_ (.A1(_07924_),
    .A2(_07932_),
    .Y(_07933_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _26996_ (.A(\cpu.spi.r_bits[2] ),
    .B(_11687_),
    .C(_07931_),
    .D(_07924_),
    .X(_07934_));
 sg13g2_o21ai_1 _26997_ (.B1(net629),
    .Y(_02550_),
    .A1(_07933_),
    .A2(_07934_));
 sg13g2_buf_1 _26998_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_07935_));
 sg13g2_inv_1 _26999_ (.Y(_07936_),
    .A(net1063));
 sg13g2_a21oi_1 _27000_ (.A1(_09134_),
    .A2(_09104_),
    .Y(_07937_),
    .B1(_06866_));
 sg13g2_inv_1 _27001_ (.Y(_07938_),
    .A(\cpu.spi.r_state[3] ));
 sg13g2_nand2_1 _27002_ (.Y(_07939_),
    .A(_07938_),
    .B(_09106_));
 sg13g2_nand2_1 _27003_ (.Y(_07940_),
    .A(_09140_),
    .B(_07939_));
 sg13g2_nor3_1 _27004_ (.A(_09177_),
    .B(_09139_),
    .C(_07939_),
    .Y(_07941_));
 sg13g2_a21oi_1 _27005_ (.A1(_11696_),
    .A2(net867),
    .Y(_07942_),
    .B1(_09009_));
 sg13g2_nor3_1 _27006_ (.A(_00278_),
    .B(_07941_),
    .C(_07942_),
    .Y(_07943_));
 sg13g2_a21oi_1 _27007_ (.A1(_00278_),
    .A2(_07940_),
    .Y(_07944_),
    .B1(_07943_));
 sg13g2_nand2b_1 _27008_ (.Y(_07945_),
    .B(_07944_),
    .A_N(_07937_));
 sg13g2_nor3_1 _27009_ (.A(_11690_),
    .B(net867),
    .C(_07945_),
    .Y(_07946_));
 sg13g2_inv_1 _27010_ (.Y(_07947_),
    .A(_07945_));
 sg13g2_a21oi_1 _27011_ (.A1(_07939_),
    .A2(_07947_),
    .Y(_07948_),
    .B1(net779));
 sg13g2_o21ai_1 _27012_ (.B1(_07948_),
    .Y(_02583_),
    .A1(_07936_),
    .A2(_07946_));
 sg13g2_buf_1 _27013_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_07949_));
 sg13g2_nand3_1 _27014_ (.B(_11707_),
    .C(_07947_),
    .A(_11704_),
    .Y(_07950_));
 sg13g2_nand2_1 _27015_ (.Y(_07951_),
    .A(net1062),
    .B(_07950_));
 sg13g2_nand2_1 _27016_ (.Y(_02584_),
    .A(_07948_),
    .B(_07951_));
 sg13g2_buf_1 _27017_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_07952_));
 sg13g2_inv_1 _27018_ (.Y(_07953_),
    .A(net1061));
 sg13g2_nor3_1 _27019_ (.A(_11704_),
    .B(_11707_),
    .C(_07945_),
    .Y(_07954_));
 sg13g2_o21ai_1 _27020_ (.B1(_07948_),
    .Y(_02585_),
    .A1(_07953_),
    .A2(_07954_));
 sg13g2_or2_1 _27021_ (.X(_07955_),
    .B(_09104_),
    .A(_06866_));
 sg13g2_o21ai_1 _27022_ (.B1(_06867_),
    .Y(_07956_),
    .A1(_09191_),
    .A2(_07955_));
 sg13g2_nand2_1 _27023_ (.Y(_07957_),
    .A(net377),
    .B(_09172_));
 sg13g2_a22oi_1 _27024_ (.Y(_07958_),
    .B1(_07957_),
    .B2(net1029),
    .A2(_07956_),
    .A1(_09121_));
 sg13g2_buf_1 _27025_ (.A(_07958_),
    .X(_07959_));
 sg13g2_o21ai_1 _27026_ (.B1(_07959_),
    .Y(_07960_),
    .A1(_09116_),
    .A2(net1028));
 sg13g2_a22oi_1 _27027_ (.Y(_07961_),
    .B1(_07960_),
    .B2(_09038_),
    .A2(_07959_),
    .A1(_09137_));
 sg13g2_nor2_1 _27028_ (.A(net564),
    .B(_07961_),
    .Y(_02594_));
 sg13g2_nand2b_1 _27029_ (.Y(_07962_),
    .B(_09009_),
    .A_N(\cpu.spi.r_ready ));
 sg13g2_nand2_1 _27030_ (.Y(_07963_),
    .A(_07938_),
    .B(_07922_));
 sg13g2_nand4_1 _27031_ (.B(_09135_),
    .C(_07959_),
    .A(_07938_),
    .Y(_07964_),
    .D(_07963_));
 sg13g2_a21oi_1 _27032_ (.A1(_07962_),
    .A2(_07964_),
    .Y(_07965_),
    .B1(net1029));
 sg13g2_a21oi_1 _27033_ (.A1(_07959_),
    .A2(_07963_),
    .Y(_07966_),
    .B1(\cpu.spi.r_ready ));
 sg13g2_o21ai_1 _27034_ (.B1(net629),
    .Y(_02609_),
    .A1(_07965_),
    .A2(_07966_));
 sg13g2_nand2_1 _27035_ (.Y(_07967_),
    .A(_09175_),
    .B(_07924_));
 sg13g2_nand2_1 _27036_ (.Y(_07968_),
    .A(\cpu.spi.r_searching ),
    .B(_07967_));
 sg13g2_or3_1 _27037_ (.A(net801),
    .B(_09095_),
    .C(_07967_),
    .X(_07969_));
 sg13g2_a21oi_1 _27038_ (.A1(_07968_),
    .A2(_07969_),
    .Y(_02610_),
    .B1(net561));
 sg13g2_and3_1 _27039_ (.X(_07970_),
    .A(net864),
    .B(_07167_),
    .C(_06234_));
 sg13g2_buf_1 _27040_ (.A(_07970_),
    .X(_07971_));
 sg13g2_and2_1 _27041_ (.A(_04948_),
    .B(_07971_),
    .X(_07972_));
 sg13g2_buf_2 _27042_ (.A(_07972_),
    .X(_07973_));
 sg13g2_nand2_1 _27043_ (.Y(_07974_),
    .A(net959),
    .B(_07973_));
 sg13g2_nand2_1 _27044_ (.Y(_07975_),
    .A(_04948_),
    .B(_07971_));
 sg13g2_buf_2 _27045_ (.A(_07975_),
    .X(_07976_));
 sg13g2_nand2_1 _27046_ (.Y(_07977_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_07976_));
 sg13g2_nand3_1 _27047_ (.B(_07974_),
    .C(_07977_),
    .A(net680),
    .Y(_02632_));
 sg13g2_and2_1 _27048_ (.A(_04894_),
    .B(_07971_),
    .X(_07978_));
 sg13g2_buf_2 _27049_ (.A(_07978_),
    .X(_07979_));
 sg13g2_nand2_1 _27050_ (.Y(_07980_),
    .A(net855),
    .B(_07979_));
 sg13g2_nand2b_1 _27051_ (.Y(_07981_),
    .B(_09802_),
    .A_N(_07979_));
 sg13g2_a21oi_1 _27052_ (.A1(_07980_),
    .A2(_07981_),
    .Y(_02633_),
    .B1(net561));
 sg13g2_nand2_1 _27053_ (.Y(_07982_),
    .A(net1017),
    .B(_07979_));
 sg13g2_nand2b_1 _27054_ (.Y(_07983_),
    .B(\cpu.uart.r_div_value[11] ),
    .A_N(_07979_));
 sg13g2_a21oi_1 _27055_ (.A1(_07982_),
    .A2(_07983_),
    .Y(_02634_),
    .B1(net561));
 sg13g2_nand2_1 _27056_ (.Y(_07984_),
    .A(net1019),
    .B(_07973_));
 sg13g2_nand2_1 _27057_ (.Y(_07985_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27058_ (.A1(_07984_),
    .A2(_07985_),
    .Y(_02635_),
    .B1(net561));
 sg13g2_nand2_1 _27059_ (.Y(_07986_),
    .A(net855),
    .B(_07973_));
 sg13g2_nand2_1 _27060_ (.Y(_07987_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27061_ (.A1(_07986_),
    .A2(_07987_),
    .Y(_02636_),
    .B1(net561));
 sg13g2_nand2_1 _27062_ (.Y(_07988_),
    .A(net1017),
    .B(_07973_));
 sg13g2_nand2_1 _27063_ (.Y(_07989_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27064_ (.A1(_07988_),
    .A2(_07989_),
    .Y(_02637_),
    .B1(net561));
 sg13g2_nand2_1 _27065_ (.Y(_07990_),
    .A(net1016),
    .B(_07973_));
 sg13g2_nand2_1 _27066_ (.Y(_07991_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27067_ (.A1(_07990_),
    .A2(_07991_),
    .Y(_02638_),
    .B1(net626));
 sg13g2_nand2_1 _27068_ (.Y(_07992_),
    .A(net1015),
    .B(_07973_));
 sg13g2_nand2_1 _27069_ (.Y(_07993_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27070_ (.A1(_07992_),
    .A2(_07993_),
    .Y(_02639_),
    .B1(net626));
 sg13g2_nand2_1 _27071_ (.Y(_07994_),
    .A(net1014),
    .B(_07973_));
 sg13g2_nand2_1 _27072_ (.Y(_07995_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27073_ (.A1(_07994_),
    .A2(_07995_),
    .Y(_02640_),
    .B1(net626));
 sg13g2_nand2_1 _27074_ (.Y(_07996_),
    .A(net1012),
    .B(_07973_));
 sg13g2_nand2_1 _27075_ (.Y(_07997_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_07976_));
 sg13g2_a21oi_1 _27076_ (.A1(_07996_),
    .A2(_07997_),
    .Y(_02641_),
    .B1(net626));
 sg13g2_nand2_1 _27077_ (.Y(_07998_),
    .A(net1020),
    .B(_07979_));
 sg13g2_nand2b_1 _27078_ (.Y(_07999_),
    .B(\cpu.uart.r_div_value[8] ),
    .A_N(_07979_));
 sg13g2_a21oi_1 _27079_ (.A1(_07998_),
    .A2(_07999_),
    .Y(_02642_),
    .B1(net626));
 sg13g2_nand2_1 _27080_ (.Y(_08000_),
    .A(net1019),
    .B(_07979_));
 sg13g2_nand2b_1 _27081_ (.Y(_08001_),
    .B(\cpu.uart.r_div_value[9] ),
    .A_N(_07979_));
 sg13g2_a21oi_1 _27082_ (.A1(_08000_),
    .A2(_08001_),
    .Y(_02643_),
    .B1(net626));
 sg13g2_nand3_1 _27083_ (.B(_04870_),
    .C(_07971_),
    .A(_09904_),
    .Y(_08002_));
 sg13g2_nand3_1 _27084_ (.B(_07167_),
    .C(_11721_),
    .A(_05043_),
    .Y(_08003_));
 sg13g2_or3_1 _27085_ (.A(net953),
    .B(_09096_),
    .C(_08003_),
    .X(_08004_));
 sg13g2_nand4_1 _27086_ (.B(net781),
    .C(_08002_),
    .A(_09034_),
    .Y(_08005_),
    .D(_08004_));
 sg13g2_nand2b_1 _27087_ (.Y(_02667_),
    .B(_08005_),
    .A_N(_07166_));
 sg13g2_and2_1 _27088_ (.A(net461),
    .B(_07971_),
    .X(_08006_));
 sg13g2_buf_1 _27089_ (.A(_08006_),
    .X(_08007_));
 sg13g2_nand2_1 _27090_ (.Y(_08008_),
    .A(net1019),
    .B(_08007_));
 sg13g2_nand2b_1 _27091_ (.Y(_08009_),
    .B(\cpu.uart.r_r_invert ),
    .A_N(_08007_));
 sg13g2_a21oi_1 _27092_ (.A1(_08008_),
    .A2(_08009_),
    .Y(_02668_),
    .B1(net626));
 sg13g2_a21oi_1 _27093_ (.A1(_07158_),
    .A2(net342),
    .Y(_08010_),
    .B1(net1067));
 sg13g2_a21oi_1 _27094_ (.A1(_07159_),
    .A2(net342),
    .Y(_08011_),
    .B1(_07228_));
 sg13g2_a221oi_1 _27095_ (.B2(_08010_),
    .C1(_08011_),
    .B1(_07157_),
    .A1(_07156_),
    .Y(_08012_),
    .A2(net1067));
 sg13g2_a21oi_1 _27096_ (.A1(_07150_),
    .A2(_08012_),
    .Y(_08013_),
    .B1(_07225_));
 sg13g2_buf_2 _27097_ (.A(_08013_),
    .X(_08014_));
 sg13g2_o21ai_1 _27098_ (.B1(_08014_),
    .Y(_08015_),
    .A1(net923),
    .A2(_07228_));
 sg13g2_xnor2_1 _27099_ (.Y(_08016_),
    .A(_07159_),
    .B(_08015_));
 sg13g2_nor2_1 _27100_ (.A(net618),
    .B(_08016_),
    .Y(_02671_));
 sg13g2_o21ai_1 _27101_ (.B1(_08014_),
    .Y(_08017_),
    .A1(_07158_),
    .A2(_07153_));
 sg13g2_nand2_1 _27102_ (.Y(_08018_),
    .A(net1066),
    .B(_08017_));
 sg13g2_nand2b_1 _27103_ (.Y(_08019_),
    .B(net923),
    .A_N(_07153_));
 sg13g2_o21ai_1 _27104_ (.B1(_08019_),
    .Y(_08020_),
    .A1(net923),
    .A2(_07227_));
 sg13g2_nand3_1 _27105_ (.B(_08014_),
    .C(_08020_),
    .A(_07226_),
    .Y(_08021_));
 sg13g2_a21oi_1 _27106_ (.A1(_08018_),
    .A2(_08021_),
    .Y(_02672_),
    .B1(_07391_));
 sg13g2_nand2_1 _27107_ (.Y(_08022_),
    .A(_07158_),
    .B(net1066));
 sg13g2_nor3_1 _27108_ (.A(net923),
    .B(net924),
    .C(_08022_),
    .Y(_08023_));
 sg13g2_o21ai_1 _27109_ (.B1(_08014_),
    .Y(_08024_),
    .A1(net924),
    .A2(_07236_));
 sg13g2_a22oi_1 _27110_ (.Y(_08025_),
    .B1(_08024_),
    .B2(net923),
    .A2(_08023_),
    .A1(_08014_));
 sg13g2_nor2_1 _27111_ (.A(net618),
    .B(_08025_),
    .Y(_02673_));
 sg13g2_a21oi_1 _27112_ (.A1(_07236_),
    .A2(_08014_),
    .Y(_08026_),
    .B1(net924));
 sg13g2_nor2b_1 _27113_ (.A(net923),
    .B_N(net1066),
    .Y(_08027_));
 sg13g2_a21oi_1 _27114_ (.A1(_08014_),
    .A2(_08027_),
    .Y(_08028_),
    .B1(_09183_));
 sg13g2_nor2b_1 _27115_ (.A(_08026_),
    .B_N(_08028_),
    .Y(_02674_));
 sg13g2_a21oi_1 _27116_ (.A1(net342),
    .A2(_07188_),
    .Y(_08029_),
    .B1(_09033_));
 sg13g2_a21oi_1 _27117_ (.A1(_09895_),
    .A2(_04870_),
    .Y(_08030_),
    .B1(net402));
 sg13g2_o21ai_1 _27118_ (.B1(_09033_),
    .Y(_08031_),
    .A1(_07168_),
    .A2(_08030_));
 sg13g2_o21ai_1 _27119_ (.B1(_08031_),
    .Y(_08032_),
    .A1(net922),
    .A2(_08029_));
 sg13g2_o21ai_1 _27120_ (.B1(net666),
    .Y(_08033_),
    .A1(_00223_),
    .A2(_04867_));
 sg13g2_nand4_1 _27121_ (.B(_07971_),
    .C(_07181_),
    .A(_04851_),
    .Y(_08034_),
    .D(_08033_));
 sg13g2_nor2b_1 _27122_ (.A(_07177_),
    .B_N(_09033_),
    .Y(_08035_));
 sg13g2_a22oi_1 _27123_ (.Y(_08036_),
    .B1(_08034_),
    .B2(_08035_),
    .A2(_08032_),
    .A1(_07177_));
 sg13g2_nor2_1 _27124_ (.A(net618),
    .B(_08036_),
    .Y(_02676_));
 sg13g2_nand2_1 _27125_ (.Y(_08037_),
    .A(net1020),
    .B(_08007_));
 sg13g2_nand2b_1 _27126_ (.Y(_08038_),
    .B(\cpu.uart.r_x_invert ),
    .A_N(_08007_));
 sg13g2_a21oi_1 _27127_ (.A1(_08037_),
    .A2(_08038_),
    .Y(_02677_),
    .B1(net626));
 sg13g2_nand2_1 _27128_ (.Y(_08039_),
    .A(_07172_),
    .B(net922));
 sg13g2_nor3_1 _27129_ (.A(_07246_),
    .B(_07169_),
    .C(_08039_),
    .Y(_08040_));
 sg13g2_a21o_1 _27130_ (.A2(_07254_),
    .A1(net920),
    .B1(_08040_),
    .X(_08041_));
 sg13g2_o21ai_1 _27131_ (.B1(_07261_),
    .Y(_08042_),
    .A1(_07169_),
    .A2(_07266_));
 sg13g2_a21oi_1 _27132_ (.A1(_07258_),
    .A2(_08041_),
    .Y(_08043_),
    .B1(_08042_));
 sg13g2_buf_1 _27133_ (.A(_08043_),
    .X(_08044_));
 sg13g2_inv_1 _27134_ (.Y(_08045_),
    .A(_08044_));
 sg13g2_o21ai_1 _27135_ (.B1(net922),
    .Y(_08046_),
    .A1(_07190_),
    .A2(_07263_));
 sg13g2_nor3_1 _27136_ (.A(_07274_),
    .B(_08045_),
    .C(_08046_),
    .Y(_08047_));
 sg13g2_o21ai_1 _27137_ (.B1(net781),
    .Y(_08048_),
    .A1(net922),
    .A2(_08044_));
 sg13g2_nor2_1 _27138_ (.A(_08047_),
    .B(_08048_),
    .Y(_02680_));
 sg13g2_o21ai_1 _27139_ (.B1(_08044_),
    .Y(_08049_),
    .A1(net922),
    .A2(_07274_));
 sg13g2_nor2b_1 _27140_ (.A(_07172_),
    .B_N(net922),
    .Y(_08050_));
 sg13g2_nor2_1 _27141_ (.A(_07274_),
    .B(_08045_),
    .Y(_08051_));
 sg13g2_a22oi_1 _27142_ (.Y(_08052_),
    .B1(_08050_),
    .B2(_08051_),
    .A2(_08049_),
    .A1(_07172_));
 sg13g2_nor2_1 _27143_ (.A(net618),
    .B(_08052_),
    .Y(_02681_));
 sg13g2_inv_1 _27144_ (.Y(_08053_),
    .A(_08039_));
 sg13g2_nand3b_1 _27145_ (.B(_08053_),
    .C(_08044_),
    .Y(_08054_),
    .A_N(net920));
 sg13g2_nand2_1 _27146_ (.Y(_08055_),
    .A(net920),
    .B(_08039_));
 sg13g2_a21oi_1 _27147_ (.A1(_08054_),
    .A2(_08055_),
    .Y(_08056_),
    .B1(net921));
 sg13g2_a221oi_1 _27148_ (.B2(net920),
    .C1(_08056_),
    .B1(_08045_),
    .A1(_07190_),
    .Y(_08057_),
    .A2(_07265_));
 sg13g2_nor2_1 _27149_ (.A(net618),
    .B(_08057_),
    .Y(_02682_));
 sg13g2_nand2_1 _27150_ (.Y(_08058_),
    .A(_07190_),
    .B(_07265_));
 sg13g2_o21ai_1 _27151_ (.B1(_08058_),
    .Y(_08059_),
    .A1(_07248_),
    .A2(_08039_));
 sg13g2_o21ai_1 _27152_ (.B1(_08044_),
    .Y(_08060_),
    .A1(net920),
    .A2(_08053_));
 sg13g2_a22oi_1 _27153_ (.Y(_08061_),
    .B1(_08060_),
    .B2(net921),
    .A2(_08059_),
    .A1(_08044_));
 sg13g2_nor2_1 _27154_ (.A(net618),
    .B(_08061_),
    .Y(_02683_));
 sg13g2_nand2_1 _27155_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .A(_07464_),
    .B(_07458_));
 sg13g2_nand2_1 _27156_ (.Y(_08062_),
    .A(_06601_),
    .B(_07892_));
 sg13g2_nor4_1 _27157_ (.A(_09662_),
    .B(_06719_),
    .C(_06713_),
    .D(_08062_),
    .Y(_08063_));
 sg13g2_nand2_1 _27158_ (.Y(_08064_),
    .A(_06745_),
    .B(_08063_));
 sg13g2_o21ai_1 _27159_ (.B1(_09676_),
    .Y(\cpu.qspi.c_rstrobe_d ),
    .A1(_09679_),
    .A2(_08064_));
 sg13g2_nor3_1 _27160_ (.A(_09738_),
    .B(_09677_),
    .C(net671),
    .Y(_08065_));
 sg13g2_a22oi_1 _27161_ (.Y(_08066_),
    .B1(_08063_),
    .B2(_08065_),
    .A2(net671),
    .A1(_09671_));
 sg13g2_nor2_1 _27162_ (.A(net927),
    .B(_08066_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27163_ (.A(_00189_),
    .B(_08066_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27164_ (.S0(_04916_),
    .A0(_09051_),
    .A1(_09043_),
    .A2(_09045_),
    .A3(_09055_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08067_));
 sg13g2_mux4_1 _27165_ (.S0(_04916_),
    .A0(_09065_),
    .A1(_09061_),
    .A2(_09067_),
    .A3(_09063_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08068_));
 sg13g2_mux2_1 _27166_ (.A0(_08067_),
    .A1(_08068_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27167_ (.S0(_04919_),
    .A0(net1084),
    .A1(net1085),
    .A2(net1063),
    .A3(net1062),
    .S1(_05323_),
    .X(_08069_));
 sg13g2_mux4_1 _27168_ (.S0(_04919_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_05323_),
    .X(_08070_));
 sg13g2_nor2b_1 _27169_ (.A(_05389_),
    .B_N(_08070_),
    .Y(_08071_));
 sg13g2_a21oi_1 _27170_ (.A1(_05389_),
    .A2(_08069_),
    .Y(_08072_),
    .B1(_08071_));
 sg13g2_nand2b_1 _27171_ (.Y(_08073_),
    .B(net1061),
    .A_N(_04919_));
 sg13g2_nand3_1 _27172_ (.B(_05323_),
    .C(net1064),
    .A(_04919_),
    .Y(_08074_));
 sg13g2_o21ai_1 _27173_ (.B1(_08074_),
    .Y(_08075_),
    .A1(_05323_),
    .A2(_08073_));
 sg13g2_nand3_1 _27174_ (.B(_00187_),
    .C(_08075_),
    .A(_05425_),
    .Y(_08076_));
 sg13g2_o21ai_1 _27175_ (.B1(_08076_),
    .Y(net15),
    .A1(_05425_),
    .A2(_08072_));
 sg13g2_mux4_1 _27176_ (.S0(_05509_),
    .A0(net1084),
    .A1(net1085),
    .A2(net1063),
    .A3(net1062),
    .S1(_05572_),
    .X(_08077_));
 sg13g2_mux4_1 _27177_ (.S0(_05509_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_05572_),
    .X(_08078_));
 sg13g2_nor2b_1 _27178_ (.A(_05661_),
    .B_N(_08078_),
    .Y(_08079_));
 sg13g2_a21oi_1 _27179_ (.A1(_05661_),
    .A2(_08077_),
    .Y(_08080_),
    .B1(_08079_));
 sg13g2_nand2b_1 _27180_ (.Y(_08081_),
    .B(net1061),
    .A_N(_05509_));
 sg13g2_nand3_1 _27181_ (.B(_05572_),
    .C(net1064),
    .A(_05509_),
    .Y(_08082_));
 sg13g2_o21ai_1 _27182_ (.B1(_08082_),
    .Y(_08083_),
    .A1(_05572_),
    .A2(_08081_));
 sg13g2_nand3_1 _27183_ (.B(_00186_),
    .C(_08083_),
    .A(_05003_),
    .Y(_08084_));
 sg13g2_o21ai_1 _27184_ (.B1(_08084_),
    .Y(net16),
    .A1(_05003_),
    .A2(_08080_));
 sg13g2_mux4_1 _27185_ (.S0(_04925_),
    .A0(net1084),
    .A1(net1085),
    .A2(net1063),
    .A3(net1062),
    .S1(_06252_),
    .X(_08085_));
 sg13g2_mux4_1 _27186_ (.S0(_04925_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_06252_),
    .X(_08086_));
 sg13g2_nor2b_1 _27187_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08086_),
    .Y(_08087_));
 sg13g2_a21oi_1 _27188_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08085_),
    .Y(_08088_),
    .B1(_08087_));
 sg13g2_nand2b_1 _27189_ (.Y(_08089_),
    .B(net1061),
    .A_N(_04925_));
 sg13g2_nand3_1 _27190_ (.B(net1064),
    .C(_06252_),
    .A(_04925_),
    .Y(_08090_));
 sg13g2_o21ai_1 _27191_ (.B1(_08090_),
    .Y(_08091_),
    .A1(_06252_),
    .A2(_08089_));
 sg13g2_nand3_1 _27192_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08091_),
    .A(_00106_),
    .Y(_08092_));
 sg13g2_o21ai_1 _27193_ (.B1(_08092_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08088_));
 sg13g2_mux4_1 _27194_ (.S0(_05496_),
    .A0(net1084),
    .A1(net1085),
    .A2(net1063),
    .A3(net1062),
    .S1(_06253_),
    .X(_08093_));
 sg13g2_mux4_1 _27195_ (.S0(_05496_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_06253_),
    .X(_08094_));
 sg13g2_nor2b_1 _27196_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08094_),
    .Y(_08095_));
 sg13g2_a21oi_1 _27197_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08093_),
    .Y(_08096_),
    .B1(_08095_));
 sg13g2_nand2b_1 _27198_ (.Y(_08097_),
    .B(net1061),
    .A_N(_05496_));
 sg13g2_nand3_1 _27199_ (.B(net1064),
    .C(_06253_),
    .A(_05496_),
    .Y(_08098_));
 sg13g2_o21ai_1 _27200_ (.B1(_08098_),
    .Y(_08099_),
    .A1(_06253_),
    .A2(_08097_));
 sg13g2_nand3_1 _27201_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08099_),
    .A(_00146_),
    .Y(_08100_));
 sg13g2_o21ai_1 _27202_ (.B1(_08100_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08096_));
 sg13g2_xor2_1 _27203_ (.B(clknet_leaf_72_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27204_ (.S0(_05493_),
    .A0(net1084),
    .A1(net1085),
    .A2(net1063),
    .A3(net1062),
    .S1(_06255_),
    .X(_08101_));
 sg13g2_mux4_1 _27205_ (.S0(_05493_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_06255_),
    .X(_08102_));
 sg13g2_nor2b_1 _27206_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08102_),
    .Y(_08103_));
 sg13g2_a21oi_1 _27207_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08101_),
    .Y(_08104_),
    .B1(_08103_));
 sg13g2_nand2b_1 _27208_ (.Y(_08105_),
    .B(net1061),
    .A_N(_05493_));
 sg13g2_nand3_1 _27209_ (.B(net1064),
    .C(_06255_),
    .A(_05493_),
    .Y(_08106_));
 sg13g2_o21ai_1 _27210_ (.B1(_08106_),
    .Y(_08107_),
    .A1(_06255_),
    .A2(_08105_));
 sg13g2_nand3_1 _27211_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08107_),
    .A(_00149_),
    .Y(_08108_));
 sg13g2_o21ai_1 _27212_ (.B1(_08108_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08104_));
 sg13g2_mux4_1 _27213_ (.S0(_04943_),
    .A0(net1084),
    .A1(net1085),
    .A2(_07935_),
    .A3(_07949_),
    .S1(_06258_),
    .X(_08109_));
 sg13g2_mux4_1 _27214_ (.S0(_04943_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(_07252_),
    .A2(_11758_),
    .A3(_11741_),
    .S1(_06258_),
    .X(_08110_));
 sg13g2_nor2b_1 _27215_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08110_),
    .Y(_08111_));
 sg13g2_a21oi_1 _27216_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08109_),
    .Y(_08112_),
    .B1(_08111_));
 sg13g2_nand2b_1 _27217_ (.Y(_08113_),
    .B(net1061),
    .A_N(_04943_));
 sg13g2_nand3_1 _27218_ (.B(net1064),
    .C(_06258_),
    .A(_04943_),
    .Y(_08114_));
 sg13g2_o21ai_1 _27219_ (.B1(_08114_),
    .Y(_08115_),
    .A1(_06258_),
    .A2(_08113_));
 sg13g2_nand3_1 _27220_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08115_),
    .A(_00108_),
    .Y(_08116_));
 sg13g2_o21ai_1 _27221_ (.B1(_08116_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08112_));
 sg13g2_mux4_1 _27222_ (.S0(_05511_),
    .A0(net1084),
    .A1(net1085),
    .A2(_07935_),
    .A3(_07949_),
    .S1(_06259_),
    .X(_08117_));
 sg13g2_mux4_1 _27223_ (.S0(_05511_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(_07252_),
    .A2(_11758_),
    .A3(_11741_),
    .S1(_06259_),
    .X(_08118_));
 sg13g2_nor2b_1 _27224_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08118_),
    .Y(_08119_));
 sg13g2_a21oi_1 _27225_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08117_),
    .Y(_08120_),
    .B1(_08119_));
 sg13g2_nand2b_1 _27226_ (.Y(_08121_),
    .B(net1061),
    .A_N(_05511_));
 sg13g2_nand3_1 _27227_ (.B(net1064),
    .C(_06259_),
    .A(_05511_),
    .Y(_08122_));
 sg13g2_o21ai_1 _27228_ (.B1(_08122_),
    .Y(_08123_),
    .A1(_06259_),
    .A2(_08121_));
 sg13g2_nand3_1 _27229_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08123_),
    .A(_00148_),
    .Y(_08124_));
 sg13g2_o21ai_1 _27230_ (.B1(_08124_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08120_));
 sg13g2_mux4_1 _27231_ (.S0(_04937_),
    .A0(_11739_),
    .A1(_11736_),
    .A2(net1063),
    .A3(net1062),
    .S1(_07797_),
    .X(_08125_));
 sg13g2_mux4_1 _27232_ (.S0(_04937_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_07797_),
    .X(_08126_));
 sg13g2_nor2b_1 _27233_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08126_),
    .Y(_08127_));
 sg13g2_a21oi_1 _27234_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08125_),
    .Y(_08128_),
    .B1(_08127_));
 sg13g2_nand2b_1 _27235_ (.Y(_08129_),
    .B(_07952_),
    .A_N(_04937_));
 sg13g2_nand3_1 _27236_ (.B(_07889_),
    .C(_07797_),
    .A(_04937_),
    .Y(_08130_));
 sg13g2_o21ai_1 _27237_ (.B1(_08130_),
    .Y(_08131_),
    .A1(_07797_),
    .A2(_08129_));
 sg13g2_nand3_1 _27238_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08131_),
    .A(_00107_),
    .Y(_08132_));
 sg13g2_o21ai_1 _27239_ (.B1(_08132_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08128_));
 sg13g2_mux4_1 _27240_ (.S0(_05498_),
    .A0(net1084),
    .A1(net1085),
    .A2(net1063),
    .A3(net1062),
    .S1(_06261_),
    .X(_08133_));
 sg13g2_mux4_1 _27241_ (.S0(_05498_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1065),
    .A2(net1082),
    .A3(net1083),
    .S1(_06261_),
    .X(_08134_));
 sg13g2_nor2b_1 _27242_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08134_),
    .Y(_08135_));
 sg13g2_a21oi_1 _27243_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08133_),
    .Y(_08136_),
    .B1(_08135_));
 sg13g2_nand2b_1 _27244_ (.Y(_08137_),
    .B(_07952_),
    .A_N(_05498_));
 sg13g2_nand3_1 _27245_ (.B(net1064),
    .C(_06261_),
    .A(_05498_),
    .Y(_08138_));
 sg13g2_o21ai_1 _27246_ (.B1(_08138_),
    .Y(_08139_),
    .A1(_06261_),
    .A2(_08137_));
 sg13g2_nand3_1 _27247_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08139_),
    .A(_00147_),
    .Y(_08140_));
 sg13g2_o21ai_1 _27248_ (.B1(_08140_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08136_));
 sg13g2_dfrbp_1 _27249_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1118),
    .D(_00317_),
    .Q_N(_14749_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27250_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1119),
    .D(_00318_),
    .Q_N(_14748_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27251_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1120),
    .D(_00319_),
    .Q_N(_14747_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27252_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1121),
    .D(_00320_),
    .Q_N(_14746_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27253_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1122),
    .D(_00321_),
    .Q_N(_14745_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27255_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27256_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1123),
    .D(_00322_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1124),
    .D(_00323_),
    .Q_N(_00103_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1125),
    .D(_00324_),
    .Q_N(_00113_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1126),
    .D(_00325_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1127),
    .D(_00326_),
    .Q_N(_00131_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1128),
    .D(_00327_),
    .Q_N(_00143_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1129),
    .D(_00328_),
    .Q_N(_00155_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1130),
    .D(_00329_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1131),
    .D(_00330_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1132),
    .D(_00331_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1133),
    .D(_00332_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1134),
    .D(_00333_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1135),
    .D(_00334_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1136),
    .D(_00335_),
    .Q_N(_00129_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1137),
    .D(_00336_),
    .Q_N(_00141_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1138),
    .D(_00337_),
    .Q_N(_00153_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1139),
    .D(_00338_),
    .Q_N(_00311_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1140),
    .D(_00339_),
    .Q_N(_00092_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1141),
    .D(_00340_),
    .Q_N(_00102_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1142),
    .D(_00341_),
    .Q_N(_00112_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1143),
    .D(_00342_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1144),
    .D(_00343_),
    .Q_N(_00130_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1145),
    .D(_00344_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1146),
    .D(_00345_),
    .Q_N(_00142_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1147),
    .D(_00346_),
    .Q_N(_00154_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1148),
    .D(_00347_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1149),
    .D(_00348_),
    .Q_N(_00121_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1150),
    .D(_00349_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1151),
    .D(_00350_),
    .Q_N(_00140_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1152),
    .D(_00351_),
    .Q_N(_00152_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1153),
    .D(_00352_),
    .Q_N(_00312_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1154),
    .D(_00353_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1155),
    .D(_00354_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1156),
    .D(_00355_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1157),
    .D(_00356_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1158),
    .D(_00357_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1159),
    .D(_00358_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1160),
    .D(_00359_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1161),
    .D(_00360_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1162),
    .D(_00361_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1163),
    .D(_00362_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1164),
    .D(_00363_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1165),
    .D(_00364_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1166),
    .D(_00365_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1167),
    .D(_00366_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1168),
    .D(_00367_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1169),
    .D(_00368_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1170),
    .D(_00369_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1171),
    .D(_00370_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1172),
    .D(_00371_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1173),
    .D(_00372_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1174),
    .D(_00373_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1175),
    .D(_00374_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1176),
    .D(_00375_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1177),
    .D(_00376_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1178),
    .D(_00377_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1179),
    .D(_00378_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1180),
    .D(_00379_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1181),
    .D(_00380_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1182),
    .D(_00381_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1183),
    .D(_00382_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1184),
    .D(_00383_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1185),
    .D(_00384_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1186),
    .D(_00385_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1187),
    .D(_00386_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1188),
    .D(_00387_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1189),
    .D(_00388_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1190),
    .D(_00389_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1191),
    .D(_00390_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1192),
    .D(_00391_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1193),
    .D(_00392_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1194),
    .D(_00393_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1195),
    .D(_00394_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1196),
    .D(_00395_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1197),
    .D(_00396_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1198),
    .D(_00397_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1199),
    .D(_00398_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1200),
    .D(_00399_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1201),
    .D(_00400_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1202),
    .D(_00401_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1203),
    .D(_00402_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1204),
    .D(_00403_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1205),
    .D(_00404_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1206),
    .D(_00405_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1207),
    .D(_00406_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1208),
    .D(_00407_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1209),
    .D(_00408_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1210),
    .D(_00409_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1211),
    .D(_00410_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1212),
    .D(_00411_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1213),
    .D(_00412_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1214),
    .D(_00413_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1215),
    .D(_00414_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1216),
    .D(_00415_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1217),
    .D(_00416_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1218),
    .D(_00417_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1219),
    .D(_00418_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1220),
    .D(_00419_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1221),
    .D(_00420_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1222),
    .D(_00421_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1223),
    .D(_00422_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1224),
    .D(_00423_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1225),
    .D(_00424_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1226),
    .D(_00425_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1227),
    .D(_00426_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1228),
    .D(_00427_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1229),
    .D(_00428_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1230),
    .D(_00429_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1231),
    .D(_00430_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1232),
    .D(_00431_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1233),
    .D(_00432_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1234),
    .D(_00433_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1235),
    .D(_00434_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1236),
    .D(_00435_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1237),
    .D(_00436_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1238),
    .D(_00437_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1239),
    .D(_00438_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1240),
    .D(_00439_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1241),
    .D(_00440_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1242),
    .D(_00441_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1243),
    .D(_00442_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1244),
    .D(_00443_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1245),
    .D(_00444_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1246),
    .D(_00445_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1247),
    .D(_00446_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1248),
    .D(_00447_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1249),
    .D(_00448_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1250),
    .D(_00449_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1251),
    .D(_00450_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1252),
    .D(_00451_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1253),
    .D(_00452_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1254),
    .D(_00453_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1255),
    .D(_00454_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1256),
    .D(_00455_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1257),
    .D(_00456_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1258),
    .D(_00457_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1259),
    .D(_00458_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1260),
    .D(_00459_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1261),
    .D(_00460_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1262),
    .D(_00461_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1263),
    .D(_00462_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1264),
    .D(_00463_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1265),
    .D(_00464_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1266),
    .D(_00465_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1267),
    .D(_00466_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1268),
    .D(_00467_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1269),
    .D(_00468_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1270),
    .D(_00469_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1271),
    .D(_00470_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1272),
    .D(_00471_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1273),
    .D(_00472_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1274),
    .D(_00473_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1275),
    .D(_00474_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1276),
    .D(_00475_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1277),
    .D(_00476_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1278),
    .D(_00477_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1279),
    .D(_00478_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1280),
    .D(_00479_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1281),
    .D(_00480_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1282),
    .D(_00481_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1283),
    .D(_00482_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1284),
    .D(_00483_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1285),
    .D(_00484_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1286),
    .D(_00485_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1287),
    .D(_00486_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1288),
    .D(_00487_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1289),
    .D(_00488_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1290),
    .D(_00489_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1291),
    .D(_00490_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1292),
    .D(_00491_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1293),
    .D(_00492_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1294),
    .D(_00493_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1295),
    .D(_00494_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1296),
    .D(_00495_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1297),
    .D(_00496_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1298),
    .D(_00497_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1299),
    .D(_00498_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1300),
    .D(_00499_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1301),
    .D(_00500_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1302),
    .D(_00501_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1303),
    .D(_00502_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1304),
    .D(_00503_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1305),
    .D(_00504_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1306),
    .D(_00505_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1307),
    .D(_00506_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1308),
    .D(_00507_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1309),
    .D(_00508_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1310),
    .D(_00509_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1311),
    .D(_00510_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1312),
    .D(_00511_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1313),
    .D(_00512_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1314),
    .D(_00513_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1315),
    .D(_00514_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1316),
    .D(_00515_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1317),
    .D(_00516_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1318),
    .D(_00517_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1319),
    .D(_00518_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1320),
    .D(_00519_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1321),
    .D(_00520_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1322),
    .D(_00521_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1323),
    .D(_00522_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1324),
    .D(_00523_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1325),
    .D(_00524_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1326),
    .D(_00525_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1327),
    .D(_00526_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1328),
    .D(_00527_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1329),
    .D(_00528_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1330),
    .D(_00529_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1331),
    .D(_00530_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1332),
    .D(_00531_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1333),
    .D(_00532_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1334),
    .D(_00533_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1335),
    .D(_00534_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1336),
    .D(_00535_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1337),
    .D(_00536_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1338),
    .D(_00537_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1339),
    .D(_00538_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1340),
    .D(_00539_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1341),
    .D(_00540_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1342),
    .D(_00541_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1343),
    .D(_00542_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1344),
    .D(_00543_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1345),
    .D(_00544_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1346),
    .D(_00545_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1347),
    .D(_00546_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1348),
    .D(_00547_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1349),
    .D(_00548_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1350),
    .D(_00549_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1351),
    .D(_00550_),
    .Q_N(_14543_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1352),
    .D(_00551_),
    .Q_N(_14542_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1353),
    .D(_00552_),
    .Q_N(_14541_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1354),
    .D(_00553_),
    .Q_N(_14540_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1355),
    .D(_00554_),
    .Q_N(_14539_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1356),
    .D(_00555_),
    .Q_N(_14538_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1357),
    .D(_00556_),
    .Q_N(_14537_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1358),
    .D(_00557_),
    .Q_N(_14536_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1359),
    .D(_00558_),
    .Q_N(_14535_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1360),
    .D(_00559_),
    .Q_N(_14534_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1361),
    .D(_00560_),
    .Q_N(_14533_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1362),
    .D(_00561_),
    .Q_N(_14532_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1363),
    .D(_00562_),
    .Q_N(_14531_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1364),
    .D(_00563_),
    .Q_N(_14530_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1365),
    .D(_00564_),
    .Q_N(_14529_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1366),
    .D(_00565_),
    .Q_N(_14528_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1367),
    .D(_00566_),
    .Q_N(_14527_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1368),
    .D(_00567_),
    .Q_N(_14526_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1369),
    .D(_00568_),
    .Q_N(_14525_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1370),
    .D(_00569_),
    .Q_N(_14524_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1371),
    .D(_00570_),
    .Q_N(_14523_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1372),
    .D(_00571_),
    .Q_N(_14522_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1373),
    .D(_00572_),
    .Q_N(_14521_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1374),
    .D(_00573_),
    .Q_N(_14520_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1375),
    .D(_00574_),
    .Q_N(_14519_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1376),
    .D(_00575_),
    .Q_N(_14518_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1377),
    .D(_00576_),
    .Q_N(_14517_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1378),
    .D(_00577_),
    .Q_N(_14516_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1379),
    .D(_00578_),
    .Q_N(_14515_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1380),
    .D(_00579_),
    .Q_N(_14514_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1381),
    .D(_00580_),
    .Q_N(_14513_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1382),
    .D(_00581_),
    .Q_N(_14512_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1383),
    .D(_00582_),
    .Q_N(_14511_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1384),
    .D(_00583_),
    .Q_N(_14510_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1385),
    .D(_00584_),
    .Q_N(_14509_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1386),
    .D(_00585_),
    .Q_N(_14508_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1387),
    .D(_00586_),
    .Q_N(_00315_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1388),
    .D(_00587_),
    .Q_N(_14507_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1389),
    .D(_00588_),
    .Q_N(_00276_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1390),
    .D(_00589_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1391),
    .D(_00590_),
    .Q_N(_00246_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1392),
    .D(_00591_),
    .Q_N(_00247_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1393),
    .D(_00592_),
    .Q_N(_00248_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1394),
    .D(_00593_),
    .Q_N(_00249_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1395),
    .D(_00594_),
    .Q_N(_00250_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1396),
    .D(_00595_),
    .Q_N(_14506_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1397),
    .D(_00596_),
    .Q_N(_14505_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1398),
    .D(_00597_),
    .Q_N(_14504_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1399),
    .D(_00598_),
    .Q_N(_00251_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1400),
    .D(_00599_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1401),
    .D(_00600_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1402),
    .D(_00601_),
    .Q_N(_00236_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1403),
    .D(_00602_),
    .Q_N(_00238_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1404),
    .D(_00603_),
    .Q_N(_00240_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1405),
    .D(_00604_),
    .Q_N(_00242_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1406),
    .D(_00605_),
    .Q_N(_00243_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1407),
    .D(_00606_),
    .Q_N(_00244_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1408),
    .D(_00607_),
    .Q_N(_00245_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1409),
    .D(_00608_),
    .Q_N(_14503_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1410),
    .D(_00609_),
    .Q_N(_14502_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1411),
    .D(_00610_),
    .Q_N(_14501_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1412),
    .D(_00611_),
    .Q_N(_14500_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1413),
    .D(_00612_),
    .Q_N(_14499_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1414),
    .D(_00613_),
    .Q_N(_14498_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1415),
    .D(_00614_),
    .Q_N(_14497_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1416),
    .D(_00615_),
    .Q_N(_14496_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1417),
    .D(_00616_),
    .Q_N(_14495_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1418),
    .D(_00617_),
    .Q_N(_14494_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1419),
    .D(_00618_),
    .Q_N(_14493_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1420),
    .D(_00619_),
    .Q_N(_14492_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1421),
    .D(_00620_),
    .Q_N(_14491_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1422),
    .D(_00621_),
    .Q_N(_14490_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1423),
    .D(_00622_),
    .Q_N(_14489_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1424),
    .D(_00623_),
    .Q_N(_14488_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1425),
    .D(_00624_),
    .Q_N(_14487_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1426),
    .D(_00625_),
    .Q_N(_14486_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1427),
    .D(_00626_),
    .Q_N(_14485_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1428),
    .D(_00627_),
    .Q_N(_14484_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1429),
    .D(_00628_),
    .Q_N(_14483_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1430),
    .D(_00629_),
    .Q_N(_14482_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1431),
    .D(_00630_),
    .Q_N(_14481_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1432),
    .D(_00631_),
    .Q_N(_14480_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1433),
    .D(_00632_),
    .Q_N(_14479_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1434),
    .D(_00633_),
    .Q_N(_14478_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1435),
    .D(_00634_),
    .Q_N(_14477_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1436),
    .D(_00635_),
    .Q_N(_14476_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1437),
    .D(_00636_),
    .Q_N(_14475_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1438),
    .D(_00637_),
    .Q_N(_14474_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1439),
    .D(_00638_),
    .Q_N(_14473_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1440),
    .D(_00639_),
    .Q_N(_14472_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1441),
    .D(_00640_),
    .Q_N(_14471_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1442),
    .D(_00641_),
    .Q_N(_14470_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1443),
    .D(_00642_),
    .Q_N(_14469_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1444),
    .D(_00643_),
    .Q_N(_14468_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1445),
    .D(_00644_),
    .Q_N(_14467_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1446),
    .D(_00645_),
    .Q_N(_14466_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1447),
    .D(_00646_),
    .Q_N(_14465_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1448),
    .D(_00647_),
    .Q_N(_14464_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1449),
    .D(_00648_),
    .Q_N(_14463_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1450),
    .D(_00649_),
    .Q_N(_14462_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1451),
    .D(_00650_),
    .Q_N(_14461_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1452),
    .D(_00651_),
    .Q_N(_14460_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1453),
    .D(_00652_),
    .Q_N(_14459_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1454),
    .D(_00653_),
    .Q_N(_14458_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1455),
    .D(_00654_),
    .Q_N(_14457_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1456),
    .D(_00655_),
    .Q_N(_14456_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1457),
    .D(_00656_),
    .Q_N(_14455_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1458),
    .D(_00657_),
    .Q_N(_14454_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1459),
    .D(_00658_),
    .Q_N(_14453_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1460),
    .D(_00659_),
    .Q_N(_14452_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1461),
    .D(_00660_),
    .Q_N(_14451_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1462),
    .D(_00661_),
    .Q_N(_14450_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1463),
    .D(_00662_),
    .Q_N(_14449_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1464),
    .D(_00663_),
    .Q_N(_14448_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1465),
    .D(_00664_),
    .Q_N(_14447_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1466),
    .D(_00665_),
    .Q_N(_14446_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1467),
    .D(_00666_),
    .Q_N(_14445_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1468),
    .D(_00667_),
    .Q_N(_14444_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1469),
    .D(_00668_),
    .Q_N(_14443_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1470),
    .D(_00669_),
    .Q_N(_14442_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1471),
    .D(_00670_),
    .Q_N(_14441_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1472),
    .D(_00671_),
    .Q_N(_14440_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1473),
    .D(_00672_),
    .Q_N(_14439_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1474),
    .D(_00673_),
    .Q_N(_14438_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1475),
    .D(_00674_),
    .Q_N(_14437_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1476),
    .D(_00675_),
    .Q_N(_14436_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1477),
    .D(_00676_),
    .Q_N(_14435_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1478),
    .D(_00677_),
    .Q_N(_14434_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1479),
    .D(_00678_),
    .Q_N(_14433_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1480),
    .D(_00679_),
    .Q_N(_14432_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1481),
    .D(_00680_),
    .Q_N(_14431_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1482),
    .D(_00681_),
    .Q_N(_14430_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1483),
    .D(_00682_),
    .Q_N(_14429_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1484),
    .D(_00683_),
    .Q_N(_14428_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1485),
    .D(_00684_),
    .Q_N(_14427_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1486),
    .D(_00685_),
    .Q_N(_14426_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1487),
    .D(_00686_),
    .Q_N(_14425_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1488),
    .D(_00687_),
    .Q_N(_14424_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1489),
    .D(_00688_),
    .Q_N(_14423_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1490),
    .D(_00689_),
    .Q_N(_14422_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1491),
    .D(_00690_),
    .Q_N(_14421_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1492),
    .D(_00691_),
    .Q_N(_14420_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1493),
    .D(_00692_),
    .Q_N(_14419_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1494),
    .D(_00693_),
    .Q_N(_14418_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1495),
    .D(_00694_),
    .Q_N(_14417_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1496),
    .D(_00695_),
    .Q_N(_14416_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1497),
    .D(_00696_),
    .Q_N(_14415_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1498),
    .D(_00697_),
    .Q_N(_14414_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1499),
    .D(_00698_),
    .Q_N(_14413_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1500),
    .D(_00699_),
    .Q_N(_14412_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1501),
    .D(_00700_),
    .Q_N(_14411_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1502),
    .D(_00701_),
    .Q_N(_14410_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1503),
    .D(_00702_),
    .Q_N(_14409_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1504),
    .D(_00703_),
    .Q_N(_14408_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1505),
    .D(_00704_),
    .Q_N(_14407_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1506),
    .D(_00705_),
    .Q_N(_14406_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1507),
    .D(_00706_),
    .Q_N(_14405_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1508),
    .D(_00707_),
    .Q_N(_14404_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1509),
    .D(_00708_),
    .Q_N(_14403_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1510),
    .D(_00709_),
    .Q_N(_14402_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1511),
    .D(_00710_),
    .Q_N(_14401_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1512),
    .D(_00711_),
    .Q_N(_14400_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1513),
    .D(_00712_),
    .Q_N(_14399_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1514),
    .D(_00713_),
    .Q_N(_14398_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1515),
    .D(_00714_),
    .Q_N(_14397_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1516),
    .D(_00715_),
    .Q_N(_14396_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1517),
    .D(_00716_),
    .Q_N(_14395_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1518),
    .D(_00717_),
    .Q_N(_14394_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1519),
    .D(_00718_),
    .Q_N(_14393_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1520),
    .D(_00719_),
    .Q_N(_14392_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1521),
    .D(_00720_),
    .Q_N(_14391_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1522),
    .D(_00721_),
    .Q_N(_14390_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1523),
    .D(_00722_),
    .Q_N(_14389_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1524),
    .D(_00723_),
    .Q_N(_14388_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1525),
    .D(_00724_),
    .Q_N(_14387_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1526),
    .D(_00725_),
    .Q_N(_14386_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1527),
    .D(_00726_),
    .Q_N(_14385_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1528),
    .D(_00727_),
    .Q_N(_14384_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1529),
    .D(_00728_),
    .Q_N(_14383_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1530),
    .D(_00729_),
    .Q_N(_14382_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1531),
    .D(_00730_),
    .Q_N(_14381_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1532),
    .D(_00731_),
    .Q_N(_14380_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1533),
    .D(_00732_),
    .Q_N(_14379_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1534),
    .D(_00733_),
    .Q_N(_14378_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1535),
    .D(_00734_),
    .Q_N(_14377_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1536),
    .D(_00735_),
    .Q_N(_14376_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1537),
    .D(_00736_),
    .Q_N(_14375_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1538),
    .D(_00737_),
    .Q_N(_14374_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1539),
    .D(_00738_),
    .Q_N(_14373_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1540),
    .D(_00739_),
    .Q_N(_14372_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1541),
    .D(_00740_),
    .Q_N(_14371_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1542),
    .D(_00741_),
    .Q_N(_14370_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1543),
    .D(_00742_),
    .Q_N(_14369_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1544),
    .D(_00743_),
    .Q_N(_14368_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1545),
    .D(_00744_),
    .Q_N(_14367_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1546),
    .D(_00745_),
    .Q_N(_14366_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1547),
    .D(_00746_),
    .Q_N(_14365_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1548),
    .D(_00747_),
    .Q_N(_14364_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1549),
    .D(_00748_),
    .Q_N(_14363_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1550),
    .D(_00749_),
    .Q_N(_14362_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1551),
    .D(_00750_),
    .Q_N(_00298_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1552),
    .D(_00751_),
    .Q_N(_14361_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1553),
    .D(_00752_),
    .Q_N(_00273_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1554),
    .D(_00753_),
    .Q_N(_14360_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1555),
    .D(_00754_),
    .Q_N(_14359_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1556),
    .D(_00755_),
    .Q_N(_14358_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1557),
    .D(_00756_),
    .Q_N(_14357_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1558),
    .D(_00757_),
    .Q_N(_14356_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1559),
    .D(_00758_),
    .Q_N(_14355_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1560),
    .D(_00759_),
    .Q_N(_14354_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1561),
    .D(_00760_),
    .Q_N(_14353_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1562),
    .D(_00761_),
    .Q_N(_14352_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1563),
    .D(_00762_),
    .Q_N(_14351_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1564),
    .D(_00763_),
    .Q_N(_14350_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1565),
    .D(_00764_),
    .Q_N(_14349_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1566),
    .D(_00765_),
    .Q_N(_14348_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1567),
    .D(_00766_),
    .Q_N(_14347_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1568),
    .D(_00767_),
    .Q_N(_14346_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1569),
    .D(_00768_),
    .Q_N(_14345_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1570),
    .D(_00769_),
    .Q_N(_14344_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1571),
    .D(_00770_),
    .Q_N(_14343_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1572),
    .D(_00771_),
    .Q_N(_14342_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1573),
    .D(_00772_),
    .Q_N(_14341_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1574),
    .D(_00773_),
    .Q_N(_14340_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1575),
    .D(_00774_),
    .Q_N(_00258_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1576),
    .D(_00775_),
    .Q_N(_14339_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1577),
    .D(_00776_),
    .Q_N(_14338_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1578),
    .D(_00777_),
    .Q_N(_14750_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1579),
    .D(_00011_),
    .Q_N(_14751_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1580),
    .D(_00012_),
    .Q_N(_14752_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1581),
    .D(_00013_),
    .Q_N(_14753_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1582),
    .D(_00014_),
    .Q_N(_14754_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1583),
    .D(_00015_),
    .Q_N(_14755_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1584),
    .D(_00016_),
    .Q_N(_14756_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1585),
    .D(_00017_),
    .Q_N(_14757_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1586),
    .D(_00018_),
    .Q_N(_14758_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1587),
    .D(_00019_),
    .Q_N(_14759_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1588),
    .D(_00020_),
    .Q_N(_14337_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1589),
    .D(_00778_),
    .Q_N(_14336_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1590),
    .D(_00779_),
    .Q_N(_14335_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1591),
    .D(_00780_),
    .Q_N(_14334_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1592),
    .D(_00781_),
    .Q_N(_14760_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1593),
    .D(_00052_),
    .Q_N(_14333_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1594),
    .D(_00782_),
    .Q_N(_14332_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1595),
    .D(_00783_),
    .Q_N(_14331_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1596),
    .D(_00784_),
    .Q_N(_14330_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1597),
    .D(_00785_),
    .Q_N(_14329_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1598),
    .D(_00786_),
    .Q_N(_14328_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1599),
    .D(_00787_),
    .Q_N(_14327_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1600),
    .D(_00788_),
    .Q_N(_14326_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1601),
    .D(_00789_),
    .Q_N(_14325_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_inv$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1602),
    .D(_00790_),
    .Q_N(_14324_),
    .Q(\cpu.dec.r_rs2_inv ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1603),
    .D(_00791_),
    .Q_N(_14323_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1604),
    .D(_00792_),
    .Q_N(_14322_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1605),
    .D(_00793_),
    .Q_N(_00310_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1606),
    .D(_00794_),
    .Q_N(_14321_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1607),
    .D(_00795_),
    .Q_N(_00274_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1608),
    .D(_00796_),
    .Q_N(_14320_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1609),
    .D(_00797_),
    .Q_N(_14319_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1610),
    .D(_00798_),
    .Q_N(_00192_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1611),
    .D(_00799_),
    .Q_N(_14761_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1612),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00193_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1613),
    .D(_00800_),
    .Q_N(_14318_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1614),
    .D(_00801_),
    .Q_N(_14317_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1615),
    .D(_00802_),
    .Q_N(_14316_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1616),
    .D(_00803_),
    .Q_N(_14315_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1617),
    .D(_00804_),
    .Q_N(_14314_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1618),
    .D(_00805_),
    .Q_N(_14313_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1619),
    .D(_00806_),
    .Q_N(_14312_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1620),
    .D(_00807_),
    .Q_N(_14311_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1621),
    .D(_00808_),
    .Q_N(_14310_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1622),
    .D(_00809_),
    .Q_N(_14309_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1623),
    .D(_00810_),
    .Q_N(_14308_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1624),
    .D(_00811_),
    .Q_N(_14307_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1625),
    .D(_00812_),
    .Q_N(_14306_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1626),
    .D(_00813_),
    .Q_N(_14305_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1627),
    .D(_00814_),
    .Q_N(_14304_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1628),
    .D(_00815_),
    .Q_N(_14303_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1629),
    .D(_00816_),
    .Q_N(_14302_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1630),
    .D(_00817_),
    .Q_N(_14301_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1631),
    .D(_00818_),
    .Q_N(_14300_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1632),
    .D(_00819_),
    .Q_N(_14299_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1633),
    .D(_00820_),
    .Q_N(_14298_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1634),
    .D(_00821_),
    .Q_N(_14297_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1635),
    .D(_00822_),
    .Q_N(_14296_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1636),
    .D(_00823_),
    .Q_N(_14295_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1637),
    .D(_00824_),
    .Q_N(_14294_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1638),
    .D(_00825_),
    .Q_N(_14293_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1639),
    .D(_00826_),
    .Q_N(_14292_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1640),
    .D(_00827_),
    .Q_N(_14291_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1641),
    .D(_00828_),
    .Q_N(_14290_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1642),
    .D(_00829_),
    .Q_N(_14289_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1643),
    .D(_00830_),
    .Q_N(_14288_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1644),
    .D(_00831_),
    .Q_N(_14287_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1645),
    .D(_00832_),
    .Q_N(_14286_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1646),
    .D(_00833_),
    .Q_N(_14285_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1647),
    .D(_00834_),
    .Q_N(_14284_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1648),
    .D(_00835_),
    .Q_N(_14283_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1649),
    .D(_00836_),
    .Q_N(_14282_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1650),
    .D(_00837_),
    .Q_N(_14281_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1651),
    .D(_00838_),
    .Q_N(_14280_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1652),
    .D(_00839_),
    .Q_N(_14279_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1653),
    .D(_00840_),
    .Q_N(_14278_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1654),
    .D(_00841_),
    .Q_N(_14277_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1655),
    .D(_00842_),
    .Q_N(_14276_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1656),
    .D(_00843_),
    .Q_N(_14275_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1657),
    .D(_00844_),
    .Q_N(_14274_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1658),
    .D(_00845_),
    .Q_N(_14273_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1659),
    .D(_00846_),
    .Q_N(_14272_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1660),
    .D(_00847_),
    .Q_N(_14271_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1661),
    .D(_00848_),
    .Q_N(_14270_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1662),
    .D(_00849_),
    .Q_N(_14269_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1663),
    .D(_00850_),
    .Q_N(_14268_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1664),
    .D(_00851_),
    .Q_N(_14267_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1665),
    .D(_00852_),
    .Q_N(_14266_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1666),
    .D(_00853_),
    .Q_N(_14265_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1667),
    .D(_00854_),
    .Q_N(_14264_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1668),
    .D(_00855_),
    .Q_N(_14263_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1669),
    .D(_00856_),
    .Q_N(_14262_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1670),
    .D(_00857_),
    .Q_N(_14261_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1671),
    .D(_00858_),
    .Q_N(_14260_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1672),
    .D(_00859_),
    .Q_N(_14259_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1673),
    .D(_00860_),
    .Q_N(_14258_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1674),
    .D(_00861_),
    .Q_N(_14257_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1675),
    .D(_00862_),
    .Q_N(_14256_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1676),
    .D(_00863_),
    .Q_N(_14255_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1677),
    .D(_00864_),
    .Q_N(_14254_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1678),
    .D(_00865_),
    .Q_N(_14253_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1679),
    .D(_00866_),
    .Q_N(_14252_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1680),
    .D(_00867_),
    .Q_N(_14251_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1681),
    .D(_00868_),
    .Q_N(_14250_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1682),
    .D(_00869_),
    .Q_N(_14249_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1683),
    .D(_00870_),
    .Q_N(_14248_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1684),
    .D(_00871_),
    .Q_N(_14247_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1685),
    .D(_00872_),
    .Q_N(_14246_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1686),
    .D(_00873_),
    .Q_N(_14245_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1687),
    .D(_00874_),
    .Q_N(_14244_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1688),
    .D(_00875_),
    .Q_N(_14243_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1689),
    .D(_00876_),
    .Q_N(_14242_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1690),
    .D(_00877_),
    .Q_N(_14241_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1691),
    .D(_00878_),
    .Q_N(_14240_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1692),
    .D(_00879_),
    .Q_N(_14239_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1693),
    .D(_00880_),
    .Q_N(_14238_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1694),
    .D(_00881_),
    .Q_N(_14237_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1695),
    .D(_00882_),
    .Q_N(_00268_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1696),
    .D(_00883_),
    .Q_N(_00269_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1697),
    .D(_00884_),
    .Q_N(_00270_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1698),
    .D(_00885_),
    .Q_N(_00271_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1699),
    .D(_00886_),
    .Q_N(_00272_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1700),
    .D(_00887_),
    .Q_N(_14236_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1701),
    .D(_00888_),
    .Q_N(_00259_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1702),
    .D(_00889_),
    .Q_N(_00260_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1703),
    .D(_00890_),
    .Q_N(_00261_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1704),
    .D(_00891_),
    .Q_N(_00262_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1705),
    .D(_00892_),
    .Q_N(_00263_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1706),
    .D(_00893_),
    .Q_N(_00264_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1707),
    .D(_00894_),
    .Q_N(_00265_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1708),
    .D(_00895_),
    .Q_N(_00266_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1709),
    .D(_00896_),
    .Q_N(_00267_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1710),
    .D(_00897_),
    .Q_N(_14235_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1711),
    .D(_00898_),
    .Q_N(_14234_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1712),
    .D(_00899_),
    .Q_N(_14233_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1713),
    .D(_00900_),
    .Q_N(_14232_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1714),
    .D(_00901_),
    .Q_N(_14231_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1715),
    .D(_00902_),
    .Q_N(_14230_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1716),
    .D(_00903_),
    .Q_N(_14229_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1717),
    .D(_00904_),
    .Q_N(_14228_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1718),
    .D(_00905_),
    .Q_N(_14227_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1719),
    .D(_00906_),
    .Q_N(_14226_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1720),
    .D(_00907_),
    .Q_N(_14225_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1721),
    .D(_00908_),
    .Q_N(_14224_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1722),
    .D(_00909_),
    .Q_N(_14223_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1723),
    .D(_00910_),
    .Q_N(_14222_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1724),
    .D(_00911_),
    .Q_N(_14221_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1725),
    .D(_00912_),
    .Q_N(_14220_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1726),
    .D(_00913_),
    .Q_N(_14219_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1727),
    .D(_00914_),
    .Q_N(_14218_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1728),
    .D(_00915_),
    .Q_N(_14217_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1729),
    .D(_00916_),
    .Q_N(_14216_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1730),
    .D(_00917_),
    .Q_N(_14215_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1731),
    .D(_00918_),
    .Q_N(_14214_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1732),
    .D(_00919_),
    .Q_N(_14213_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1733),
    .D(_00920_),
    .Q_N(_14212_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1734),
    .D(_00921_),
    .Q_N(_14211_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1735),
    .D(_00922_),
    .Q_N(_14210_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1736),
    .D(_00923_),
    .Q_N(_14209_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1737),
    .D(_00924_),
    .Q_N(_14208_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1738),
    .D(_00925_),
    .Q_N(_14207_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1739),
    .D(_00926_),
    .Q_N(_14206_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1740),
    .D(_00927_),
    .Q_N(_14205_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1741),
    .D(_00928_),
    .Q_N(_14762_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1742),
    .D(_00053_),
    .Q_N(_14204_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_cc$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1743),
    .D(_00929_),
    .Q_N(_14203_),
    .Q(\cpu.ex.r_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1744),
    .D(_00930_),
    .Q_N(_14763_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1745),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14202_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1746),
    .D(_00931_),
    .Q_N(_14201_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1747),
    .D(_00932_),
    .Q_N(_14200_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1748),
    .D(_00933_),
    .Q_N(_14199_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1749),
    .D(_00934_),
    .Q_N(_14198_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1750),
    .D(_00935_),
    .Q_N(_14197_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1751),
    .D(_00936_),
    .Q_N(_14196_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1752),
    .D(_00937_),
    .Q_N(_14195_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1753),
    .D(_00938_),
    .Q_N(_14194_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1754),
    .D(_00939_),
    .Q_N(_14193_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1755),
    .D(_00940_),
    .Q_N(_14192_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1756),
    .D(_00941_),
    .Q_N(_14191_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1757),
    .D(_00942_),
    .Q_N(_14190_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1758),
    .D(_00943_),
    .Q_N(_14189_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1759),
    .D(_00944_),
    .Q_N(_14188_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1760),
    .D(_00945_),
    .Q_N(_14187_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1761),
    .D(_00946_),
    .Q_N(_00189_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1762),
    .D(_00947_),
    .Q_N(_14186_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1763),
    .D(_00948_),
    .Q_N(_14185_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1764),
    .D(_00949_),
    .Q_N(_14184_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1765),
    .D(_00950_),
    .Q_N(_00197_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1766),
    .D(_00951_),
    .Q_N(_14183_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1767),
    .D(_00952_),
    .Q_N(_14182_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1768),
    .D(_00953_),
    .Q_N(_14181_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1769),
    .D(_00954_),
    .Q_N(_14180_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1770),
    .D(_00955_),
    .Q_N(_14179_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1771),
    .D(_00956_),
    .Q_N(_14178_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1772),
    .D(_00957_),
    .Q_N(_14177_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1773),
    .D(_00958_),
    .Q_N(_14176_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1774),
    .D(_00959_),
    .Q_N(_14175_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1775),
    .D(_00960_),
    .Q_N(_14174_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1776),
    .D(_00961_),
    .Q_N(_14173_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1777),
    .D(_00962_),
    .Q_N(_14172_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1778),
    .D(_00963_),
    .Q_N(_14171_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1779),
    .D(_00964_),
    .Q_N(_14170_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1780),
    .D(_00965_),
    .Q_N(_14764_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1781),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14765_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1782),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_00167_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1783),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_00168_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1784),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_00169_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1785),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_00170_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1786),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00171_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1787),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14169_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1788),
    .D(_00966_),
    .Q_N(_00309_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1789),
    .D(_00967_),
    .Q_N(_00308_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1790),
    .D(_00968_),
    .Q_N(_00307_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1791),
    .D(_00969_),
    .Q_N(_00306_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1792),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14168_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1793),
    .D(_00970_),
    .Q_N(_00305_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1794),
    .D(_00971_),
    .Q_N(_00304_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1795),
    .D(_00972_),
    .Q_N(_14167_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1796),
    .D(_00973_),
    .Q_N(_00303_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1797),
    .D(_00974_),
    .Q_N(_00302_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1798),
    .D(_00975_),
    .Q_N(_00301_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1799),
    .D(_00976_),
    .Q_N(_14166_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1800),
    .D(_00977_),
    .Q_N(_00300_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1801),
    .D(_00978_),
    .Q_N(_14165_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1802),
    .D(_00979_),
    .Q_N(_14766_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1803),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_00120_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1804),
    .D(_00980_),
    .Q_N(_00299_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1805),
    .D(_00981_),
    .Q_N(_14767_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1806),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_00127_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1807),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_00139_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1808),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_00151_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1809),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_00163_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1810),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_00164_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1811),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_00165_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1812),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_00166_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1813),
    .D(net495),
    .Q_N(_14768_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1814),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14769_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1815),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14770_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1816),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14771_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1817),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00199_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1818),
    .D(_00982_),
    .Q_N(_00200_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1819),
    .D(_00983_),
    .Q_N(_00290_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1820),
    .D(_00984_),
    .Q_N(_00289_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1821),
    .D(_00985_),
    .Q_N(_00196_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1822),
    .D(_00986_),
    .Q_N(_00195_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1823),
    .D(_00987_),
    .Q_N(_00194_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1824),
    .D(_00988_),
    .Q_N(_00297_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1825),
    .D(_00989_),
    .Q_N(_00191_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1826),
    .D(_00990_),
    .Q_N(_00190_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1827),
    .D(_00991_),
    .Q_N(_00296_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1828),
    .D(_00992_),
    .Q_N(_00295_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1829),
    .D(_00993_),
    .Q_N(_00294_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1830),
    .D(_00994_),
    .Q_N(_00293_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1831),
    .D(_00995_),
    .Q_N(_00292_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1832),
    .D(_00996_),
    .Q_N(_00291_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1833),
    .D(_00997_),
    .Q_N(_14164_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1834),
    .D(_00998_),
    .Q_N(_00198_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_set_cc$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1835),
    .D(_00999_),
    .Q_N(_14163_),
    .Q(\cpu.ex.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1836),
    .D(_01000_),
    .Q_N(_14162_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1837),
    .D(_01001_),
    .Q_N(_14161_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1838),
    .D(_01002_),
    .Q_N(_14160_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1839),
    .D(_01003_),
    .Q_N(_14159_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1840),
    .D(_01004_),
    .Q_N(_14158_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1841),
    .D(_01005_),
    .Q_N(_14157_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1842),
    .D(_01006_),
    .Q_N(_14156_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1843),
    .D(_01007_),
    .Q_N(_14155_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1844),
    .D(_01008_),
    .Q_N(_14154_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1845),
    .D(_01009_),
    .Q_N(_14153_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1846),
    .D(_01010_),
    .Q_N(_14152_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1847),
    .D(_01011_),
    .Q_N(_14151_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1848),
    .D(_01012_),
    .Q_N(_14150_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1849),
    .D(_01013_),
    .Q_N(_14149_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1850),
    .D(_01014_),
    .Q_N(_14148_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1851),
    .D(_01015_),
    .Q_N(_14147_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1852),
    .D(_01016_),
    .Q_N(_14146_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1853),
    .D(_01017_),
    .Q_N(_14145_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1854),
    .D(_01018_),
    .Q_N(_14144_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1855),
    .D(_01019_),
    .Q_N(_14143_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1856),
    .D(_01020_),
    .Q_N(_14142_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1857),
    .D(_01021_),
    .Q_N(_14141_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1858),
    .D(_01022_),
    .Q_N(_14140_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1859),
    .D(_01023_),
    .Q_N(_14139_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1860),
    .D(_01024_),
    .Q_N(_14138_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1861),
    .D(_01025_),
    .Q_N(_14137_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1862),
    .D(_01026_),
    .Q_N(_14136_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1863),
    .D(_01027_),
    .Q_N(_14135_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1864),
    .D(_01028_),
    .Q_N(_14134_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1865),
    .D(_01029_),
    .Q_N(_14133_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1866),
    .D(_01030_),
    .Q_N(_14132_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1867),
    .D(_01031_),
    .Q_N(_00257_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1868),
    .D(_01032_),
    .Q_N(_00239_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1869),
    .D(_01033_),
    .Q_N(_00241_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1870),
    .D(_01034_),
    .Q_N(_14131_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1871),
    .D(_01035_),
    .Q_N(_14130_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1872),
    .D(_01036_),
    .Q_N(_14129_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1873),
    .D(_01037_),
    .Q_N(_14128_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1874),
    .D(_01038_),
    .Q_N(_00275_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1875),
    .D(_01039_),
    .Q_N(_14127_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1876),
    .D(_01040_),
    .Q_N(_00228_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1877),
    .D(_01041_),
    .Q_N(_00227_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1878),
    .D(_01042_),
    .Q_N(_00229_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1879),
    .D(_01043_),
    .Q_N(_00231_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1880),
    .D(_01044_),
    .Q_N(_00233_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1881),
    .D(_01045_),
    .Q_N(_00235_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1882),
    .D(_01046_),
    .Q_N(_00237_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1883),
    .D(_01047_),
    .Q_N(_14126_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1884),
    .D(_01048_),
    .Q_N(_14125_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1885),
    .D(_01049_),
    .Q_N(_14124_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1886),
    .D(_01050_),
    .Q_N(_14123_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1887),
    .D(_01051_),
    .Q_N(_14772_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1888),
    .D(_00054_),
    .Q_N(_00256_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1889),
    .D(_01052_),
    .Q_N(_00223_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1890),
    .D(_01053_),
    .Q_N(_14122_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1891),
    .D(_01054_),
    .Q_N(_14121_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1892),
    .D(_01055_),
    .Q_N(_14120_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1893),
    .D(_01056_),
    .Q_N(_14119_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1894),
    .D(_01057_),
    .Q_N(_14118_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1895),
    .D(_01058_),
    .Q_N(_14117_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1896),
    .D(_01059_),
    .Q_N(_00178_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1897),
    .D(_01060_),
    .Q_N(_00179_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1898),
    .D(_01061_),
    .Q_N(_00287_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1899),
    .D(_01062_),
    .Q_N(_00180_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1900),
    .D(_01063_),
    .Q_N(_00181_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1901),
    .D(_01064_),
    .Q_N(_00182_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1902),
    .D(_01065_),
    .Q_N(_00281_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1903),
    .D(_01066_),
    .Q_N(_14116_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1904),
    .D(_01067_),
    .Q_N(_14115_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1905),
    .D(_01068_),
    .Q_N(_14114_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1906),
    .D(_01069_),
    .Q_N(_14113_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1907),
    .D(_01070_),
    .Q_N(_00288_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1908),
    .D(_01071_),
    .Q_N(_14112_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1909),
    .D(_01072_),
    .Q_N(_00188_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1910),
    .D(_01073_),
    .Q_N(_14111_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1911),
    .D(_01074_),
    .Q_N(_00255_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1912),
    .D(_01075_),
    .Q_N(_14110_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1913),
    .D(_01076_),
    .Q_N(_14109_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1914),
    .D(_01077_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1915),
    .D(_01078_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1916),
    .D(_01079_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1917),
    .D(_01080_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1918),
    .D(_01081_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1919),
    .D(_01082_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1920),
    .D(_01083_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1921),
    .D(_01084_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1922),
    .D(_01085_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1923),
    .D(_01086_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1924),
    .D(_01087_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1925),
    .D(_01088_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1926),
    .D(_01089_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1927),
    .D(_01090_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1928),
    .D(_01091_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1929),
    .D(_01092_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1930),
    .D(_01093_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1931),
    .D(_01094_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1932),
    .D(_01095_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1933),
    .D(_01096_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1934),
    .D(_01097_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1935),
    .D(_01098_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1936),
    .D(_01099_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1937),
    .D(_01100_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1938),
    .D(_01101_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1939),
    .D(_01102_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1940),
    .D(_01103_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1941),
    .D(_01104_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1942),
    .D(_01105_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1943),
    .D(_01106_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1944),
    .D(_01107_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1945),
    .D(_01108_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1946),
    .D(_01109_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1947),
    .D(_01110_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1948),
    .D(_01111_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1949),
    .D(_01112_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1950),
    .D(_01113_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1951),
    .D(_01114_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1952),
    .D(_01115_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1953),
    .D(_01116_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1954),
    .D(_01117_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1955),
    .D(_01118_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1956),
    .D(_01119_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1957),
    .D(_01120_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1958),
    .D(_01121_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1959),
    .D(_01122_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1960),
    .D(_01123_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1961),
    .D(_01124_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1962),
    .D(_01125_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1963),
    .D(_01126_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1964),
    .D(_01127_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1965),
    .D(_01128_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1966),
    .D(_01129_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1967),
    .D(_01130_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1968),
    .D(_01131_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1969),
    .D(_01132_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1970),
    .D(_01133_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1971),
    .D(_01134_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1972),
    .D(_01135_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1973),
    .D(_01136_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1974),
    .D(_01137_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1975),
    .D(_01138_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1976),
    .D(_01139_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1977),
    .D(_01140_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1978),
    .D(_01141_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1979),
    .D(_01142_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1980),
    .D(_01143_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1981),
    .D(_01144_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1982),
    .D(_01145_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1983),
    .D(_01146_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1984),
    .D(_01147_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1985),
    .D(_01148_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1986),
    .D(_01149_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1987),
    .D(_01150_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1988),
    .D(_01151_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1989),
    .D(_01152_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1990),
    .D(_01153_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1991),
    .D(_01154_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1992),
    .D(_01155_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1993),
    .D(_01156_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1994),
    .D(_01157_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1995),
    .D(_01158_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1996),
    .D(_01159_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1997),
    .D(_01160_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1998),
    .D(_01161_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1999),
    .D(_01162_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2000),
    .D(_01163_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2001),
    .D(_01164_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2002),
    .D(_01165_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2003),
    .D(_01166_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2004),
    .D(_01167_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2005),
    .D(_01168_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2006),
    .D(_01169_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2007),
    .D(_01170_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2008),
    .D(_01171_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2009),
    .D(_01172_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2010),
    .D(_01173_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2011),
    .D(_01174_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2012),
    .D(_01175_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2013),
    .D(_01176_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2014),
    .D(_01177_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2015),
    .D(_01178_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2016),
    .D(_01179_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2017),
    .D(_01180_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2018),
    .D(_01181_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2019),
    .D(_01182_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2020),
    .D(_01183_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2021),
    .D(_01184_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2022),
    .D(_01185_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2023),
    .D(_01186_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2024),
    .D(_01187_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2025),
    .D(_01188_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2026),
    .D(_01189_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2027),
    .D(_01190_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2028),
    .D(_01191_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2029),
    .D(_01192_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2030),
    .D(_01193_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2031),
    .D(_01194_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2032),
    .D(_01195_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2033),
    .D(_01196_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2034),
    .D(_01197_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2035),
    .D(_01198_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2036),
    .D(_01199_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2037),
    .D(_01200_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2038),
    .D(_01201_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2039),
    .D(_01202_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2040),
    .D(_01203_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2041),
    .D(_01204_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2042),
    .D(_01205_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2043),
    .D(_01206_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2044),
    .D(_01207_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2045),
    .D(_01208_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2046),
    .D(_01209_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2047),
    .D(_01210_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2048),
    .D(_01211_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2049),
    .D(_01212_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2050),
    .D(_01213_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2051),
    .D(_01214_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2052),
    .D(_01215_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2053),
    .D(_01216_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2054),
    .D(_01217_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2055),
    .D(_01218_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2056),
    .D(_01219_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2057),
    .D(_01220_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2058),
    .D(_01221_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2059),
    .D(_01222_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2060),
    .D(_01223_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2061),
    .D(_01224_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2062),
    .D(_01225_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2063),
    .D(_01226_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2064),
    .D(_01227_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2065),
    .D(_01228_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2066),
    .D(_01229_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2067),
    .D(_01230_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2068),
    .D(_01231_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2069),
    .D(_01232_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2070),
    .D(_01233_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2071),
    .D(_01234_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2072),
    .D(_01235_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2073),
    .D(_01236_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2074),
    .D(_01237_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2075),
    .D(_01238_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2076),
    .D(_01239_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2077),
    .D(_01240_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2078),
    .D(_01241_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2079),
    .D(_01242_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2080),
    .D(_01243_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2081),
    .D(_01244_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2082),
    .D(_01245_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2083),
    .D(_01246_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2084),
    .D(_01247_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2085),
    .D(_01248_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2086),
    .D(_01249_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2087),
    .D(_01250_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2088),
    .D(_01251_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2089),
    .D(_01252_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2090),
    .D(_01253_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2091),
    .D(_01254_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2092),
    .D(_01255_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2093),
    .D(_01256_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2094),
    .D(_01257_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2095),
    .D(_01258_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2096),
    .D(_01259_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2097),
    .D(_01260_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2098),
    .D(_01261_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2099),
    .D(_01262_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2100),
    .D(_01263_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2101),
    .D(_01264_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2102),
    .D(_01265_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2103),
    .D(_01266_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2104),
    .D(_01267_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2105),
    .D(_01268_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2106),
    .D(_01269_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2107),
    .D(_01270_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2108),
    .D(_01271_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2109),
    .D(_01272_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2110),
    .D(_01273_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2111),
    .D(_01274_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2112),
    .D(_01275_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2113),
    .D(_01276_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2114),
    .D(_01277_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2115),
    .D(_01278_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2116),
    .D(_01279_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2117),
    .D(_01280_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2118),
    .D(_01281_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2119),
    .D(_01282_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2120),
    .D(_01283_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2121),
    .D(_01284_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2122),
    .D(_01285_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2123),
    .D(_01286_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2124),
    .D(_01287_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2125),
    .D(_01288_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2126),
    .D(_01289_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2127),
    .D(_01290_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2128),
    .D(_01291_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2129),
    .D(_01292_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2130),
    .D(_01293_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2131),
    .D(_01294_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2132),
    .D(_01295_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2133),
    .D(_01296_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2134),
    .D(_01297_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2135),
    .D(_01298_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2136),
    .D(_01299_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2137),
    .D(_01300_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2138),
    .D(_01301_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2139),
    .D(_01302_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2140),
    .D(_01303_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2141),
    .D(_01304_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2142),
    .D(_01305_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2143),
    .D(_01306_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2144),
    .D(_01307_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2145),
    .D(_01308_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2146),
    .D(_01309_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2147),
    .D(_01310_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2148),
    .D(_01311_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2149),
    .D(_01312_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2150),
    .D(_01313_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2151),
    .D(_01314_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2152),
    .D(_01315_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2153),
    .D(_01316_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2154),
    .D(_01317_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2155),
    .D(_01318_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2156),
    .D(_01319_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2157),
    .D(_01320_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2158),
    .D(_01321_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2159),
    .D(_01322_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2160),
    .D(_01323_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2161),
    .D(_01324_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2162),
    .D(_01325_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2163),
    .D(_01326_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2164),
    .D(_01327_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2165),
    .D(_01328_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2166),
    .D(_01329_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2167),
    .D(_01330_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2168),
    .D(_01331_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2169),
    .D(_01332_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2170),
    .D(_01333_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2171),
    .D(_01334_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2172),
    .D(_01335_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2173),
    .D(_01336_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2174),
    .D(_01337_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2175),
    .D(_01338_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2176),
    .D(_01339_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2177),
    .D(_01340_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2178),
    .D(_01341_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2179),
    .D(_01342_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2180),
    .D(_01343_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2181),
    .D(_01344_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2182),
    .D(_01345_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2183),
    .D(_01346_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2184),
    .D(_01347_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2185),
    .D(_01348_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2186),
    .D(_01349_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2187),
    .D(_01350_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2188),
    .D(_01351_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2189),
    .D(_01352_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2190),
    .D(_01353_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2191),
    .D(_01354_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2192),
    .D(_01355_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2193),
    .D(_01356_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2194),
    .D(_01357_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2195),
    .D(_01358_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2196),
    .D(_01359_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2197),
    .D(_01360_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2198),
    .D(_01361_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2199),
    .D(_01362_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2200),
    .D(_01363_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2201),
    .D(_01364_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2202),
    .D(_01365_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2203),
    .D(_01366_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2204),
    .D(_01367_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2205),
    .D(_01368_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2206),
    .D(_01369_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2207),
    .D(_01370_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2208),
    .D(_01371_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2209),
    .D(_01372_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2210),
    .D(_01373_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2211),
    .D(_01374_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2212),
    .D(_01375_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2213),
    .D(_01376_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2214),
    .D(_01377_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2215),
    .D(_01378_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2216),
    .D(_01379_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2217),
    .D(_01380_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2218),
    .D(_01381_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2219),
    .D(_01382_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2220),
    .D(_01383_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2221),
    .D(_01384_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2222),
    .D(_01385_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2223),
    .D(_01386_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2224),
    .D(_01387_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2225),
    .D(_01388_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2226),
    .D(_01389_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2227),
    .D(_01390_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2228),
    .D(_01391_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2229),
    .D(_01392_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2230),
    .D(_01393_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2231),
    .D(_01394_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2232),
    .D(_01395_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2233),
    .D(_01396_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2234),
    .D(_01397_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2235),
    .D(_01398_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2236),
    .D(_01399_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2237),
    .D(_01400_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2238),
    .D(_01401_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2239),
    .D(_01402_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2240),
    .D(_01403_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2241),
    .D(_01404_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2242),
    .D(_01405_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2243),
    .D(_01406_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2244),
    .D(_01407_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2245),
    .D(_01408_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2246),
    .D(_01409_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2247),
    .D(_01410_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2248),
    .D(_01411_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2249),
    .D(_01412_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2250),
    .D(_01413_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2251),
    .D(_01414_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2252),
    .D(_01415_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2253),
    .D(_01416_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2254),
    .D(_01417_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2255),
    .D(_01418_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2256),
    .D(_01419_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2257),
    .D(_01420_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2258),
    .D(_01421_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2259),
    .D(_01422_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2260),
    .D(_01423_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2261),
    .D(_01424_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2262),
    .D(_01425_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2263),
    .D(_01426_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2264),
    .D(_01427_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2265),
    .D(_01428_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2266),
    .D(_01429_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2267),
    .D(_01430_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2268),
    .D(_01431_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2269),
    .D(_01432_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2270),
    .D(_01433_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2271),
    .D(_01434_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2272),
    .D(_01435_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2273),
    .D(_01436_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2274),
    .D(_01437_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2275),
    .D(_01438_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2276),
    .D(_01439_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2277),
    .D(_01440_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2278),
    .D(_01441_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2279),
    .D(_01442_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2280),
    .D(_01443_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2281),
    .D(_01444_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2282),
    .D(_01445_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2283),
    .D(_01446_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2284),
    .D(_01447_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2285),
    .D(_01448_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2286),
    .D(_01449_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2287),
    .D(_01450_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2288),
    .D(_01451_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2289),
    .D(_01452_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2290),
    .D(_01453_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2291),
    .D(_01454_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2292),
    .D(_01455_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2293),
    .D(_01456_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2294),
    .D(_01457_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2295),
    .D(_01458_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2296),
    .D(_01459_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2297),
    .D(_01460_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2298),
    .D(_01461_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2299),
    .D(_01462_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2300),
    .D(_01463_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2301),
    .D(_01464_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2302),
    .D(_01465_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2303),
    .D(_01466_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2304),
    .D(_01467_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2305),
    .D(_01468_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2306),
    .D(_01469_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2307),
    .D(_01470_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2308),
    .D(_01471_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2309),
    .D(_01472_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2310),
    .D(_01473_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2311),
    .D(_01474_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2312),
    .D(_01475_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2313),
    .D(_01476_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2314),
    .D(_01477_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2315),
    .D(_01478_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2316),
    .D(_01479_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2317),
    .D(_01480_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2318),
    .D(_01481_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2319),
    .D(_01482_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2320),
    .D(_01483_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2321),
    .D(_01484_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2322),
    .D(_01485_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2323),
    .D(_01486_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2324),
    .D(_01487_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2325),
    .D(_01488_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2326),
    .D(_01489_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2327),
    .D(_01490_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2328),
    .D(_01491_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2329),
    .D(_01492_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2330),
    .D(_01493_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2331),
    .D(_01494_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2332),
    .D(_01495_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2333),
    .D(_01496_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2334),
    .D(_01497_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2335),
    .D(_01498_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2336),
    .D(_01499_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2337),
    .D(_01500_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2338),
    .D(_01501_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2339),
    .D(_01502_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2340),
    .D(_01503_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2341),
    .D(_01504_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2342),
    .D(_01505_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2343),
    .D(_01506_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2344),
    .D(_01507_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2345),
    .D(_01508_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2346),
    .D(_01509_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2347),
    .D(_01510_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2348),
    .D(_01511_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2349),
    .D(_01512_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2350),
    .D(_01513_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2351),
    .D(_01514_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2352),
    .D(_01515_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2353),
    .D(_01516_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2354),
    .D(_01517_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2355),
    .D(_01518_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2356),
    .D(_01519_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2357),
    .D(_01520_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2358),
    .D(_01521_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2359),
    .D(_01522_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2360),
    .D(_01523_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net2361),
    .D(_01524_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2362),
    .D(_01525_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2363),
    .D(_01526_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2364),
    .D(_01527_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2365),
    .D(_01528_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2366),
    .D(_01529_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2367),
    .D(_01530_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2368),
    .D(_01531_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2369),
    .D(_01532_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2370),
    .D(_01533_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2371),
    .D(_01534_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2372),
    .D(_01535_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2373),
    .D(_01536_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2374),
    .D(_01537_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2375),
    .D(_01538_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2376),
    .D(_01539_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2377),
    .D(_01540_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2378),
    .D(_01541_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2379),
    .D(_01542_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2380),
    .D(_01543_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2381),
    .D(_01544_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2382),
    .D(_01545_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2383),
    .D(_01546_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2384),
    .D(_01547_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2385),
    .D(_01548_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2386),
    .D(_01549_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2387),
    .D(_01550_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2388),
    .D(_01551_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2389),
    .D(_01552_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2390),
    .D(_01553_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2391),
    .D(_01554_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2392),
    .D(_01555_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2393),
    .D(_01556_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2394),
    .D(_01557_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2395),
    .D(_01558_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2396),
    .D(_01559_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2397),
    .D(_01560_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2398),
    .D(_01561_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2399),
    .D(_01562_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2400),
    .D(_01563_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2401),
    .D(_01564_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2402),
    .D(_01565_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2403),
    .D(_01566_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2404),
    .D(_01567_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2405),
    .D(_01568_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2406),
    .D(_01569_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2407),
    .D(_01570_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2408),
    .D(_01571_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2409),
    .D(_01572_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2410),
    .D(_01573_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2411),
    .D(_01574_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2412),
    .D(_01575_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2413),
    .D(_01576_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2414),
    .D(_01577_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2415),
    .D(_01578_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2416),
    .D(_01579_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2417),
    .D(_01580_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2418),
    .D(_01581_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2419),
    .D(_01582_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2420),
    .D(_01583_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2421),
    .D(_01584_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2422),
    .D(_01585_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2423),
    .D(_01586_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2424),
    .D(_01587_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2425),
    .D(_01588_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2426),
    .D(_01589_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2427),
    .D(_01590_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2428),
    .D(_01591_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2429),
    .D(_01592_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2430),
    .D(_01593_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2431),
    .D(_01594_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2432),
    .D(_01595_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2433),
    .D(_01596_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2434),
    .D(_01597_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2435),
    .D(_01598_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2436),
    .D(_01599_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2437),
    .D(_01600_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2438),
    .D(_01601_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2439),
    .D(_01602_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2440),
    .D(_01603_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2441),
    .D(_01604_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2442),
    .D(_01605_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2443),
    .D(_01606_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2444),
    .D(_01607_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2445),
    .D(_01608_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2446),
    .D(_01609_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2447),
    .D(_01610_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2448),
    .D(_01611_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2449),
    .D(_01612_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2450),
    .D(_01613_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2451),
    .D(_01614_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2452),
    .D(_01615_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2453),
    .D(_01616_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2454),
    .D(_01617_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2455),
    .D(_01618_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2456),
    .D(_01619_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2457),
    .D(_01620_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2458),
    .D(_01621_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2459),
    .D(_01622_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2460),
    .D(_01623_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2461),
    .D(_01624_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2462),
    .D(_01625_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2463),
    .D(_01626_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2464),
    .D(_01627_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2465),
    .D(_01628_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2466),
    .D(_01629_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2467),
    .D(_01630_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2468),
    .D(_01631_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2469),
    .D(_01632_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2470),
    .D(_01633_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2471),
    .D(_01634_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2472),
    .D(_01635_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2473),
    .D(_01636_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2474),
    .D(_01637_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2475),
    .D(_01638_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2476),
    .D(_01639_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2477),
    .D(_01640_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2478),
    .D(_01641_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2479),
    .D(_01642_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2480),
    .D(_01643_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2481),
    .D(_01644_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2482),
    .D(_01645_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2483),
    .D(_01646_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2484),
    .D(_01647_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2485),
    .D(_01648_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2486),
    .D(_01649_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2487),
    .D(_01650_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2488),
    .D(_01651_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2489),
    .D(_01652_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2490),
    .D(_01653_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2491),
    .D(_01654_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2492),
    .D(_01655_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2493),
    .D(_01656_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2494),
    .D(_01657_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2495),
    .D(_01658_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2496),
    .D(_01659_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2497),
    .D(_01660_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2498),
    .D(_01661_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2499),
    .D(_01662_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2500),
    .D(_01663_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2501),
    .D(_01664_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2502),
    .D(_01665_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2503),
    .D(_01666_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2504),
    .D(_01667_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2505),
    .D(_01668_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2506),
    .D(_01669_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2507),
    .D(_01670_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2508),
    .D(_01671_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2509),
    .D(_01672_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2510),
    .D(_01673_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2511),
    .D(_01674_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2512),
    .D(_01675_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2513),
    .D(_01676_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2514),
    .D(_01677_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2515),
    .D(_01678_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2516),
    .D(_01679_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2517),
    .D(_01680_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2518),
    .D(_01681_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2519),
    .D(_01682_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2520),
    .D(_01683_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2521),
    .D(_01684_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2522),
    .D(_01685_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2523),
    .D(_01686_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2524),
    .D(_01687_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2525),
    .D(_01688_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2526),
    .D(_01689_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2527),
    .D(_01690_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2528),
    .D(_01691_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2529),
    .D(_01692_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2530),
    .D(_01693_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2531),
    .D(_01694_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2532),
    .D(_01695_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2533),
    .D(_01696_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2534),
    .D(_01697_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2535),
    .D(_01698_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2536),
    .D(_01699_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2537),
    .D(_01700_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2538),
    .D(_01701_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2539),
    .D(_01702_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2540),
    .D(_01703_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2541),
    .D(_01704_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2542),
    .D(_01705_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2543),
    .D(_01706_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2544),
    .D(_01707_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2545),
    .D(_01708_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2546),
    .D(_01709_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2547),
    .D(_01710_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2548),
    .D(_01711_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2549),
    .D(_01712_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2550),
    .D(_01713_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2551),
    .D(_01714_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2552),
    .D(_01715_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2553),
    .D(_01716_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2554),
    .D(_01717_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2555),
    .D(_01718_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2556),
    .D(_01719_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2557),
    .D(_01720_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2558),
    .D(_01721_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2559),
    .D(_01722_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2560),
    .D(_01723_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2561),
    .D(_01724_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2562),
    .D(_01725_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2563),
    .D(_01726_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2564),
    .D(_01727_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2565),
    .D(_01728_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2566),
    .D(_01729_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2567),
    .D(_01730_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2568),
    .D(_01731_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2569),
    .D(_01732_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2570),
    .D(_01733_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2571),
    .D(_01734_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2572),
    .D(_01735_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2573),
    .D(_01736_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2574),
    .D(_01737_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2575),
    .D(_01738_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2576),
    .D(_01739_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2577),
    .D(_01740_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2578),
    .D(_01741_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2579),
    .D(_01742_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2580),
    .D(_01743_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2581),
    .D(_01744_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2582),
    .D(_01745_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2583),
    .D(_01746_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2584),
    .D(_01747_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2585),
    .D(_01748_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2586),
    .D(_01749_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2587),
    .D(_01750_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2588),
    .D(_01751_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2589),
    .D(_01752_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2590),
    .D(_01753_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2591),
    .D(_01754_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2592),
    .D(_01755_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2593),
    .D(_01756_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2594),
    .D(_01757_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2595),
    .D(_01758_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2596),
    .D(_01759_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2597),
    .D(_01760_),
    .Q_N(_13425_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2598),
    .D(_01761_),
    .Q_N(_13424_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2599),
    .D(_01762_),
    .Q_N(_13423_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2600),
    .D(_01763_),
    .Q_N(_13422_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2601),
    .D(_01764_),
    .Q_N(_13421_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2602),
    .D(_01765_),
    .Q_N(_13420_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2603),
    .D(_01766_),
    .Q_N(_13419_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2604),
    .D(_01767_),
    .Q_N(_13418_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2605),
    .D(_01768_),
    .Q_N(_13417_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2606),
    .D(_01769_),
    .Q_N(_13416_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2607),
    .D(_01770_),
    .Q_N(_13415_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2608),
    .D(_01771_),
    .Q_N(_13414_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2609),
    .D(_01772_),
    .Q_N(_13413_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2610),
    .D(_01773_),
    .Q_N(_13412_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2611),
    .D(_01774_),
    .Q_N(_13411_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2612),
    .D(_01775_),
    .Q_N(_13410_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2613),
    .D(_01776_),
    .Q_N(_13409_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2614),
    .D(_01777_),
    .Q_N(_13408_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2615),
    .D(_01778_),
    .Q_N(_13407_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2616),
    .D(_01779_),
    .Q_N(_13406_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2617),
    .D(_01780_),
    .Q_N(_13405_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2618),
    .D(_01781_),
    .Q_N(_13404_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2619),
    .D(_01782_),
    .Q_N(_13403_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2620),
    .D(_01783_),
    .Q_N(_13402_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2621),
    .D(_01784_),
    .Q_N(_13401_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2622),
    .D(_01785_),
    .Q_N(_13400_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2623),
    .D(_01786_),
    .Q_N(_13399_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2624),
    .D(_01787_),
    .Q_N(_13398_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2625),
    .D(_01788_),
    .Q_N(_13397_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2626),
    .D(_01789_),
    .Q_N(_13396_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2627),
    .D(_01790_),
    .Q_N(_13395_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2628),
    .D(_01791_),
    .Q_N(_13394_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2629),
    .D(_01792_),
    .Q_N(_13393_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2630),
    .D(_01793_),
    .Q_N(_13392_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2631),
    .D(_01794_),
    .Q_N(_13391_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2632),
    .D(_01795_),
    .Q_N(_13390_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2633),
    .D(_01796_),
    .Q_N(_13389_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2634),
    .D(_01797_),
    .Q_N(_13388_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2635),
    .D(_01798_),
    .Q_N(_13387_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2636),
    .D(_01799_),
    .Q_N(_13386_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2637),
    .D(_01800_),
    .Q_N(_13385_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2638),
    .D(_01801_),
    .Q_N(_13384_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2639),
    .D(_01802_),
    .Q_N(_13383_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2640),
    .D(_01803_),
    .Q_N(_13382_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2641),
    .D(_01804_),
    .Q_N(_13381_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2642),
    .D(_01805_),
    .Q_N(_13380_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2643),
    .D(_01806_),
    .Q_N(_13379_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2644),
    .D(_01807_),
    .Q_N(_13378_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2645),
    .D(_01808_),
    .Q_N(_13377_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2646),
    .D(_01809_),
    .Q_N(_13376_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2647),
    .D(_01810_),
    .Q_N(_13375_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2648),
    .D(_01811_),
    .Q_N(_13374_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2649),
    .D(_01812_),
    .Q_N(_13373_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2650),
    .D(_01813_),
    .Q_N(_13372_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2651),
    .D(_01814_),
    .Q_N(_13371_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2652),
    .D(_01815_),
    .Q_N(_13370_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2653),
    .D(_01816_),
    .Q_N(_13369_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2654),
    .D(_01817_),
    .Q_N(_13368_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2655),
    .D(_01818_),
    .Q_N(_13367_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2656),
    .D(_01819_),
    .Q_N(_13366_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2657),
    .D(_01820_),
    .Q_N(_13365_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2658),
    .D(_01821_),
    .Q_N(_13364_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2659),
    .D(_01822_),
    .Q_N(_13363_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2660),
    .D(_01823_),
    .Q_N(_13362_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2661),
    .D(_01824_),
    .Q_N(_13361_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2662),
    .D(_01825_),
    .Q_N(_13360_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2663),
    .D(_01826_),
    .Q_N(_13359_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2664),
    .D(_01827_),
    .Q_N(_13358_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2665),
    .D(_01828_),
    .Q_N(_13357_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2666),
    .D(_01829_),
    .Q_N(_13356_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2667),
    .D(_01830_),
    .Q_N(_13355_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2668),
    .D(_01831_),
    .Q_N(_13354_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2669),
    .D(_01832_),
    .Q_N(_13353_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2670),
    .D(_01833_),
    .Q_N(_13352_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2671),
    .D(_01834_),
    .Q_N(_13351_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2672),
    .D(_01835_),
    .Q_N(_13350_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2673),
    .D(_01836_),
    .Q_N(_13349_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2674),
    .D(_01837_),
    .Q_N(_13348_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2675),
    .D(_01838_),
    .Q_N(_13347_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2676),
    .D(_01839_),
    .Q_N(_13346_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2677),
    .D(_01840_),
    .Q_N(_13345_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2678),
    .D(_01841_),
    .Q_N(_13344_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2679),
    .D(_01842_),
    .Q_N(_13343_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2680),
    .D(_01843_),
    .Q_N(_13342_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2681),
    .D(_01844_),
    .Q_N(_13341_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2682),
    .D(_01845_),
    .Q_N(_13340_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2683),
    .D(_01846_),
    .Q_N(_13339_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2684),
    .D(_01847_),
    .Q_N(_13338_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2685),
    .D(_01848_),
    .Q_N(_13337_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2686),
    .D(_01849_),
    .Q_N(_13336_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2687),
    .D(_01850_),
    .Q_N(_13335_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2688),
    .D(_01851_),
    .Q_N(_13334_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2689),
    .D(_01852_),
    .Q_N(_13333_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2690),
    .D(_01853_),
    .Q_N(_13332_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2691),
    .D(_01854_),
    .Q_N(_13331_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2692),
    .D(_01855_),
    .Q_N(_13330_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2693),
    .D(_01856_),
    .Q_N(_13329_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2694),
    .D(_01857_),
    .Q_N(_13328_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2695),
    .D(_01858_),
    .Q_N(_13327_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2696),
    .D(_01859_),
    .Q_N(_13326_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2697),
    .D(_01860_),
    .Q_N(_13325_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2698),
    .D(_01861_),
    .Q_N(_13324_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2699),
    .D(_01862_),
    .Q_N(_13323_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2700),
    .D(_01863_),
    .Q_N(_13322_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2701),
    .D(_01864_),
    .Q_N(_13321_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2702),
    .D(_01865_),
    .Q_N(_13320_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2703),
    .D(_01866_),
    .Q_N(_13319_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2704),
    .D(_01867_),
    .Q_N(_13318_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2705),
    .D(_01868_),
    .Q_N(_13317_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2706),
    .D(_01869_),
    .Q_N(_13316_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2707),
    .D(_01870_),
    .Q_N(_13315_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2708),
    .D(_01871_),
    .Q_N(_13314_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2709),
    .D(_01872_),
    .Q_N(_13313_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2710),
    .D(_01873_),
    .Q_N(_13312_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2711),
    .D(_01874_),
    .Q_N(_13311_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2712),
    .D(_01875_),
    .Q_N(_13310_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2713),
    .D(_01876_),
    .Q_N(_13309_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2714),
    .D(_01877_),
    .Q_N(_13308_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2715),
    .D(_01878_),
    .Q_N(_13307_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2716),
    .D(_01879_),
    .Q_N(_13306_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2717),
    .D(_01880_),
    .Q_N(_13305_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2718),
    .D(_01881_),
    .Q_N(_13304_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2719),
    .D(_01882_),
    .Q_N(_13303_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2720),
    .D(_01883_),
    .Q_N(_13302_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2721),
    .D(_01884_),
    .Q_N(_13301_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2722),
    .D(_01885_),
    .Q_N(_13300_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2723),
    .D(_01886_),
    .Q_N(_13299_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2724),
    .D(_01887_),
    .Q_N(_13298_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2725),
    .D(_01888_),
    .Q_N(_13297_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2726),
    .D(_01889_),
    .Q_N(_13296_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2727),
    .D(_01890_),
    .Q_N(_13295_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2728),
    .D(_01891_),
    .Q_N(_13294_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2729),
    .D(_01892_),
    .Q_N(_13293_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2730),
    .D(_01893_),
    .Q_N(_13292_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2731),
    .D(_01894_),
    .Q_N(_13291_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2732),
    .D(_01895_),
    .Q_N(_13290_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2733),
    .D(_01896_),
    .Q_N(_13289_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2734),
    .D(_01897_),
    .Q_N(_13288_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2735),
    .D(_01898_),
    .Q_N(_13287_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2736),
    .D(_01899_),
    .Q_N(_13286_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2737),
    .D(_01900_),
    .Q_N(_13285_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2738),
    .D(_01901_),
    .Q_N(_13284_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2739),
    .D(_01902_),
    .Q_N(_13283_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2740),
    .D(_01903_),
    .Q_N(_13282_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2741),
    .D(_01904_),
    .Q_N(_13281_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2742),
    .D(_01905_),
    .Q_N(_13280_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2743),
    .D(_01906_),
    .Q_N(_13279_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2744),
    .D(_01907_),
    .Q_N(_13278_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2745),
    .D(_01908_),
    .Q_N(_13277_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2746),
    .D(_01909_),
    .Q_N(_13276_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2747),
    .D(_01910_),
    .Q_N(_13275_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2748),
    .D(_01911_),
    .Q_N(_13274_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2749),
    .D(_01912_),
    .Q_N(_13273_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2750),
    .D(_01913_),
    .Q_N(_13272_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2751),
    .D(_01914_),
    .Q_N(_13271_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2752),
    .D(_01915_),
    .Q_N(_13270_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2753),
    .D(_01916_),
    .Q_N(_13269_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2754),
    .D(_01917_),
    .Q_N(_13268_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2755),
    .D(_01918_),
    .Q_N(_13267_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2756),
    .D(_01919_),
    .Q_N(_13266_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2757),
    .D(_01920_),
    .Q_N(_13265_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2758),
    .D(_01921_),
    .Q_N(_13264_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2759),
    .D(_01922_),
    .Q_N(_13263_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2760),
    .D(_01923_),
    .Q_N(_13262_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2761),
    .D(_01924_),
    .Q_N(_13261_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2762),
    .D(_01925_),
    .Q_N(_13260_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2763),
    .D(_01926_),
    .Q_N(_13259_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2764),
    .D(_01927_),
    .Q_N(_13258_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2765),
    .D(_01928_),
    .Q_N(_13257_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2766),
    .D(_01929_),
    .Q_N(_13256_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2767),
    .D(_01930_),
    .Q_N(_13255_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2768),
    .D(_01931_),
    .Q_N(_13254_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2769),
    .D(_01932_),
    .Q_N(_13253_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2770),
    .D(_01933_),
    .Q_N(_13252_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2771),
    .D(_01934_),
    .Q_N(_13251_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2772),
    .D(_01935_),
    .Q_N(_13250_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2773),
    .D(_01936_),
    .Q_N(_13249_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2774),
    .D(_01937_),
    .Q_N(_13248_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2775),
    .D(_01938_),
    .Q_N(_13247_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2776),
    .D(_01939_),
    .Q_N(_13246_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2777),
    .D(_01940_),
    .Q_N(_13245_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2778),
    .D(_01941_),
    .Q_N(_13244_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2779),
    .D(_01942_),
    .Q_N(_13243_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2780),
    .D(_01943_),
    .Q_N(_13242_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2781),
    .D(_01944_),
    .Q_N(_13241_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2782),
    .D(_01945_),
    .Q_N(_13240_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2783),
    .D(_01946_),
    .Q_N(_13239_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2784),
    .D(_01947_),
    .Q_N(_13238_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2785),
    .D(_01948_),
    .Q_N(_13237_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2786),
    .D(_01949_),
    .Q_N(_13236_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2787),
    .D(_01950_),
    .Q_N(_13235_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2788),
    .D(_01951_),
    .Q_N(_13234_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2789),
    .D(_01952_),
    .Q_N(_13233_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2790),
    .D(_01953_),
    .Q_N(_13232_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2791),
    .D(_01954_),
    .Q_N(_13231_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2792),
    .D(_01955_),
    .Q_N(_13230_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2793),
    .D(_01956_),
    .Q_N(_13229_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2794),
    .D(_01957_),
    .Q_N(_13228_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2795),
    .D(_01958_),
    .Q_N(_13227_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2796),
    .D(_01959_),
    .Q_N(_13226_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2797),
    .D(_01960_),
    .Q_N(_13225_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2798),
    .D(_01961_),
    .Q_N(_13224_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2799),
    .D(_01962_),
    .Q_N(_13223_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2800),
    .D(_01963_),
    .Q_N(_13222_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2801),
    .D(_01964_),
    .Q_N(_13221_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2802),
    .D(_01965_),
    .Q_N(_13220_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2803),
    .D(_01966_),
    .Q_N(_13219_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2804),
    .D(_01967_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2805),
    .D(_01968_),
    .Q_N(_00110_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2806),
    .D(_01969_),
    .Q_N(_00119_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2807),
    .D(_01970_),
    .Q_N(_13218_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2808),
    .D(_01971_),
    .Q_N(_00138_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2809),
    .D(_01972_),
    .Q_N(_00150_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2810),
    .D(_01973_),
    .Q_N(_00162_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2811),
    .D(_01974_),
    .Q_N(_13217_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2812),
    .D(_01975_),
    .Q_N(_13216_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2813),
    .D(_01976_),
    .Q_N(_00187_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2814),
    .D(_01977_),
    .Q_N(_13215_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2815),
    .D(_01978_),
    .Q_N(_13214_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2816),
    .D(_01979_),
    .Q_N(_13213_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2817),
    .D(_01980_),
    .Q_N(_00186_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2818),
    .D(_01981_),
    .Q_N(_13212_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2819),
    .D(_01982_),
    .Q_N(_13211_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2820),
    .D(_01983_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2821),
    .D(_01984_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2822),
    .D(_01985_),
    .Q_N(_00116_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2823),
    .D(_01986_),
    .Q_N(_13210_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2824),
    .D(_01987_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2825),
    .D(_01988_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2826),
    .D(_01989_),
    .Q_N(_00158_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2827),
    .D(_01990_),
    .Q_N(_13209_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2828),
    .D(_01991_),
    .Q_N(_00137_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2829),
    .D(_01992_),
    .Q_N(_00149_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2830),
    .D(_01993_),
    .Q_N(_00161_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2831),
    .D(_01994_),
    .Q_N(_13208_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2832),
    .D(_01995_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2833),
    .D(_01996_),
    .Q_N(_00108_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2834),
    .D(_01997_),
    .Q_N(_00118_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2835),
    .D(_01998_),
    .Q_N(_13207_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2836),
    .D(_01999_),
    .Q_N(_00136_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2837),
    .D(_02000_),
    .Q_N(_00148_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2838),
    .D(_02001_),
    .Q_N(_00160_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2839),
    .D(_02002_),
    .Q_N(_13206_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2840),
    .D(_02003_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2841),
    .D(_02004_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2842),
    .D(_02005_),
    .Q_N(_00117_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2843),
    .D(_02006_),
    .Q_N(_13205_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2844),
    .D(_02007_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2845),
    .D(_02008_),
    .Q_N(_00147_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2846),
    .D(_02009_),
    .Q_N(_00159_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2847),
    .D(_02010_),
    .Q_N(_13204_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2848),
    .D(_02011_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net2849),
    .D(_02012_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2850),
    .D(_02013_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2851),
    .D(_02014_),
    .Q_N(_00205_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2852),
    .D(_02015_),
    .Q_N(_00207_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2853),
    .D(_02016_),
    .Q_N(_00213_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2854),
    .D(_02017_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2855),
    .D(_02018_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2856),
    .D(_02019_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2857),
    .D(_02020_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2858),
    .D(_02021_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2859),
    .D(_02022_),
    .Q_N(_00216_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2860),
    .D(_02023_),
    .Q_N(_00218_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2861),
    .D(_02024_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2862),
    .D(_02025_),
    .Q_N(_00220_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2863),
    .D(_02026_),
    .Q_N(_00210_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2864),
    .D(_02027_),
    .Q_N(_00212_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2865),
    .D(_02028_),
    .Q_N(_00173_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2866),
    .D(_02029_),
    .Q_N(_00175_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2867),
    .D(_02030_),
    .Q_N(_00177_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2868),
    .D(_02031_),
    .Q_N(_00206_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2869),
    .D(_02032_),
    .Q_N(_00208_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2870),
    .D(_02033_),
    .Q_N(_00214_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2871),
    .D(_02034_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2872),
    .D(_02035_),
    .Q_N(_00215_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2873),
    .D(_02036_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2874),
    .D(_02037_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2875),
    .D(_02038_),
    .Q_N(_00217_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2876),
    .D(_02039_),
    .Q_N(_00219_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2877),
    .D(_02040_),
    .Q_N(_00209_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2878),
    .D(_02041_),
    .Q_N(_00211_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2879),
    .D(_02042_),
    .Q_N(_00172_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2880),
    .D(_02043_),
    .Q_N(_00174_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2881),
    .D(_02044_),
    .Q_N(_00176_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2882),
    .D(_02045_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2883),
    .D(_02046_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2884),
    .D(_02047_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2885),
    .D(_02048_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2886),
    .D(_02049_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2887),
    .D(_02050_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2888),
    .D(_02051_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2889),
    .D(_02052_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2890),
    .D(_02053_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2891),
    .D(_02054_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2892),
    .D(_02055_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2893),
    .D(_02056_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2894),
    .D(_02057_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2895),
    .D(_02058_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2896),
    .D(_02059_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2897),
    .D(_02060_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2898),
    .D(_02061_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2899),
    .D(_02062_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2900),
    .D(_02063_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2901),
    .D(_02064_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2902),
    .D(_02065_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2903),
    .D(_02066_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2904),
    .D(_02067_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2905),
    .D(_02068_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2906),
    .D(_02069_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2907),
    .D(_02070_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2908),
    .D(_02071_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2909),
    .D(_02072_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2910),
    .D(_02073_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2911),
    .D(_02074_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2912),
    .D(_02075_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2913),
    .D(_02076_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2914),
    .D(_02077_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2915),
    .D(_02078_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2916),
    .D(_02079_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2917),
    .D(_02080_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2918),
    .D(_02081_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2919),
    .D(_02082_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2920),
    .D(_02083_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2921),
    .D(_02084_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2922),
    .D(_02085_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2923),
    .D(_02086_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2924),
    .D(_02087_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2925),
    .D(_02088_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2926),
    .D(_02089_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2927),
    .D(_02090_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2928),
    .D(_02091_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2929),
    .D(_02092_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2930),
    .D(_02093_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2931),
    .D(_02094_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2932),
    .D(_02095_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2933),
    .D(_02096_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2934),
    .D(_02097_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2935),
    .D(_02098_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2936),
    .D(_02099_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2937),
    .D(_02100_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2938),
    .D(_02101_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2939),
    .D(_02102_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2940),
    .D(_02103_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2941),
    .D(_02104_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2942),
    .D(_02105_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2943),
    .D(_02106_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2944),
    .D(_02107_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2945),
    .D(_02108_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2946),
    .D(_02109_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2947),
    .D(_02110_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2948),
    .D(_02111_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2949),
    .D(_02112_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2950),
    .D(_02113_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2951),
    .D(_02114_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2952),
    .D(_02115_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2953),
    .D(_02116_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2954),
    .D(_02117_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2955),
    .D(_02118_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2956),
    .D(_02119_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2957),
    .D(_02120_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2958),
    .D(_02121_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2959),
    .D(_02122_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2960),
    .D(_02123_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2961),
    .D(_02124_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2962),
    .D(_02125_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2963),
    .D(_02126_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2964),
    .D(_02127_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2965),
    .D(_02128_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2966),
    .D(_02129_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2967),
    .D(_02130_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2968),
    .D(_02131_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2969),
    .D(_02132_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2970),
    .D(_02133_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2971),
    .D(_02134_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2972),
    .D(_02135_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2973),
    .D(_02136_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2974),
    .D(_02137_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2975),
    .D(_02138_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2976),
    .D(_02139_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2977),
    .D(_02140_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2978),
    .D(_02141_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2979),
    .D(_02142_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2980),
    .D(_02143_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2981),
    .D(_02144_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2982),
    .D(_02145_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2983),
    .D(_02146_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2984),
    .D(_02147_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2985),
    .D(_02148_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2986),
    .D(_02149_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2987),
    .D(_02150_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2988),
    .D(_02151_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2989),
    .D(_02152_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2990),
    .D(_02153_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2991),
    .D(_02154_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2992),
    .D(_02155_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2993),
    .D(_02156_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2994),
    .D(_02157_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2995),
    .D(_02158_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2996),
    .D(_02159_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2997),
    .D(_02160_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2998),
    .D(_02161_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2999),
    .D(_02162_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3000),
    .D(_02163_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3001),
    .D(_02164_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3002),
    .D(_02165_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3003),
    .D(_02166_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3004),
    .D(_02167_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3005),
    .D(_02168_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3006),
    .D(_02169_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3007),
    .D(_02170_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3008),
    .D(_02171_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3009),
    .D(_02172_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3010),
    .D(_02173_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3011),
    .D(_02174_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3012),
    .D(_02175_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3013),
    .D(_02176_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3014),
    .D(_02177_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3015),
    .D(_02178_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3016),
    .D(_02179_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3017),
    .D(_02180_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3018),
    .D(_02181_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3019),
    .D(_02182_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3020),
    .D(_02183_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3021),
    .D(_02184_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3022),
    .D(_02185_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3023),
    .D(_02186_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3024),
    .D(_02187_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3025),
    .D(_02188_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3026),
    .D(_02189_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3027),
    .D(_02190_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3028),
    .D(_02191_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3029),
    .D(_02192_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3030),
    .D(_02193_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3031),
    .D(_02194_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3032),
    .D(_02195_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3033),
    .D(_02196_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3034),
    .D(_02197_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3035),
    .D(_02198_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3036),
    .D(_02199_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3037),
    .D(_02200_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3038),
    .D(_02201_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3039),
    .D(_02202_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3040),
    .D(_02203_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3041),
    .D(_02204_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3042),
    .D(_02205_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3043),
    .D(_02206_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3044),
    .D(_02207_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3045),
    .D(_02208_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3046),
    .D(_02209_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3047),
    .D(_02210_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3048),
    .D(_02211_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3049),
    .D(_02212_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3050),
    .D(_02213_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3051),
    .D(_02214_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3052),
    .D(_02215_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3053),
    .D(_02216_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3054),
    .D(_02217_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3055),
    .D(_02218_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3056),
    .D(_02219_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3057),
    .D(_02220_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3058),
    .D(_02221_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3059),
    .D(_02222_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3060),
    .D(_02223_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3061),
    .D(_02224_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3062),
    .D(_02225_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3063),
    .D(_02226_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3064),
    .D(_02227_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3065),
    .D(_02228_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3066),
    .D(_02229_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3067),
    .D(_02230_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3068),
    .D(_02231_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3069),
    .D(_02232_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3070),
    .D(_02233_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3071),
    .D(_02234_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3072),
    .D(_02235_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3073),
    .D(_02236_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3074),
    .D(_02237_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3075),
    .D(_02238_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3076),
    .D(_02239_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3077),
    .D(_02240_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3078),
    .D(_02241_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3079),
    .D(_02242_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3080),
    .D(_02243_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3081),
    .D(_02244_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3082),
    .D(_02245_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3083),
    .D(_02246_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3084),
    .D(_02247_),
    .Q_N(_12995_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3085),
    .D(_02248_),
    .Q_N(_12994_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3086),
    .D(_02249_),
    .Q_N(_12993_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3087),
    .D(_02250_),
    .Q_N(_12992_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3088),
    .D(_02251_),
    .Q_N(_12991_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3089),
    .D(_02252_),
    .Q_N(_12990_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3090),
    .D(_02253_),
    .Q_N(_12989_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3091),
    .D(_02254_),
    .Q_N(_12988_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3092),
    .D(_02255_),
    .Q_N(_12987_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3093),
    .D(_02256_),
    .Q_N(_12986_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3094),
    .D(_02257_),
    .Q_N(_12985_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3095),
    .D(_02258_),
    .Q_N(_12984_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3096),
    .D(_02259_),
    .Q_N(_12983_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3097),
    .D(_02260_),
    .Q_N(_12982_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3098),
    .D(_02261_),
    .Q_N(_12981_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3099),
    .D(_02262_),
    .Q_N(_12980_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3100),
    .D(_02263_),
    .Q_N(_12979_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3101),
    .D(_02264_),
    .Q_N(_12978_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3102),
    .D(_02265_),
    .Q_N(_12977_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3103),
    .D(_02266_),
    .Q_N(_12976_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3104),
    .D(_02267_),
    .Q_N(_12975_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3105),
    .D(_02268_),
    .Q_N(_12974_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3106),
    .D(_02269_),
    .Q_N(_00316_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3107),
    .D(_02270_),
    .Q_N(_12973_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3108),
    .D(_02271_),
    .Q_N(_00254_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3109),
    .D(_02272_),
    .Q_N(_12972_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3110),
    .D(_02273_),
    .Q_N(_12971_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3111),
    .D(_02274_),
    .Q_N(_12970_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3112),
    .D(_02275_),
    .Q_N(_12969_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3113),
    .D(_02276_),
    .Q_N(_12968_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3114),
    .D(_02277_),
    .Q_N(_12967_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3115),
    .D(_02278_),
    .Q_N(_12966_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3116),
    .D(_02279_),
    .Q_N(_12965_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3117),
    .D(_02280_),
    .Q_N(_12964_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3118),
    .D(_02281_),
    .Q_N(_12963_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3119),
    .D(_02282_),
    .Q_N(_12962_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3120),
    .D(_02283_),
    .Q_N(_12961_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3121),
    .D(_02284_),
    .Q_N(_12960_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3122),
    .D(_02285_),
    .Q_N(_12959_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3123),
    .D(_02286_),
    .Q_N(_12958_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3124),
    .D(_02287_),
    .Q_N(_12957_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3125),
    .D(_02288_),
    .Q_N(_12956_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3126),
    .D(_02289_),
    .Q_N(_12955_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3127),
    .D(_02290_),
    .Q_N(_12954_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3128),
    .D(_02291_),
    .Q_N(_12953_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3129),
    .D(_02292_),
    .Q_N(_12952_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3130),
    .D(_02293_),
    .Q_N(_12951_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3131),
    .D(_02294_),
    .Q_N(_12950_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3132),
    .D(_02295_),
    .Q_N(_12949_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3133),
    .D(_02296_),
    .Q_N(_12948_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3134),
    .D(_02297_),
    .Q_N(_12947_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3135),
    .D(_02298_),
    .Q_N(_12946_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3136),
    .D(_02299_),
    .Q_N(_12945_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3137),
    .D(_02300_),
    .Q_N(_12944_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3138),
    .D(_02301_),
    .Q_N(_12943_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3139),
    .D(_02302_),
    .Q_N(_12942_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3140),
    .D(_02303_),
    .Q_N(_12941_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3141),
    .D(_02304_),
    .Q_N(_12940_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3142),
    .D(_02305_),
    .Q_N(_12939_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3143),
    .D(_02306_),
    .Q_N(_12938_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3144),
    .D(_02307_),
    .Q_N(_12937_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3145),
    .D(_02308_),
    .Q_N(_12936_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3146),
    .D(_02309_),
    .Q_N(_12935_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3147),
    .D(_02310_),
    .Q_N(_12934_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3148),
    .D(_02311_),
    .Q_N(_12933_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3149),
    .D(_02312_),
    .Q_N(_12932_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3150),
    .D(_02313_),
    .Q_N(_12931_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3151),
    .D(_02314_),
    .Q_N(_12930_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3152),
    .D(_02315_),
    .Q_N(_12929_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3153),
    .D(_02316_),
    .Q_N(_12928_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3154),
    .D(_02317_),
    .Q_N(_12927_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3155),
    .D(_02318_),
    .Q_N(_12926_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3156),
    .D(_02319_),
    .Q_N(_12925_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3157),
    .D(_02320_),
    .Q_N(_12924_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3158),
    .D(_02321_),
    .Q_N(_12923_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3159),
    .D(_02322_),
    .Q_N(_12922_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3160),
    .D(_02323_),
    .Q_N(_12921_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3161),
    .D(_02324_),
    .Q_N(_12920_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3162),
    .D(_02325_),
    .Q_N(_12919_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3163),
    .D(_02326_),
    .Q_N(_12918_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3164),
    .D(_02327_),
    .Q_N(_12917_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3165),
    .D(_02328_),
    .Q_N(_12916_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3166),
    .D(_02329_),
    .Q_N(_12915_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3167),
    .D(_02330_),
    .Q_N(_12914_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3168),
    .D(_02331_),
    .Q_N(_12913_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3169),
    .D(_02332_),
    .Q_N(_12912_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3170),
    .D(_02333_),
    .Q_N(_12911_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3171),
    .D(_02334_),
    .Q_N(_12910_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3172),
    .D(_02335_),
    .Q_N(_12909_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3173),
    .D(_02336_),
    .Q_N(_12908_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3174),
    .D(_02337_),
    .Q_N(_12907_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3175),
    .D(_02338_),
    .Q_N(_12906_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3176),
    .D(_02339_),
    .Q_N(_12905_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3177),
    .D(_02340_),
    .Q_N(_12904_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3178),
    .D(_02341_),
    .Q_N(_12903_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3179),
    .D(_02342_),
    .Q_N(_12902_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3180),
    .D(_02343_),
    .Q_N(_12901_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3181),
    .D(_02344_),
    .Q_N(_12900_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3182),
    .D(_02345_),
    .Q_N(_12899_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3183),
    .D(_02346_),
    .Q_N(_12898_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3184),
    .D(_02347_),
    .Q_N(_12897_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3185),
    .D(_02348_),
    .Q_N(_12896_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3186),
    .D(_02349_),
    .Q_N(_12895_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3187),
    .D(_02350_),
    .Q_N(_12894_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3188),
    .D(_02351_),
    .Q_N(_12893_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3189),
    .D(_02352_),
    .Q_N(_12892_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3190),
    .D(_02353_),
    .Q_N(_12891_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3191),
    .D(_02354_),
    .Q_N(_12890_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3192),
    .D(_02355_),
    .Q_N(_12889_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3193),
    .D(_02356_),
    .Q_N(_12888_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3194),
    .D(_02357_),
    .Q_N(_12887_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3195),
    .D(_02358_),
    .Q_N(_12886_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3196),
    .D(_02359_),
    .Q_N(_12885_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3197),
    .D(_02360_),
    .Q_N(_12884_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3198),
    .D(_02361_),
    .Q_N(_12883_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3199),
    .D(_02362_),
    .Q_N(_12882_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3200),
    .D(_02363_),
    .Q_N(_12881_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3201),
    .D(_02364_),
    .Q_N(_12880_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3202),
    .D(_02365_),
    .Q_N(_12879_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3203),
    .D(_02366_),
    .Q_N(_12878_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3204),
    .D(_02367_),
    .Q_N(_12877_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3205),
    .D(_02368_),
    .Q_N(_12876_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3206),
    .D(_02369_),
    .Q_N(_12875_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3207),
    .D(_02370_),
    .Q_N(_12874_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3208),
    .D(_02371_),
    .Q_N(_12873_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3209),
    .D(_02372_),
    .Q_N(_12872_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3210),
    .D(_02373_),
    .Q_N(_12871_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3211),
    .D(_02374_),
    .Q_N(_12870_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3212),
    .D(_02375_),
    .Q_N(_12869_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3213),
    .D(_02376_),
    .Q_N(_12868_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3214),
    .D(_02377_),
    .Q_N(_12867_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3215),
    .D(_02378_),
    .Q_N(_12866_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3216),
    .D(_02379_),
    .Q_N(_12865_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3217),
    .D(_02380_),
    .Q_N(_12864_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3218),
    .D(_02381_),
    .Q_N(_12863_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net3219),
    .D(_02382_),
    .Q_N(_12862_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3220),
    .D(_02383_),
    .Q_N(_12861_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3221),
    .D(_02384_),
    .Q_N(_12860_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3222),
    .D(_02385_),
    .Q_N(_12859_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3223),
    .D(_02386_),
    .Q_N(_12858_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3224),
    .D(_02387_),
    .Q_N(_12857_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3225),
    .D(_02388_),
    .Q_N(_12856_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3226),
    .D(_02389_),
    .Q_N(_12855_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3227),
    .D(_02390_),
    .Q_N(_12854_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3228),
    .D(_02391_),
    .Q_N(_12853_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3229),
    .D(_02392_),
    .Q_N(_12852_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net3230),
    .D(_02393_),
    .Q_N(_12851_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3231),
    .D(_02394_),
    .Q_N(_12850_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3232),
    .D(_02395_),
    .Q_N(_12849_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3233),
    .D(_02396_),
    .Q_N(_12848_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3234),
    .D(_02397_),
    .Q_N(_12847_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3235),
    .D(_02398_),
    .Q_N(_12846_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net3236),
    .D(_02399_),
    .Q_N(_12845_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3237),
    .D(_02400_),
    .Q_N(_12844_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3238),
    .D(_02401_),
    .Q_N(_12843_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3239),
    .D(_02402_),
    .Q_N(_12842_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net3240),
    .D(_02403_),
    .Q_N(_12841_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3241),
    .D(_02404_),
    .Q_N(_12840_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3242),
    .D(_02405_),
    .Q_N(_12839_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3243),
    .D(_02406_),
    .Q_N(_12838_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3244),
    .D(_02407_),
    .Q_N(_12837_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3245),
    .D(_02408_),
    .Q_N(_12836_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3246),
    .D(_02409_),
    .Q_N(_12835_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net3247),
    .D(_02410_),
    .Q_N(_12834_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net3248),
    .D(_02411_),
    .Q_N(_12833_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3249),
    .D(_02412_),
    .Q_N(_12832_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3250),
    .D(_02413_),
    .Q_N(_12831_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3251),
    .D(_02414_),
    .Q_N(_12830_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3252),
    .D(_02415_),
    .Q_N(_12829_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3253),
    .D(_02416_),
    .Q_N(_12828_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net3254),
    .D(_02417_),
    .Q_N(_12827_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3255),
    .D(_02418_),
    .Q_N(_12826_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3256),
    .D(_02419_),
    .Q_N(_12825_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3257),
    .D(_02420_),
    .Q_N(_12824_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3258),
    .D(_02421_),
    .Q_N(_12823_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3259),
    .D(_02422_),
    .Q_N(_12822_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3260),
    .D(_02423_),
    .Q_N(_12821_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3261),
    .D(_02424_),
    .Q_N(_12820_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3262),
    .D(_02425_),
    .Q_N(_12819_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3263),
    .D(_02426_),
    .Q_N(_12818_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3264),
    .D(_02427_),
    .Q_N(_12817_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3265),
    .D(_02428_),
    .Q_N(_12816_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3266),
    .D(_02429_),
    .Q_N(_12815_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3267),
    .D(_02430_),
    .Q_N(_12814_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3268),
    .D(_02431_),
    .Q_N(_12813_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3269),
    .D(_02432_),
    .Q_N(_12812_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3270),
    .D(_02433_),
    .Q_N(_12811_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3271),
    .D(_02434_),
    .Q_N(_12810_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3272),
    .D(_02435_),
    .Q_N(_12809_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3273),
    .D(_02436_),
    .Q_N(_12808_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3274),
    .D(_02437_),
    .Q_N(_12807_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3275),
    .D(_02438_),
    .Q_N(_12806_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3276),
    .D(_02439_),
    .Q_N(_12805_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3277),
    .D(_02440_),
    .Q_N(_12804_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3278),
    .D(_02441_),
    .Q_N(_12803_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3279),
    .D(_02442_),
    .Q_N(_12802_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3280),
    .D(_02443_),
    .Q_N(_12801_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3281),
    .D(_02444_),
    .Q_N(_12800_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3282),
    .D(_02445_),
    .Q_N(_12799_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3283),
    .D(_02446_),
    .Q_N(_12798_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3284),
    .D(_02447_),
    .Q_N(_12797_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3285),
    .D(_02448_),
    .Q_N(_12796_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3286),
    .D(_02449_),
    .Q_N(_12795_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3287),
    .D(_02450_),
    .Q_N(_12794_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3288),
    .D(_02451_),
    .Q_N(_12793_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3289),
    .D(_02452_),
    .Q_N(_12792_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3290),
    .D(_02453_),
    .Q_N(_12791_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3291),
    .D(_02454_),
    .Q_N(_12790_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3292),
    .D(_02455_),
    .Q_N(_12789_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3293),
    .D(_02456_),
    .Q_N(_12788_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3294),
    .D(_02457_),
    .Q_N(_12787_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3295),
    .D(_02458_),
    .Q_N(_12786_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3296),
    .D(_02459_),
    .Q_N(_12785_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3297),
    .D(_02460_),
    .Q_N(_12784_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3298),
    .D(_02461_),
    .Q_N(_12783_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3299),
    .D(_02462_),
    .Q_N(_12782_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3300),
    .D(_02463_),
    .Q_N(_12781_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3301),
    .D(_02464_),
    .Q_N(_14773_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3302),
    .D(_00036_),
    .Q_N(_00286_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3303),
    .D(_00037_),
    .Q_N(_14774_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3304),
    .D(_00038_),
    .Q_N(_14775_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3305),
    .D(_00039_),
    .Q_N(_14776_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3306),
    .D(_00040_),
    .Q_N(_14777_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3307),
    .D(_00041_),
    .Q_N(_14778_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3308),
    .D(_00042_),
    .Q_N(_12780_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3309),
    .D(_02465_),
    .Q_N(_12779_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3310),
    .D(_02466_),
    .Q_N(_12778_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3311),
    .D(_02467_),
    .Q_N(_12777_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3312),
    .D(_02468_),
    .Q_N(_14779_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3313),
    .D(_00043_),
    .Q_N(_12776_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3314),
    .D(_02469_),
    .Q_N(_12775_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net3315),
    .D(_02470_),
    .Q_N(_12774_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3316),
    .D(_02471_),
    .Q_N(_12773_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3317),
    .D(_02472_),
    .Q_N(_12772_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3318),
    .D(_02473_),
    .Q_N(_12771_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3319),
    .D(_02474_),
    .Q_N(_12770_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3320),
    .D(_02475_),
    .Q_N(_12769_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3321),
    .D(_02476_),
    .Q_N(_12768_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3322),
    .D(_02477_),
    .Q_N(_12767_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3323),
    .D(_02478_),
    .Q_N(_14780_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3324),
    .D(_00044_),
    .Q_N(_12766_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3325),
    .D(_02479_),
    .Q_N(_12765_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3326),
    .D(_02480_),
    .Q_N(_14781_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3327),
    .D(_00045_),
    .Q_N(_14782_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3328),
    .D(_00046_),
    .Q_N(_14783_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3329),
    .D(_00047_),
    .Q_N(_14784_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3330),
    .D(_00048_),
    .Q_N(_14785_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3331),
    .D(_00049_),
    .Q_N(_14786_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3332),
    .D(_00050_),
    .Q_N(_14787_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3333),
    .D(_00051_),
    .Q_N(_12764_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3334),
    .D(_02481_),
    .Q_N(_12763_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3335),
    .D(_02482_),
    .Q_N(_12762_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3336),
    .D(_02483_),
    .Q_N(_12761_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3337),
    .D(_02484_),
    .Q_N(_12760_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3338),
    .D(_02485_),
    .Q_N(_12759_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3339),
    .D(_02486_),
    .Q_N(_12758_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3340),
    .D(_02487_),
    .Q_N(_14788_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3341),
    .D(_00055_),
    .Q_N(_00285_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3342),
    .D(_00056_),
    .Q_N(_14789_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3343),
    .D(_00057_),
    .Q_N(_14790_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3344),
    .D(_00058_),
    .Q_N(_14791_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3345),
    .D(_00059_),
    .Q_N(_14792_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3346),
    .D(_00060_),
    .Q_N(_14793_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3347),
    .D(_00061_),
    .Q_N(_14794_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3348),
    .D(_00062_),
    .Q_N(_14795_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3349),
    .D(_00063_),
    .Q_N(_14796_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3350),
    .D(_00064_),
    .Q_N(_14797_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3351),
    .D(_00065_),
    .Q_N(_14798_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3352),
    .D(_00066_),
    .Q_N(_14799_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3353),
    .D(_00067_),
    .Q_N(_14800_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3354),
    .D(_00068_),
    .Q_N(_14801_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3355),
    .D(_00069_),
    .Q_N(_14802_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3356),
    .D(_00070_),
    .Q_N(_14803_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3357),
    .D(_00071_),
    .Q_N(_14804_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3358),
    .D(_00072_),
    .Q_N(_14805_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3359),
    .D(_00073_),
    .Q_N(_14806_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3360),
    .D(_00074_),
    .Q_N(_14807_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3361),
    .D(_00075_),
    .Q_N(_14808_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3362),
    .D(_00076_),
    .Q_N(_14809_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3363),
    .D(_00077_),
    .Q_N(_14810_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3364),
    .D(_00078_),
    .Q_N(_12757_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3365),
    .D(_02488_),
    .Q_N(_12756_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3366),
    .D(_02489_),
    .Q_N(_12755_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net3367),
    .D(_02490_),
    .Q_N(_12754_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3368),
    .D(_02491_),
    .Q_N(_12753_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3369),
    .D(_02492_),
    .Q_N(_12752_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net3370),
    .D(_02493_),
    .Q_N(_12751_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net3371),
    .D(_02494_),
    .Q_N(_12750_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3372),
    .D(_02495_),
    .Q_N(_12749_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3373),
    .D(_02496_),
    .Q_N(_12748_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3374),
    .D(_02497_),
    .Q_N(_12747_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3375),
    .D(_02498_),
    .Q_N(_12746_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3376),
    .D(_02499_),
    .Q_N(_12745_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3377),
    .D(_02500_),
    .Q_N(_12744_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3378),
    .D(_02501_),
    .Q_N(_12743_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3379),
    .D(_02502_),
    .Q_N(_12742_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3380),
    .D(_02503_),
    .Q_N(_12741_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3381),
    .D(_02504_),
    .Q_N(_12740_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net3382),
    .D(_02505_),
    .Q_N(_12739_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3383),
    .D(_02506_),
    .Q_N(_12738_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3384),
    .D(_02507_),
    .Q_N(_12737_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3385),
    .D(_02508_),
    .Q_N(_12736_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3386),
    .D(_02509_),
    .Q_N(_12735_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3387),
    .D(_02510_),
    .Q_N(_12734_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net3388),
    .D(_02511_),
    .Q_N(_12733_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3389),
    .D(_02512_),
    .Q_N(_00183_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3390),
    .D(_02513_),
    .Q_N(_12732_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3391),
    .D(_02514_),
    .Q_N(_00184_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3392),
    .D(_02515_),
    .Q_N(_12731_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net3393),
    .D(_02516_),
    .Q_N(_00252_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3394),
    .D(_02517_),
    .Q_N(_12730_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3395),
    .D(_02518_),
    .Q_N(_12729_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3396),
    .D(_02519_),
    .Q_N(_12728_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net3397),
    .D(_02520_),
    .Q_N(_12727_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3398),
    .D(_02521_),
    .Q_N(_12726_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3399),
    .D(_02522_),
    .Q_N(_12725_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3400),
    .D(_02523_),
    .Q_N(_12724_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3401),
    .D(_02524_),
    .Q_N(_12723_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3402),
    .D(_02525_),
    .Q_N(_12722_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3403),
    .D(_02526_),
    .Q_N(_12721_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3404),
    .D(_02527_),
    .Q_N(_12720_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3405),
    .D(_02528_),
    .Q_N(_12719_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net3406),
    .D(_02529_),
    .Q_N(_12718_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3407),
    .D(_02530_),
    .Q_N(_12717_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3408),
    .D(_02531_),
    .Q_N(_12716_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3409),
    .D(_02532_),
    .Q_N(_12715_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3410),
    .D(_02533_),
    .Q_N(_12714_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3411),
    .D(_02534_),
    .Q_N(_12713_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3412),
    .D(_02535_),
    .Q_N(_12712_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net3413),
    .D(_02536_),
    .Q_N(_12711_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3414),
    .D(_02537_),
    .Q_N(_12710_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net3415),
    .D(_02538_),
    .Q_N(_12709_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3416),
    .D(_02539_),
    .Q_N(_12708_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3417),
    .D(_02540_),
    .Q_N(_14811_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3418),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14812_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3419),
    .D(_00021_),
    .Q_N(_00277_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3420),
    .D(_00008_),
    .Q_N(_14813_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3421),
    .D(_00022_),
    .Q_N(_14814_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3422),
    .D(_00023_),
    .Q_N(_14815_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3423),
    .D(_00009_),
    .Q_N(_14816_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net3424),
    .D(_00024_),
    .Q_N(_14817_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3425),
    .D(_00010_),
    .Q_N(_14818_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3426),
    .D(_00025_),
    .Q_N(_14819_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3427),
    .D(_00026_),
    .Q_N(_14820_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net3428),
    .D(_00001_),
    .Q_N(_14821_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net3429),
    .D(_00027_),
    .Q_N(_14822_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net3430),
    .D(_00002_),
    .Q_N(_14823_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net3431),
    .D(_00028_),
    .Q_N(_14824_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3432),
    .D(_00003_),
    .Q_N(_14825_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3433),
    .D(_00004_),
    .Q_N(_14826_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net3434),
    .D(_00005_),
    .Q_N(_14827_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3435),
    .D(_00006_),
    .Q_N(_00185_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3436),
    .D(_00007_),
    .Q_N(_12707_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net3437),
    .D(_02541_),
    .Q_N(_12706_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net3438),
    .D(_02542_),
    .Q_N(_12705_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3439),
    .D(_02543_),
    .Q_N(_12704_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3440),
    .D(_02544_),
    .Q_N(_12703_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3441),
    .D(_02545_),
    .Q_N(_12702_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net3442),
    .D(_02546_),
    .Q_N(_14828_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net3443),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_14829_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3444),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00253_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3445),
    .D(_02547_),
    .Q_N(_12701_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3446),
    .D(_02548_),
    .Q_N(_12700_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3447),
    .D(_02549_),
    .Q_N(_12699_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3448),
    .D(_02550_),
    .Q_N(_12698_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3449),
    .D(_02551_),
    .Q_N(_00314_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3450),
    .D(_02552_),
    .Q_N(_00095_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3451),
    .D(_02553_),
    .Q_N(_00105_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3452),
    .D(_02554_),
    .Q_N(_00115_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3453),
    .D(_02555_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3454),
    .D(_02556_),
    .Q_N(_00133_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3455),
    .D(_02557_),
    .Q_N(_00145_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3456),
    .D(_02558_),
    .Q_N(_00157_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3457),
    .D(_02559_),
    .Q_N(_00313_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3458),
    .D(_02560_),
    .Q_N(_00094_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3459),
    .D(_02561_),
    .Q_N(_00104_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3460),
    .D(_02562_),
    .Q_N(_00114_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3461),
    .D(_02563_),
    .Q_N(_00125_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3462),
    .D(_02564_),
    .Q_N(_00132_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3463),
    .D(_02565_),
    .Q_N(_00144_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3464),
    .D(_02566_),
    .Q_N(_00156_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3465),
    .D(_02567_),
    .Q_N(_12697_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3466),
    .D(_02568_),
    .Q_N(_12696_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3467),
    .D(_02569_),
    .Q_N(_12695_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3468),
    .D(_02570_),
    .Q_N(_12694_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3469),
    .D(_02571_),
    .Q_N(_12693_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3470),
    .D(_02572_),
    .Q_N(_12692_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3471),
    .D(_02573_),
    .Q_N(_12691_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3472),
    .D(_02574_),
    .Q_N(_12690_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3473),
    .D(_02575_),
    .Q_N(_12689_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3474),
    .D(_02576_),
    .Q_N(_12688_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3475),
    .D(_02577_),
    .Q_N(_12687_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3476),
    .D(_02578_),
    .Q_N(_12686_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3477),
    .D(_02579_),
    .Q_N(_12685_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3478),
    .D(_02580_),
    .Q_N(_12684_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3479),
    .D(_02581_),
    .Q_N(_12683_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3480),
    .D(_02582_),
    .Q_N(_12682_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3481),
    .D(_02583_),
    .Q_N(_12681_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3482),
    .D(_02584_),
    .Q_N(_12680_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3483),
    .D(_02585_),
    .Q_N(_12679_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3484),
    .D(_02586_),
    .Q_N(_12678_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3485),
    .D(_02587_),
    .Q_N(_12677_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3486),
    .D(_02588_),
    .Q_N(_12676_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3487),
    .D(_02589_),
    .Q_N(_12675_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3488),
    .D(_02590_),
    .Q_N(_12674_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3489),
    .D(_02591_),
    .Q_N(_12673_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3490),
    .D(_02592_),
    .Q_N(_12672_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3491),
    .D(_02593_),
    .Q_N(_00222_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3492),
    .D(_02594_),
    .Q_N(_12671_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3493),
    .D(_02595_),
    .Q_N(_00224_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3494),
    .D(_02596_),
    .Q_N(_12670_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3495),
    .D(_02597_),
    .Q_N(_12669_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3496),
    .D(_02598_),
    .Q_N(_12668_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3497),
    .D(_02599_),
    .Q_N(_12667_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3498),
    .D(_02600_),
    .Q_N(_12666_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3499),
    .D(_02601_),
    .Q_N(_12665_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3500),
    .D(_02602_),
    .Q_N(_12664_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3501),
    .D(_02603_),
    .Q_N(_12663_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3502),
    .D(_02604_),
    .Q_N(_12662_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3503),
    .D(_02605_),
    .Q_N(_12661_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net3504),
    .D(_02606_),
    .Q_N(_12660_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3505),
    .D(_02607_),
    .Q_N(_12659_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3506),
    .D(_02608_),
    .Q_N(_12658_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3507),
    .D(_02609_),
    .Q_N(_12657_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3508),
    .D(_02610_),
    .Q_N(_00221_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3509),
    .D(_02611_),
    .Q_N(_12656_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3510),
    .D(_02612_),
    .Q_N(_12655_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3511),
    .D(_02613_),
    .Q_N(_00282_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3512),
    .D(_02614_),
    .Q_N(_00283_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3513),
    .D(_02615_),
    .Q_N(_14830_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3514),
    .D(_00029_),
    .Q_N(_14831_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3515),
    .D(_00030_),
    .Q_N(_00225_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3516),
    .D(_00031_),
    .Q_N(_14832_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3517),
    .D(_00032_),
    .Q_N(_14833_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3518),
    .D(_00033_),
    .Q_N(_00278_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3519),
    .D(_00034_),
    .Q_N(_14834_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3520),
    .D(_00035_),
    .Q_N(_00226_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3521),
    .D(_02616_),
    .Q_N(_12654_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3522),
    .D(_02617_),
    .Q_N(_12653_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3523),
    .D(_02618_),
    .Q_N(_12652_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3524),
    .D(_02619_),
    .Q_N(_12651_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3525),
    .D(_02620_),
    .Q_N(_12650_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3526),
    .D(_02621_),
    .Q_N(_12649_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3527),
    .D(_02622_),
    .Q_N(_12648_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3528),
    .D(_02623_),
    .Q_N(_12647_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3529),
    .D(_02624_),
    .Q_N(_00284_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3530),
    .D(_02625_),
    .Q_N(_12646_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3531),
    .D(_02626_),
    .Q_N(_12645_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3532),
    .D(_02627_),
    .Q_N(_12644_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3533),
    .D(_02628_),
    .Q_N(_12643_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3534),
    .D(_02629_),
    .Q_N(_12642_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3535),
    .D(_02630_),
    .Q_N(_12641_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3536),
    .D(_02631_),
    .Q_N(_14835_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3537),
    .D(_00079_),
    .Q_N(_00279_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3538),
    .D(_00080_),
    .Q_N(_14836_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3539),
    .D(_00081_),
    .Q_N(_14837_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3540),
    .D(_00082_),
    .Q_N(_14838_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3541),
    .D(_00083_),
    .Q_N(_14839_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3542),
    .D(_00084_),
    .Q_N(_14840_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3543),
    .D(_00085_),
    .Q_N(_14841_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3544),
    .D(_00086_),
    .Q_N(_14842_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3545),
    .D(_00087_),
    .Q_N(_14843_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3546),
    .D(_00088_),
    .Q_N(_14844_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3547),
    .D(_00089_),
    .Q_N(_14845_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3548),
    .D(_00090_),
    .Q_N(_12640_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3549),
    .D(_02632_),
    .Q_N(_12639_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3550),
    .D(_02633_),
    .Q_N(_12638_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3551),
    .D(_02634_),
    .Q_N(_12637_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3552),
    .D(_02635_),
    .Q_N(_12636_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3553),
    .D(_02636_),
    .Q_N(_12635_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3554),
    .D(_02637_),
    .Q_N(_12634_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3555),
    .D(_02638_),
    .Q_N(_12633_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3556),
    .D(_02639_),
    .Q_N(_12632_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3557),
    .D(_02640_),
    .Q_N(_12631_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3558),
    .D(_02641_),
    .Q_N(_12630_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3559),
    .D(_02642_),
    .Q_N(_12629_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3560),
    .D(_02643_),
    .Q_N(_12628_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3561),
    .D(_02644_),
    .Q_N(_12627_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3562),
    .D(_02645_),
    .Q_N(_12626_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3563),
    .D(_02646_),
    .Q_N(_12625_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3564),
    .D(_02647_),
    .Q_N(_12624_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3565),
    .D(_02648_),
    .Q_N(_12623_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3566),
    .D(_02649_),
    .Q_N(_12622_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3567),
    .D(_02650_),
    .Q_N(_12621_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3568),
    .D(_02651_),
    .Q_N(_12620_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3569),
    .D(_02652_),
    .Q_N(_12619_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3570),
    .D(_02653_),
    .Q_N(_12618_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3571),
    .D(_02654_),
    .Q_N(_12617_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3572),
    .D(_02655_),
    .Q_N(_12616_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3573),
    .D(_02656_),
    .Q_N(_12615_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3574),
    .D(_02657_),
    .Q_N(_12614_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3575),
    .D(_02658_),
    .Q_N(_12613_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3576),
    .D(_02659_),
    .Q_N(_12612_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3577),
    .D(_02660_),
    .Q_N(_12611_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3578),
    .D(_02661_),
    .Q_N(_12610_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3579),
    .D(_02662_),
    .Q_N(_12609_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3580),
    .D(_02663_),
    .Q_N(_12608_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3581),
    .D(_02664_),
    .Q_N(_12607_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3582),
    .D(_02665_),
    .Q_N(_12606_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3583),
    .D(_02666_),
    .Q_N(_14846_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3584),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12605_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3585),
    .D(_02667_),
    .Q_N(_12604_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3586),
    .D(_02668_),
    .Q_N(_12603_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3587),
    .D(_02669_),
    .Q_N(_12602_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3588),
    .D(_02670_),
    .Q_N(_12601_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3589),
    .D(_02671_),
    .Q_N(_12600_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3590),
    .D(_02672_),
    .Q_N(_12599_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3591),
    .D(_02673_),
    .Q_N(_12598_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3592),
    .D(_02674_),
    .Q_N(_12597_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3593),
    .D(_02675_),
    .Q_N(_12596_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3594),
    .D(_02676_),
    .Q_N(_12595_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3595),
    .D(_02677_),
    .Q_N(_00280_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3596),
    .D(_02678_),
    .Q_N(_12594_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3597),
    .D(_02679_),
    .Q_N(_12593_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3598),
    .D(_02680_),
    .Q_N(_12592_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3599),
    .D(_02681_),
    .Q_N(_12591_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3600),
    .D(_02682_),
    .Q_N(_12590_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3601),
    .D(_02683_),
    .Q_N(_14847_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3602),
    .D(_00000_),
    .Q_N(_12589_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_06607_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_03744_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_07120_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_06875_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_04992_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_04797_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_04137_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02826_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02787_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02767_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02759_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02706_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_12576_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_12556_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_12548_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_12489_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_12455_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_12435_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12427_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12344_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12324_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12316_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12259_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12225_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12205_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12197_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12138_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12102_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12080_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12071_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12012_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_11966_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_11936_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_11923_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_11659_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_07195_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_12383_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_11881_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_11810_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_09870_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_09859_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_09857_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_09698_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_09192_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_07288_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_07287_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_07284_),
    .X(net73));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(_06593_));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_06587_));
 sg13g2_buf_2 fanout76 (.A(_04223_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_11324_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_09966_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_09955_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_09191_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_07773_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_07283_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04127_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_04090_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_04024_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_03070_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_11394_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_11329_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_11323_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_09965_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_09762_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_08928_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_06757_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_06686_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_06646_),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_06590_));
 sg13g2_buf_2 fanout97 (.A(_04089_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_03220_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_11369_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_11328_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_10001_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_09971_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_09950_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_09899_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_09898_),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_09768_));
 sg13g2_buf_2 fanout107 (.A(_09679_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_08997_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_08893_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_08845_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_08841_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_04328_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_04257_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_04154_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_04150_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_04088_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04082_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04054_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_03485_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_03474_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_02987_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_10722_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_09957_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_09949_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_08251_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_07509_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_05340_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_05117_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_04253_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_04174_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04165_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04076_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04041_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04037_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04028_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_03654_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_03608_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_03592_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_03591_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03578_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03461_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03456_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_03111_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_02992_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02975_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_02962_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_09730_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_07600_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_07530_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_07521_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_05413_),
    .X(net151));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_05252_));
 sg13g2_buf_2 fanout153 (.A(_04983_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04796_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04252_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04249_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_03603_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_03476_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_03460_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_02976_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_02963_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_11628_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_11623_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_09729_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_08991_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_08249_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_07692_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_07674_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_07670_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_07562_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_07522_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_07502_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(_07166_));
 sg13g2_buf_2 fanout174 (.A(_04182_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_04152_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_04109_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_03955_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_03549_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_03546_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_03498_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_03186_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_11572_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_11499_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_11488_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_11318_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_11286_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_11271_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_11206_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_09731_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_08916_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_08355_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_07723_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_07700_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_07673_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_05992_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_05926_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_05882_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_03559_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_03505_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_03491_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_03453_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_03137_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_03063_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_03031_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_03014_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_02981_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_02974_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_11564_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_11393_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_11295_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_11095_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_11073_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_09783_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_07662_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_06485_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_06478_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_06461_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_06459_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_06458_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_06362_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_06361_),
    .X(net221));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(_05969_));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_05953_));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(_05950_));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_05910_));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(_05905_));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_05900_));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(_05853_));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(_05848_));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_05825_));
 sg13g2_buf_2 fanout231 (.A(_05179_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_04988_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_04318_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_04025_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_03457_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_03452_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_03057_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_02991_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_02988_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_02967_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_02964_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_11442_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_11440_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_11332_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_11316_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_11139_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_10518_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_09782_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_08990_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_06568_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_06566_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_06565_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_06524_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_06522_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_06521_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_06457_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_06439_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_06437_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_06436_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_06225_),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_06213_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_06207_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_06201_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_06195_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_06189_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_06183_));
 sg13g2_buf_2 fanout267 (.A(_06176_),
    .X(net267));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_06170_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_06164_));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_06158_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_06151_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_06145_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_06139_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_06123_));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_06116_));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(_06103_));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_06097_));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_06090_));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_06084_));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(_06078_));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_06072_));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(_06065_));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_06058_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_06047_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_06039_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_06025_));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_06018_));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_06012_));
 sg13g2_buf_2 fanout289 (.A(_06003_),
    .X(net289));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(_05989_));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_05985_));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(_05980_));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_05974_));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_05965_));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_05962_));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_05959_));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(_05956_));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(_05941_));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(_05933_));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(_05922_));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_05916_));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(_05913_));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(_05897_));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(_05891_));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(_05873_));
 sg13g2_buf_4 fanout306 (.X(net306),
    .A(_05863_));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_05859_));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(_05841_));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(_05832_));
 sg13g2_buf_2 fanout310 (.A(_05307_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_04501_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_03798_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_03451_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_03399_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_02979_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_11402_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_11383_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_11368_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_11291_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_11119_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_11037_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_11003_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_11000_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_09694_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_06564_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_06520_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_06435_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_06219_),
    .X(net328));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_06133_));
 sg13g2_buf_2 fanout330 (.A(_05907_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_05834_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_05083_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_04875_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_03770_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_03398_),
    .X(net335));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_02910_));
 sg13g2_buf_2 fanout337 (.A(_02909_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_11543_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_11389_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_11313_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_10883_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_09780_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_09724_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_09249_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_09141_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_08969_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_08838_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_08401_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_08210_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_06546_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_06544_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_06543_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_06502_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_06500_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_06499_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_06420_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_06413_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_06298_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_06297_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_05154_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_05104_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_04951_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_04948_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_04824_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_04808_),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_03397_));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_02960_));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(_02959_));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(_02955_));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(_02946_));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_02945_));
 sg13g2_buf_2 fanout372 (.A(_02888_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_10798_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_10071_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_09963_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_09316_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_09140_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_08908_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_08837_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_08564_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_08543_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_08522_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_08498_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_08477_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_08426_),
    .X(net385));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(_08341_));
 sg13g2_buf_2 fanout387 (.A(_08212_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_08209_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_06876_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_06542_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_06498_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_06009_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_05856_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_05826_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_05155_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_05110_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_04928_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_04921_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_04894_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_04891_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_04870_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_04854_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_04807_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_03759_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_03396_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_03395_),
    .X(net406));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(_02956_));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(_02952_));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(_02948_));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(_02947_));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(_02931_));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_02929_));
 sg13g2_buf_2 fanout413 (.A(_02900_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_02896_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_02893_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_02887_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_02828_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_02708_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_12261_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_11902_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_11899_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_11895_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_11888_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_11728_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_11182_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_10915_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_10891_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_10070_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_09962_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_09631_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_09609_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_09586_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_09562_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_09537_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_09515_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_09493_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_09467_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_09444_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_09342_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_08911_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_08909_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_08650_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_08628_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_08607_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_08585_),
    .X(net445));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(_08346_));
 sg13g2_buf_2 fanout447 (.A(_08214_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_08211_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_08208_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_08201_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_08173_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_08158_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_06884_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_06231_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_06229_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_06130_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_06054_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_05107_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_05082_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_05081_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_04887_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_04860_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_04823_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_04799_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_04740_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_04737_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_03695_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_03415_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_03394_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_03389_),
    .X(net470));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(_02953_));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_02939_));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_02937_));
 sg13g2_buf_2 fanout474 (.A(_02906_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_02903_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_02899_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_02895_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_02892_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_02756_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_12545_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_12492_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_12194_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_12017_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_11885_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_11877_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_11816_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_11806_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_11764_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_11719_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_11049_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_10221_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_10095_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_09274_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_09262_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(\cpu.ex.c_mult_off[0] ),
    .X(net495));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(_09094_));
 sg13g2_buf_2 fanout497 (.A(_09024_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_08450_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_08217_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_08207_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_08200_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_08189_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_08178_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_08172_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_08166_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_08157_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_06125_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_06049_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_05918_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_05855_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_05833_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_04881_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_04842_),
    .X(net513));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(_04802_));
 sg13g2_buf_2 fanout515 (.A(_04742_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_04730_),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(_04727_));
 sg13g2_buf_2 fanout518 (.A(_03808_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_03755_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_03696_),
    .X(net520));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_03440_));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(_03432_));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_03420_));
 sg13g2_buf_2 fanout524 (.A(_03416_),
    .X(net524));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(_03414_));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_03403_));
 sg13g2_buf_2 fanout527 (.A(_03391_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_03388_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_03387_),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(_03385_));
 sg13g2_buf_2 fanout531 (.A(_02905_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_02902_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_12544_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_12424_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_12140_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_11918_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_11718_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_11335_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_11121_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_10220_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_10106_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_10066_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_09976_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_09944_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_09346_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_09281_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_09273_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_09268_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_09261_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_09258_),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_09119_));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_09093_));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(_08899_));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_08894_));
 sg13g2_buf_2 fanout555 (.A(_08206_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_08199_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_08188_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_08177_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_08171_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_08165_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_07872_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_07801_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_07772_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_07737_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_07713_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_07685_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_07647_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_07613_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_07565_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_07487_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_07476_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_07415_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_06043_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_05942_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_05923_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_05906_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_05874_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_05860_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_05766_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_05098_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_04822_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_04116_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_03754_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_03710_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_03709_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_03704_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_03690_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_03689_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_03439_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_03431_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_03425_),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(_03423_));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(_03408_));
 sg13g2_buf_2 fanout594 (.A(_03390_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_03386_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_02928_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_12423_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_12378_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_12313_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_12068_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_11762_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_11753_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_11717_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_11373_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_11050_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_10725_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_10224_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_09975_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_09943_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_09710_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_09313_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_09286_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_09280_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_09267_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_09257_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_09213_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_09187_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_09184_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_09092_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_09086_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_08195_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_08183_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_08176_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_08170_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_08164_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_07391_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_06869_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_06684_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_06655_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_06128_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_06126_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_06120_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_06052_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_06050_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_05176_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_04821_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_03703_),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(_03699_));
 sg13g2_buf_2 fanout639 (.A(_03697_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_03693_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_03417_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_03393_),
    .X(net642));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(_02927_));
 sg13g2_buf_2 fanout644 (.A(_11727_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_11663_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_11372_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_11153_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_11062_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_11056_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_11052_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_10859_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_10420_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_10388_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_10320_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_10281_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_10275_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_10248_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_10245_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_10244_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_10235_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_10153_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_10144_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_10137_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_10133_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_10113_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_09959_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_09952_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_09942_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_09815_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_09814_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_09675_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_09478_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_09290_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_09245_),
    .X(net674));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_09231_));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_09228_));
 sg13g2_buf_2 fanout677 (.A(_09219_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_09212_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_09185_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_09129_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_09091_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_09085_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_08832_),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(_08516_),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(_08460_),
    .X(net685));
 sg13g2_buf_8 fanout686 (.A(_08392_),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(_08370_),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(_08363_));
 sg13g2_buf_2 fanout689 (.A(_08316_),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(_08231_));
 sg13g2_buf_2 fanout691 (.A(_08226_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_08194_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_08182_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_08163_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_07185_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_06685_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_06683_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_06178_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_06109_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_06108_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_06107_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_06105_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_06031_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_06030_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_06029_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_06027_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_05917_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_05854_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_05779_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_04984_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_04792_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_03702_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_03698_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_03692_),
    .X(net714));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_03428_));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_03427_));
 sg13g2_buf_2 fanout717 (.A(_03392_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_03378_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_03217_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_02941_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_02940_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_02938_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_02933_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_02932_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_02930_),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(_02920_));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_02918_));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_02916_));
 sg13g2_buf_2 fanout729 (.A(_02908_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_11850_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_11726_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_11371_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_10980_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_10826_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_10768_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_10742_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_10723_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_10314_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_10294_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_10277_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_10270_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_10266_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_10259_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_10255_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_10239_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_10237_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_10234_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_10231_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_10229_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_10226_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_10147_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_10143_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_10132_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_10129_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_10126_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_10122_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_10117_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_10100_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_09813_),
    .X(net759));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(_09574_));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_09549_));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(_09479_));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(_09436_));
 sg13g2_buf_8 fanout764 (.A(_09435_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_09349_),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(_09336_),
    .X(net766));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(_09331_));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_09328_));
 sg13g2_buf_8 fanout769 (.A(_09325_),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_09307_));
 sg13g2_buf_8 fanout771 (.A(_09306_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_09294_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_09270_),
    .X(net773));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_09237_));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(_09234_));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_09230_));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(_09227_));
 sg13g2_buf_8 fanout778 (.A(_09225_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_09182_),
    .X(net779));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_09131_));
 sg13g2_buf_2 fanout781 (.A(_09128_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_09118_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_09090_),
    .X(net783));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(_09084_));
 sg13g2_buf_8 fanout785 (.A(_08466_),
    .X(net785));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(_08464_));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_08459_));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(_08411_));
 sg13g2_buf_4 fanout789 (.X(net789),
    .A(_08394_));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_08391_));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(_08386_));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_08382_));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(_08374_));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(_08369_));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(_08362_));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(_08320_));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_08317_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_08233_));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(_08230_));
 sg13g2_buf_2 fanout800 (.A(_08225_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_07081_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_06378_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_06377_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_06376_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_06374_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_06358_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_06357_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_06355_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_06353_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_06322_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_06321_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_06320_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_06317_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_06314_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_06311_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_06308_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_06305_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_06285_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_06280_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_06273_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_06262_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_06112_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_06111_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_06110_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_06034_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_06033_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_06032_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_05936_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_05935_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_05934_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_05866_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_05865_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_05864_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_05807_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_05773_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_05731_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_04932_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_03433_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_03429_),
    .X(net839));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(_03426_));
 sg13g2_buf_2 fanout841 (.A(_03377_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_02944_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_02943_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_02942_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_02936_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_02935_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_02934_),
    .X(net847));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(_02926_));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(_02924_));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(_02922_));
 sg13g2_buf_2 fanout851 (.A(_02919_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_02917_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_02915_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_02878_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_02848_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_12160_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_12120_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_11981_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_11977_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_11971_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_11930_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_11856_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_11780_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_11725_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_11715_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_11714_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_11707_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_10950_),
    .X(net868));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(_10258_));
 sg13g2_buf_2 fanout870 (.A(_10238_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_10236_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_10233_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_10159_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_10151_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_10149_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_10148_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_10140_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_10131_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_10121_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_10120_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_10116_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_10076_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_09951_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_09897_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_09812_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_09656_),
    .X(net886));
 sg13g2_buf_4 fanout887 (.X(net887),
    .A(_09597_));
 sg13g2_buf_8 fanout888 (.A(_09556_),
    .X(net888));
 sg13g2_buf_8 fanout889 (.A(_09546_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_09428_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_09359_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_09351_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_09293_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_09264_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_09233_),
    .X(net895));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(_09181_));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(_09127_));
 sg13g2_buf_2 fanout898 (.A(_09117_),
    .X(net898));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(_09089_));
 sg13g2_buf_2 fanout900 (.A(_09083_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_08844_),
    .X(net901));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(_08744_));
 sg13g2_buf_2 fanout903 (.A(_08721_),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(_08463_));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_08461_));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(_08410_));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(_08393_));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(_08385_));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(_08381_));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(_08373_));
 sg13g2_buf_2 fanout911 (.A(_08368_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_08319_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_08312_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_08273_),
    .X(net914));
 sg13g2_buf_4 fanout915 (.X(net915),
    .A(_08228_));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(_08227_));
 sg13g2_buf_2 fanout917 (.A(_08224_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_08150_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_08143_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_07246_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_07178_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_07171_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_07156_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_07153_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_06894_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_06763_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_06720_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_06346_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_06345_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_06344_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_06341_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_05945_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_05944_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_05943_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_05877_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_05876_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_05875_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_05816_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_05806_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_05794_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_05777_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_05772_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_05113_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_04926_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_04798_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_04720_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_04570_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_04212_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_03424_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_02925_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_02923_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_02921_),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(_02914_));
 sg13g2_buf_2 fanout954 (.A(_02808_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_02805_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_02801_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_02797_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_02788_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_12581_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_12504_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_12500_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_12496_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_12490_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_12358_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_12297_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_12291_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_12287_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_12279_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_12181_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_12177_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_12173_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_12108_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_12087_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_12081_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_12072_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_12058_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_12013_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_12006_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_12002_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_11998_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_11994_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_11985_),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(_11974_));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_11945_));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(_11938_));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(_11925_));
 sg13g2_buf_2 fanout987 (.A(_11870_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_11868_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_11866_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_11858_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_11807_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_11770_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_11768_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_11766_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_11724_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_11697_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_11696_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_11694_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_11690_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_10227_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_10196_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_10192_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_10190_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_10161_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_10119_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_10115_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_10101_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_10098_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_10075_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_10054_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_10052_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_10000_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_09941_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_09934_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_09928_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_09922_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_09916_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_09910_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_09905_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_09896_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_09749_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_09736_),
    .X(net1022));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(_09457_));
 sg13g2_buf_2 fanout1024 (.A(_09255_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_09251_),
    .X(net1025));
 sg13g2_buf_4 fanout1026 (.X(net1026),
    .A(_09238_));
 sg13g2_buf_2 fanout1027 (.A(_09200_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_09190_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_09137_),
    .X(net1029));
 sg13g2_buf_4 fanout1030 (.X(net1030),
    .A(_09123_));
 sg13g2_buf_2 fanout1031 (.A(_09107_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_09098_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_09097_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_09088_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_09082_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_09080_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_09014_),
    .X(net1037));
 sg13g2_buf_4 fanout1038 (.X(net1038),
    .A(_09012_));
 sg13g2_buf_2 fanout1039 (.A(_08996_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_08892_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_08843_),
    .X(net1041));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(_08782_));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(_08751_));
 sg13g2_buf_4 fanout1044 (.X(net1044),
    .A(_08743_));
 sg13g2_buf_2 fanout1045 (.A(_08680_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_08670_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_08659_),
    .X(net1047));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(_08437_));
 sg13g2_buf_2 fanout1049 (.A(_08436_),
    .X(net1049));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(_08384_));
 sg13g2_buf_2 fanout1051 (.A(_08372_),
    .X(net1051));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(_08367_));
 sg13g2_buf_2 fanout1053 (.A(_08365_),
    .X(net1053));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(_08360_));
 sg13g2_buf_2 fanout1055 (.A(_08358_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_08253_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_08160_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_08147_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_08145_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_08142_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_07952_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_07949_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_07935_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_07889_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_07252_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_07154_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_07152_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_05767_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_11973_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_11959_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_11956_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_11953_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_11949_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_11944_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_11937_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_11924_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_11832_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_11812_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_11795_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_11778_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_11761_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_11758_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_11741_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_11739_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_11736_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_11150_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_11128_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_10764_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_10652_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_10363_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_10197_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_10081_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_10079_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_10078_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_10074_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_10056_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_10055_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_09915_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_09748_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_09744_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_09708_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_09686_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_09215_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_09177_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_09176_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_09079_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_09019_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_08995_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_08891_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_08769_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_08765_),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(_08749_));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(_08742_));
 sg13g2_buf_2 fanout1114 (.A(_08366_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_08364_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_08151_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_08141_),
    .X(net1117));
 sg13g2_tiehi _27249__1118 (.L_HI(net1118));
 sg13g2_tiehi _27250__1119 (.L_HI(net1119));
 sg13g2_tiehi _27251__1120 (.L_HI(net1120));
 sg13g2_tiehi _27252__1121 (.L_HI(net1121));
 sg13g2_tiehi _27253__1122 (.L_HI(net1122));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_rs2_inv$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_cc$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_set_cc$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_DFFE_PP__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_DFFE_PP__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_DFFE_PP__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_DFFE_PP__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_DFFE_PP__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_DFFE_PP__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_DFFE_PP__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_DFFE_PP__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_DFFE_PP__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_DFFE_PP__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_DFFE_PP__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_DFFE_PP__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_DFFE_PP__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_DFFE_PP__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_DFFE_PP__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_DFFE_PP__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_DFFE_PP__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_DFFE_PP__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_DFFE_PP__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_DFFE_PP__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_DFFE_PP__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_DFFE_PP__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_DFFE_PP__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_DFFE_PP__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.spi.r_count[0]$_DFFE_PP__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.spi.r_count[1]$_DFFE_PP__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.spi.r_count[2]$_DFFE_PP__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.spi.r_count[3]$_DFFE_PP__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_count[4]$_DFFE_PP__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_count[5]$_DFFE_PP__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_count[6]$_DFFE_PP__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_count[7]$_DFFE_PP__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_DFFE_PP__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_DFFE_PP__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_DFFE_PP__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_DFFE_PP__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_DFFE_PP__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_DFFE_PP__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_src[0]$_DFFE_PP__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_src[1]$_DFFE_PP__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_src[2]$_DFFE_PP__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3601  (.L_HI(net3601));
 sg13g2_tiehi \r_reset$_DFF_P__3602  (.L_HI(net3602));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_310_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00237_));
 sg13g2_antennanp ANTENNA_2 (.A(_00789_));
 sg13g2_antennanp ANTENNA_3 (.A(_00798_));
 sg13g2_antennanp ANTENNA_4 (.A(_00930_));
 sg13g2_antennanp ANTENNA_5 (.A(_02788_));
 sg13g2_antennanp ANTENNA_6 (.A(_02788_));
 sg13g2_antennanp ANTENNA_7 (.A(_02788_));
 sg13g2_antennanp ANTENNA_8 (.A(_02788_));
 sg13g2_antennanp ANTENNA_9 (.A(_02788_));
 sg13g2_antennanp ANTENNA_10 (.A(_02788_));
 sg13g2_antennanp ANTENNA_11 (.A(_02788_));
 sg13g2_antennanp ANTENNA_12 (.A(_02788_));
 sg13g2_antennanp ANTENNA_13 (.A(_02788_));
 sg13g2_antennanp ANTENNA_14 (.A(_02797_));
 sg13g2_antennanp ANTENNA_15 (.A(_02797_));
 sg13g2_antennanp ANTENNA_16 (.A(_02797_));
 sg13g2_antennanp ANTENNA_17 (.A(_02797_));
 sg13g2_antennanp ANTENNA_18 (.A(_02797_));
 sg13g2_antennanp ANTENNA_19 (.A(_02797_));
 sg13g2_antennanp ANTENNA_20 (.A(_02797_));
 sg13g2_antennanp ANTENNA_21 (.A(_02797_));
 sg13g2_antennanp ANTENNA_22 (.A(_02797_));
 sg13g2_antennanp ANTENNA_23 (.A(_02801_));
 sg13g2_antennanp ANTENNA_24 (.A(_02801_));
 sg13g2_antennanp ANTENNA_25 (.A(_02801_));
 sg13g2_antennanp ANTENNA_26 (.A(_02801_));
 sg13g2_antennanp ANTENNA_27 (.A(_02801_));
 sg13g2_antennanp ANTENNA_28 (.A(_02801_));
 sg13g2_antennanp ANTENNA_29 (.A(_02801_));
 sg13g2_antennanp ANTENNA_30 (.A(_02801_));
 sg13g2_antennanp ANTENNA_31 (.A(_02801_));
 sg13g2_antennanp ANTENNA_32 (.A(_02805_));
 sg13g2_antennanp ANTENNA_33 (.A(_02805_));
 sg13g2_antennanp ANTENNA_34 (.A(_02805_));
 sg13g2_antennanp ANTENNA_35 (.A(_02805_));
 sg13g2_antennanp ANTENNA_36 (.A(_02805_));
 sg13g2_antennanp ANTENNA_37 (.A(_02805_));
 sg13g2_antennanp ANTENNA_38 (.A(_02805_));
 sg13g2_antennanp ANTENNA_39 (.A(_02805_));
 sg13g2_antennanp ANTENNA_40 (.A(_02805_));
 sg13g2_antennanp ANTENNA_41 (.A(_02908_));
 sg13g2_antennanp ANTENNA_42 (.A(_02908_));
 sg13g2_antennanp ANTENNA_43 (.A(_02908_));
 sg13g2_antennanp ANTENNA_44 (.A(_02908_));
 sg13g2_antennanp ANTENNA_45 (.A(_02908_));
 sg13g2_antennanp ANTENNA_46 (.A(_02908_));
 sg13g2_antennanp ANTENNA_47 (.A(_02914_));
 sg13g2_antennanp ANTENNA_48 (.A(_02914_));
 sg13g2_antennanp ANTENNA_49 (.A(_02914_));
 sg13g2_antennanp ANTENNA_50 (.A(_02914_));
 sg13g2_antennanp ANTENNA_51 (.A(_02914_));
 sg13g2_antennanp ANTENNA_52 (.A(_02914_));
 sg13g2_antennanp ANTENNA_53 (.A(_02914_));
 sg13g2_antennanp ANTENNA_54 (.A(_02914_));
 sg13g2_antennanp ANTENNA_55 (.A(_02917_));
 sg13g2_antennanp ANTENNA_56 (.A(_02917_));
 sg13g2_antennanp ANTENNA_57 (.A(_02917_));
 sg13g2_antennanp ANTENNA_58 (.A(_02917_));
 sg13g2_antennanp ANTENNA_59 (.A(_02918_));
 sg13g2_antennanp ANTENNA_60 (.A(_02918_));
 sg13g2_antennanp ANTENNA_61 (.A(_02918_));
 sg13g2_antennanp ANTENNA_62 (.A(_02919_));
 sg13g2_antennanp ANTENNA_63 (.A(_02919_));
 sg13g2_antennanp ANTENNA_64 (.A(_02919_));
 sg13g2_antennanp ANTENNA_65 (.A(_02919_));
 sg13g2_antennanp ANTENNA_66 (.A(_02920_));
 sg13g2_antennanp ANTENNA_67 (.A(_02920_));
 sg13g2_antennanp ANTENNA_68 (.A(_02920_));
 sg13g2_antennanp ANTENNA_69 (.A(_02920_));
 sg13g2_antennanp ANTENNA_70 (.A(_02920_));
 sg13g2_antennanp ANTENNA_71 (.A(_02920_));
 sg13g2_antennanp ANTENNA_72 (.A(_02920_));
 sg13g2_antennanp ANTENNA_73 (.A(_02920_));
 sg13g2_antennanp ANTENNA_74 (.A(_02920_));
 sg13g2_antennanp ANTENNA_75 (.A(_02920_));
 sg13g2_antennanp ANTENNA_76 (.A(_02922_));
 sg13g2_antennanp ANTENNA_77 (.A(_02922_));
 sg13g2_antennanp ANTENNA_78 (.A(_02922_));
 sg13g2_antennanp ANTENNA_79 (.A(_02927_));
 sg13g2_antennanp ANTENNA_80 (.A(_02927_));
 sg13g2_antennanp ANTENNA_81 (.A(_02927_));
 sg13g2_antennanp ANTENNA_82 (.A(_02927_));
 sg13g2_antennanp ANTENNA_83 (.A(_02927_));
 sg13g2_antennanp ANTENNA_84 (.A(_02927_));
 sg13g2_antennanp ANTENNA_85 (.A(_02927_));
 sg13g2_antennanp ANTENNA_86 (.A(_02927_));
 sg13g2_antennanp ANTENNA_87 (.A(_02927_));
 sg13g2_antennanp ANTENNA_88 (.A(_02927_));
 sg13g2_antennanp ANTENNA_89 (.A(_02936_));
 sg13g2_antennanp ANTENNA_90 (.A(_02936_));
 sg13g2_antennanp ANTENNA_91 (.A(_02936_));
 sg13g2_antennanp ANTENNA_92 (.A(_03293_));
 sg13g2_antennanp ANTENNA_93 (.A(_03293_));
 sg13g2_antennanp ANTENNA_94 (.A(_03317_));
 sg13g2_antennanp ANTENNA_95 (.A(_03317_));
 sg13g2_antennanp ANTENNA_96 (.A(_03323_));
 sg13g2_antennanp ANTENNA_97 (.A(_03323_));
 sg13g2_antennanp ANTENNA_98 (.A(_03324_));
 sg13g2_antennanp ANTENNA_99 (.A(_03329_));
 sg13g2_antennanp ANTENNA_100 (.A(_03397_));
 sg13g2_antennanp ANTENNA_101 (.A(_03397_));
 sg13g2_antennanp ANTENNA_102 (.A(_03397_));
 sg13g2_antennanp ANTENNA_103 (.A(_03397_));
 sg13g2_antennanp ANTENNA_104 (.A(_03519_));
 sg13g2_antennanp ANTENNA_105 (.A(_03693_));
 sg13g2_antennanp ANTENNA_106 (.A(_03693_));
 sg13g2_antennanp ANTENNA_107 (.A(_03693_));
 sg13g2_antennanp ANTENNA_108 (.A(_03693_));
 sg13g2_antennanp ANTENNA_109 (.A(_03696_));
 sg13g2_antennanp ANTENNA_110 (.A(_03696_));
 sg13g2_antennanp ANTENNA_111 (.A(_03696_));
 sg13g2_antennanp ANTENNA_112 (.A(_03696_));
 sg13g2_antennanp ANTENNA_113 (.A(_03697_));
 sg13g2_antennanp ANTENNA_114 (.A(_03697_));
 sg13g2_antennanp ANTENNA_115 (.A(_03697_));
 sg13g2_antennanp ANTENNA_116 (.A(_04980_));
 sg13g2_antennanp ANTENNA_117 (.A(_05114_));
 sg13g2_antennanp ANTENNA_118 (.A(_05142_));
 sg13g2_antennanp ANTENNA_119 (.A(_05173_));
 sg13g2_antennanp ANTENNA_120 (.A(_05173_));
 sg13g2_antennanp ANTENNA_121 (.A(_05204_));
 sg13g2_antennanp ANTENNA_122 (.A(_05236_));
 sg13g2_antennanp ANTENNA_123 (.A(_05248_));
 sg13g2_antennanp ANTENNA_124 (.A(_05255_));
 sg13g2_antennanp ANTENNA_125 (.A(_05335_));
 sg13g2_antennanp ANTENNA_126 (.A(_05407_));
 sg13g2_antennanp ANTENNA_127 (.A(_05412_));
 sg13g2_antennanp ANTENNA_128 (.A(_05477_));
 sg13g2_antennanp ANTENNA_129 (.A(_05556_));
 sg13g2_antennanp ANTENNA_130 (.A(_05681_));
 sg13g2_antennanp ANTENNA_131 (.A(_05695_));
 sg13g2_antennanp ANTENNA_132 (.A(_05708_));
 sg13g2_antennanp ANTENNA_133 (.A(_05735_));
 sg13g2_antennanp ANTENNA_134 (.A(_05756_));
 sg13g2_antennanp ANTENNA_135 (.A(_06178_));
 sg13g2_antennanp ANTENNA_136 (.A(_06178_));
 sg13g2_antennanp ANTENNA_137 (.A(_06178_));
 sg13g2_antennanp ANTENNA_138 (.A(_06178_));
 sg13g2_antennanp ANTENNA_139 (.A(_06655_));
 sg13g2_antennanp ANTENNA_140 (.A(_06655_));
 sg13g2_antennanp ANTENNA_141 (.A(_06655_));
 sg13g2_antennanp ANTENNA_142 (.A(_06655_));
 sg13g2_antennanp ANTENNA_143 (.A(_07439_));
 sg13g2_antennanp ANTENNA_144 (.A(_07439_));
 sg13g2_antennanp ANTENNA_145 (.A(_07476_));
 sg13g2_antennanp ANTENNA_146 (.A(_07476_));
 sg13g2_antennanp ANTENNA_147 (.A(_07476_));
 sg13g2_antennanp ANTENNA_148 (.A(_07737_));
 sg13g2_antennanp ANTENNA_149 (.A(_07737_));
 sg13g2_antennanp ANTENNA_150 (.A(_07737_));
 sg13g2_antennanp ANTENNA_151 (.A(_07737_));
 sg13g2_antennanp ANTENNA_152 (.A(_07737_));
 sg13g2_antennanp ANTENNA_153 (.A(_07737_));
 sg13g2_antennanp ANTENNA_154 (.A(_07737_));
 sg13g2_antennanp ANTENNA_155 (.A(_07737_));
 sg13g2_antennanp ANTENNA_156 (.A(_07737_));
 sg13g2_antennanp ANTENNA_157 (.A(_07737_));
 sg13g2_antennanp ANTENNA_158 (.A(_08224_));
 sg13g2_antennanp ANTENNA_159 (.A(_08224_));
 sg13g2_antennanp ANTENNA_160 (.A(_08224_));
 sg13g2_antennanp ANTENNA_161 (.A(_08253_));
 sg13g2_antennanp ANTENNA_162 (.A(_08253_));
 sg13g2_antennanp ANTENNA_163 (.A(_08253_));
 sg13g2_antennanp ANTENNA_164 (.A(_08401_));
 sg13g2_antennanp ANTENNA_165 (.A(_08401_));
 sg13g2_antennanp ANTENNA_166 (.A(_08401_));
 sg13g2_antennanp ANTENNA_167 (.A(_08401_));
 sg13g2_antennanp ANTENNA_168 (.A(_08401_));
 sg13g2_antennanp ANTENNA_169 (.A(_08401_));
 sg13g2_antennanp ANTENNA_170 (.A(_08426_));
 sg13g2_antennanp ANTENNA_171 (.A(_08426_));
 sg13g2_antennanp ANTENNA_172 (.A(_08426_));
 sg13g2_antennanp ANTENNA_173 (.A(_08450_));
 sg13g2_antennanp ANTENNA_174 (.A(_08450_));
 sg13g2_antennanp ANTENNA_175 (.A(_08450_));
 sg13g2_antennanp ANTENNA_176 (.A(_08450_));
 sg13g2_antennanp ANTENNA_177 (.A(_08450_));
 sg13g2_antennanp ANTENNA_178 (.A(_08450_));
 sg13g2_antennanp ANTENNA_179 (.A(_08450_));
 sg13g2_antennanp ANTENNA_180 (.A(_08450_));
 sg13g2_antennanp ANTENNA_181 (.A(_08450_));
 sg13g2_antennanp ANTENNA_182 (.A(_08476_));
 sg13g2_antennanp ANTENNA_183 (.A(_08476_));
 sg13g2_antennanp ANTENNA_184 (.A(_08498_));
 sg13g2_antennanp ANTENNA_185 (.A(_08498_));
 sg13g2_antennanp ANTENNA_186 (.A(_08498_));
 sg13g2_antennanp ANTENNA_187 (.A(_08522_));
 sg13g2_antennanp ANTENNA_188 (.A(_08522_));
 sg13g2_antennanp ANTENNA_189 (.A(_08522_));
 sg13g2_antennanp ANTENNA_190 (.A(_08522_));
 sg13g2_antennanp ANTENNA_191 (.A(_08522_));
 sg13g2_antennanp ANTENNA_192 (.A(_08522_));
 sg13g2_antennanp ANTENNA_193 (.A(_08522_));
 sg13g2_antennanp ANTENNA_194 (.A(_08522_));
 sg13g2_antennanp ANTENNA_195 (.A(_08522_));
 sg13g2_antennanp ANTENNA_196 (.A(_08543_));
 sg13g2_antennanp ANTENNA_197 (.A(_08543_));
 sg13g2_antennanp ANTENNA_198 (.A(_08543_));
 sg13g2_antennanp ANTENNA_199 (.A(_08543_));
 sg13g2_antennanp ANTENNA_200 (.A(_08543_));
 sg13g2_antennanp ANTENNA_201 (.A(_08543_));
 sg13g2_antennanp ANTENNA_202 (.A(_08543_));
 sg13g2_antennanp ANTENNA_203 (.A(_08543_));
 sg13g2_antennanp ANTENNA_204 (.A(_08543_));
 sg13g2_antennanp ANTENNA_205 (.A(_08564_));
 sg13g2_antennanp ANTENNA_206 (.A(_08564_));
 sg13g2_antennanp ANTENNA_207 (.A(_08564_));
 sg13g2_antennanp ANTENNA_208 (.A(_08564_));
 sg13g2_antennanp ANTENNA_209 (.A(_08564_));
 sg13g2_antennanp ANTENNA_210 (.A(_08564_));
 sg13g2_antennanp ANTENNA_211 (.A(_08564_));
 sg13g2_antennanp ANTENNA_212 (.A(_08564_));
 sg13g2_antennanp ANTENNA_213 (.A(_08564_));
 sg13g2_antennanp ANTENNA_214 (.A(_08583_));
 sg13g2_antennanp ANTENNA_215 (.A(_08584_));
 sg13g2_antennanp ANTENNA_216 (.A(_08584_));
 sg13g2_antennanp ANTENNA_217 (.A(_08607_));
 sg13g2_antennanp ANTENNA_218 (.A(_08607_));
 sg13g2_antennanp ANTENNA_219 (.A(_08607_));
 sg13g2_antennanp ANTENNA_220 (.A(_08607_));
 sg13g2_antennanp ANTENNA_221 (.A(_08607_));
 sg13g2_antennanp ANTENNA_222 (.A(_08607_));
 sg13g2_antennanp ANTENNA_223 (.A(_08627_));
 sg13g2_antennanp ANTENNA_224 (.A(_08650_));
 sg13g2_antennanp ANTENNA_225 (.A(_08650_));
 sg13g2_antennanp ANTENNA_226 (.A(_08650_));
 sg13g2_antennanp ANTENNA_227 (.A(_08650_));
 sg13g2_antennanp ANTENNA_228 (.A(_08650_));
 sg13g2_antennanp ANTENNA_229 (.A(_08650_));
 sg13g2_antennanp ANTENNA_230 (.A(_08680_));
 sg13g2_antennanp ANTENNA_231 (.A(_08680_));
 sg13g2_antennanp ANTENNA_232 (.A(_08680_));
 sg13g2_antennanp ANTENNA_233 (.A(_08680_));
 sg13g2_antennanp ANTENNA_234 (.A(_08732_));
 sg13g2_antennanp ANTENNA_235 (.A(_08732_));
 sg13g2_antennanp ANTENNA_236 (.A(_08732_));
 sg13g2_antennanp ANTENNA_237 (.A(_08732_));
 sg13g2_antennanp ANTENNA_238 (.A(_08732_));
 sg13g2_antennanp ANTENNA_239 (.A(_08732_));
 sg13g2_antennanp ANTENNA_240 (.A(_09012_));
 sg13g2_antennanp ANTENNA_241 (.A(_09012_));
 sg13g2_antennanp ANTENNA_242 (.A(_09012_));
 sg13g2_antennanp ANTENNA_243 (.A(_09012_));
 sg13g2_antennanp ANTENNA_244 (.A(_09012_));
 sg13g2_antennanp ANTENNA_245 (.A(_09012_));
 sg13g2_antennanp ANTENNA_246 (.A(_09012_));
 sg13g2_antennanp ANTENNA_247 (.A(_09012_));
 sg13g2_antennanp ANTENNA_248 (.A(_09014_));
 sg13g2_antennanp ANTENNA_249 (.A(_09014_));
 sg13g2_antennanp ANTENNA_250 (.A(_09014_));
 sg13g2_antennanp ANTENNA_251 (.A(_09014_));
 sg13g2_antennanp ANTENNA_252 (.A(_09014_));
 sg13g2_antennanp ANTENNA_253 (.A(_09014_));
 sg13g2_antennanp ANTENNA_254 (.A(_09014_));
 sg13g2_antennanp ANTENNA_255 (.A(_09014_));
 sg13g2_antennanp ANTENNA_256 (.A(_09014_));
 sg13g2_antennanp ANTENNA_257 (.A(_09040_));
 sg13g2_antennanp ANTENNA_258 (.A(_09040_));
 sg13g2_antennanp ANTENNA_259 (.A(_09040_));
 sg13g2_antennanp ANTENNA_260 (.A(_09040_));
 sg13g2_antennanp ANTENNA_261 (.A(_09090_));
 sg13g2_antennanp ANTENNA_262 (.A(_09090_));
 sg13g2_antennanp ANTENNA_263 (.A(_09090_));
 sg13g2_antennanp ANTENNA_264 (.A(_09090_));
 sg13g2_antennanp ANTENNA_265 (.A(_09094_));
 sg13g2_antennanp ANTENNA_266 (.A(_09094_));
 sg13g2_antennanp ANTENNA_267 (.A(_09094_));
 sg13g2_antennanp ANTENNA_268 (.A(_09094_));
 sg13g2_antennanp ANTENNA_269 (.A(_09095_));
 sg13g2_antennanp ANTENNA_270 (.A(_09095_));
 sg13g2_antennanp ANTENNA_271 (.A(_09102_));
 sg13g2_antennanp ANTENNA_272 (.A(_09119_));
 sg13g2_antennanp ANTENNA_273 (.A(_09119_));
 sg13g2_antennanp ANTENNA_274 (.A(_09119_));
 sg13g2_antennanp ANTENNA_275 (.A(_09119_));
 sg13g2_antennanp ANTENNA_276 (.A(_09119_));
 sg13g2_antennanp ANTENNA_277 (.A(_09119_));
 sg13g2_antennanp ANTENNA_278 (.A(_09123_));
 sg13g2_antennanp ANTENNA_279 (.A(_09123_));
 sg13g2_antennanp ANTENNA_280 (.A(_09123_));
 sg13g2_antennanp ANTENNA_281 (.A(_09125_));
 sg13g2_antennanp ANTENNA_282 (.A(_09125_));
 sg13g2_antennanp ANTENNA_283 (.A(_09130_));
 sg13g2_antennanp ANTENNA_284 (.A(_09130_));
 sg13g2_antennanp ANTENNA_285 (.A(_09130_));
 sg13g2_antennanp ANTENNA_286 (.A(_09130_));
 sg13g2_antennanp ANTENNA_287 (.A(_09130_));
 sg13g2_antennanp ANTENNA_288 (.A(_09130_));
 sg13g2_antennanp ANTENNA_289 (.A(_09130_));
 sg13g2_antennanp ANTENNA_290 (.A(_09130_));
 sg13g2_antennanp ANTENNA_291 (.A(_09130_));
 sg13g2_antennanp ANTENNA_292 (.A(_09130_));
 sg13g2_antennanp ANTENNA_293 (.A(_09130_));
 sg13g2_antennanp ANTENNA_294 (.A(_09130_));
 sg13g2_antennanp ANTENNA_295 (.A(_09130_));
 sg13g2_antennanp ANTENNA_296 (.A(_09181_));
 sg13g2_antennanp ANTENNA_297 (.A(_09181_));
 sg13g2_antennanp ANTENNA_298 (.A(_09181_));
 sg13g2_antennanp ANTENNA_299 (.A(_09181_));
 sg13g2_antennanp ANTENNA_300 (.A(_09181_));
 sg13g2_antennanp ANTENNA_301 (.A(_09181_));
 sg13g2_antennanp ANTENNA_302 (.A(_09181_));
 sg13g2_antennanp ANTENNA_303 (.A(_09181_));
 sg13g2_antennanp ANTENNA_304 (.A(_09181_));
 sg13g2_antennanp ANTENNA_305 (.A(_09181_));
 sg13g2_antennanp ANTENNA_306 (.A(_09246_));
 sg13g2_antennanp ANTENNA_307 (.A(_09312_));
 sg13g2_antennanp ANTENNA_308 (.A(_09315_));
 sg13g2_antennanp ANTENNA_309 (.A(_09315_));
 sg13g2_antennanp ANTENNA_310 (.A(_09341_));
 sg13g2_antennanp ANTENNA_311 (.A(_09443_));
 sg13g2_antennanp ANTENNA_312 (.A(_09466_));
 sg13g2_antennanp ANTENNA_313 (.A(_09492_));
 sg13g2_antennanp ANTENNA_314 (.A(_09492_));
 sg13g2_antennanp ANTENNA_315 (.A(_09492_));
 sg13g2_antennanp ANTENNA_316 (.A(_09514_));
 sg13g2_antennanp ANTENNA_317 (.A(_09536_));
 sg13g2_antennanp ANTENNA_318 (.A(_09561_));
 sg13g2_antennanp ANTENNA_319 (.A(_09585_));
 sg13g2_antennanp ANTENNA_320 (.A(_09608_));
 sg13g2_antennanp ANTENNA_321 (.A(_09630_));
 sg13g2_antennanp ANTENNA_322 (.A(_09759_));
 sg13g2_antennanp ANTENNA_323 (.A(_09943_));
 sg13g2_antennanp ANTENNA_324 (.A(_09943_));
 sg13g2_antennanp ANTENNA_325 (.A(_09943_));
 sg13g2_antennanp ANTENNA_326 (.A(_09944_));
 sg13g2_antennanp ANTENNA_327 (.A(_09944_));
 sg13g2_antennanp ANTENNA_328 (.A(_09944_));
 sg13g2_antennanp ANTENNA_329 (.A(_09944_));
 sg13g2_antennanp ANTENNA_330 (.A(_09952_));
 sg13g2_antennanp ANTENNA_331 (.A(_09952_));
 sg13g2_antennanp ANTENNA_332 (.A(_09952_));
 sg13g2_antennanp ANTENNA_333 (.A(_09952_));
 sg13g2_antennanp ANTENNA_334 (.A(_09952_));
 sg13g2_antennanp ANTENNA_335 (.A(_09952_));
 sg13g2_antennanp ANTENNA_336 (.A(_09952_));
 sg13g2_antennanp ANTENNA_337 (.A(_09952_));
 sg13g2_antennanp ANTENNA_338 (.A(_09952_));
 sg13g2_antennanp ANTENNA_339 (.A(_09952_));
 sg13g2_antennanp ANTENNA_340 (.A(_10018_));
 sg13g2_antennanp ANTENNA_341 (.A(_10018_));
 sg13g2_antennanp ANTENNA_342 (.A(_10018_));
 sg13g2_antennanp ANTENNA_343 (.A(_10018_));
 sg13g2_antennanp ANTENNA_344 (.A(_10018_));
 sg13g2_antennanp ANTENNA_345 (.A(_10018_));
 sg13g2_antennanp ANTENNA_346 (.A(_10018_));
 sg13g2_antennanp ANTENNA_347 (.A(_10018_));
 sg13g2_antennanp ANTENNA_348 (.A(_10187_));
 sg13g2_antennanp ANTENNA_349 (.A(_10187_));
 sg13g2_antennanp ANTENNA_350 (.A(_10187_));
 sg13g2_antennanp ANTENNA_351 (.A(_10187_));
 sg13g2_antennanp ANTENNA_352 (.A(_10429_));
 sg13g2_antennanp ANTENNA_353 (.A(_10758_));
 sg13g2_antennanp ANTENNA_354 (.A(_10758_));
 sg13g2_antennanp ANTENNA_355 (.A(_10758_));
 sg13g2_antennanp ANTENNA_356 (.A(_10758_));
 sg13g2_antennanp ANTENNA_357 (.A(_10758_));
 sg13g2_antennanp ANTENNA_358 (.A(_10758_));
 sg13g2_antennanp ANTENNA_359 (.A(_11070_));
 sg13g2_antennanp ANTENNA_360 (.A(_11070_));
 sg13g2_antennanp ANTENNA_361 (.A(_11070_));
 sg13g2_antennanp ANTENNA_362 (.A(_11070_));
 sg13g2_antennanp ANTENNA_363 (.A(_11070_));
 sg13g2_antennanp ANTENNA_364 (.A(_11070_));
 sg13g2_antennanp ANTENNA_365 (.A(_11761_));
 sg13g2_antennanp ANTENNA_366 (.A(_11761_));
 sg13g2_antennanp ANTENNA_367 (.A(_11761_));
 sg13g2_antennanp ANTENNA_368 (.A(_11761_));
 sg13g2_antennanp ANTENNA_369 (.A(_11761_));
 sg13g2_antennanp ANTENNA_370 (.A(_11761_));
 sg13g2_antennanp ANTENNA_371 (.A(_11761_));
 sg13g2_antennanp ANTENNA_372 (.A(_11761_));
 sg13g2_antennanp ANTENNA_373 (.A(_11761_));
 sg13g2_antennanp ANTENNA_374 (.A(_11795_));
 sg13g2_antennanp ANTENNA_375 (.A(_11795_));
 sg13g2_antennanp ANTENNA_376 (.A(_11795_));
 sg13g2_antennanp ANTENNA_377 (.A(_11795_));
 sg13g2_antennanp ANTENNA_378 (.A(_11795_));
 sg13g2_antennanp ANTENNA_379 (.A(_11795_));
 sg13g2_antennanp ANTENNA_380 (.A(_11795_));
 sg13g2_antennanp ANTENNA_381 (.A(_11795_));
 sg13g2_antennanp ANTENNA_382 (.A(_11795_));
 sg13g2_antennanp ANTENNA_383 (.A(_11812_));
 sg13g2_antennanp ANTENNA_384 (.A(_11812_));
 sg13g2_antennanp ANTENNA_385 (.A(_11812_));
 sg13g2_antennanp ANTENNA_386 (.A(_11812_));
 sg13g2_antennanp ANTENNA_387 (.A(_11812_));
 sg13g2_antennanp ANTENNA_388 (.A(_11812_));
 sg13g2_antennanp ANTENNA_389 (.A(_11812_));
 sg13g2_antennanp ANTENNA_390 (.A(_11812_));
 sg13g2_antennanp ANTENNA_391 (.A(_11812_));
 sg13g2_antennanp ANTENNA_392 (.A(_11832_));
 sg13g2_antennanp ANTENNA_393 (.A(_11832_));
 sg13g2_antennanp ANTENNA_394 (.A(_11832_));
 sg13g2_antennanp ANTENNA_395 (.A(_11832_));
 sg13g2_antennanp ANTENNA_396 (.A(_11832_));
 sg13g2_antennanp ANTENNA_397 (.A(_11832_));
 sg13g2_antennanp ANTENNA_398 (.A(_11832_));
 sg13g2_antennanp ANTENNA_399 (.A(_11832_));
 sg13g2_antennanp ANTENNA_400 (.A(_11832_));
 sg13g2_antennanp ANTENNA_401 (.A(_11925_));
 sg13g2_antennanp ANTENNA_402 (.A(_11925_));
 sg13g2_antennanp ANTENNA_403 (.A(_11925_));
 sg13g2_antennanp ANTENNA_404 (.A(_11925_));
 sg13g2_antennanp ANTENNA_405 (.A(_11925_));
 sg13g2_antennanp ANTENNA_406 (.A(_11925_));
 sg13g2_antennanp ANTENNA_407 (.A(_11925_));
 sg13g2_antennanp ANTENNA_408 (.A(_11925_));
 sg13g2_antennanp ANTENNA_409 (.A(_11925_));
 sg13g2_antennanp ANTENNA_410 (.A(_11938_));
 sg13g2_antennanp ANTENNA_411 (.A(_11938_));
 sg13g2_antennanp ANTENNA_412 (.A(_11938_));
 sg13g2_antennanp ANTENNA_413 (.A(_11938_));
 sg13g2_antennanp ANTENNA_414 (.A(_11938_));
 sg13g2_antennanp ANTENNA_415 (.A(_11938_));
 sg13g2_antennanp ANTENNA_416 (.A(_11938_));
 sg13g2_antennanp ANTENNA_417 (.A(_11938_));
 sg13g2_antennanp ANTENNA_418 (.A(_11938_));
 sg13g2_antennanp ANTENNA_419 (.A(_11945_));
 sg13g2_antennanp ANTENNA_420 (.A(_11945_));
 sg13g2_antennanp ANTENNA_421 (.A(_11945_));
 sg13g2_antennanp ANTENNA_422 (.A(_11945_));
 sg13g2_antennanp ANTENNA_423 (.A(_11945_));
 sg13g2_antennanp ANTENNA_424 (.A(_11945_));
 sg13g2_antennanp ANTENNA_425 (.A(_11945_));
 sg13g2_antennanp ANTENNA_426 (.A(_11945_));
 sg13g2_antennanp ANTENNA_427 (.A(_11945_));
 sg13g2_antennanp ANTENNA_428 (.A(_11974_));
 sg13g2_antennanp ANTENNA_429 (.A(_11974_));
 sg13g2_antennanp ANTENNA_430 (.A(_11974_));
 sg13g2_antennanp ANTENNA_431 (.A(_11974_));
 sg13g2_antennanp ANTENNA_432 (.A(_11974_));
 sg13g2_antennanp ANTENNA_433 (.A(_11974_));
 sg13g2_antennanp ANTENNA_434 (.A(_11974_));
 sg13g2_antennanp ANTENNA_435 (.A(_11974_));
 sg13g2_antennanp ANTENNA_436 (.A(clk));
 sg13g2_antennanp ANTENNA_437 (.A(clk));
 sg13g2_antennanp ANTENNA_438 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_439 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_440 (.A(net3));
 sg13g2_antennanp ANTENNA_441 (.A(net3));
 sg13g2_antennanp ANTENNA_442 (.A(net3));
 sg13g2_antennanp ANTENNA_443 (.A(net151));
 sg13g2_antennanp ANTENNA_444 (.A(net151));
 sg13g2_antennanp ANTENNA_445 (.A(net151));
 sg13g2_antennanp ANTENNA_446 (.A(net151));
 sg13g2_antennanp ANTENNA_447 (.A(net151));
 sg13g2_antennanp ANTENNA_448 (.A(net151));
 sg13g2_antennanp ANTENNA_449 (.A(net151));
 sg13g2_antennanp ANTENNA_450 (.A(net151));
 sg13g2_antennanp ANTENNA_451 (.A(net151));
 sg13g2_antennanp ANTENNA_452 (.A(net366));
 sg13g2_antennanp ANTENNA_453 (.A(net366));
 sg13g2_antennanp ANTENNA_454 (.A(net366));
 sg13g2_antennanp ANTENNA_455 (.A(net366));
 sg13g2_antennanp ANTENNA_456 (.A(net366));
 sg13g2_antennanp ANTENNA_457 (.A(net366));
 sg13g2_antennanp ANTENNA_458 (.A(net366));
 sg13g2_antennanp ANTENNA_459 (.A(net366));
 sg13g2_antennanp ANTENNA_460 (.A(net366));
 sg13g2_antennanp ANTENNA_461 (.A(net366));
 sg13g2_antennanp ANTENNA_462 (.A(net366));
 sg13g2_antennanp ANTENNA_463 (.A(net366));
 sg13g2_antennanp ANTENNA_464 (.A(net468));
 sg13g2_antennanp ANTENNA_465 (.A(net468));
 sg13g2_antennanp ANTENNA_466 (.A(net468));
 sg13g2_antennanp ANTENNA_467 (.A(net468));
 sg13g2_antennanp ANTENNA_468 (.A(net468));
 sg13g2_antennanp ANTENNA_469 (.A(net468));
 sg13g2_antennanp ANTENNA_470 (.A(net468));
 sg13g2_antennanp ANTENNA_471 (.A(net468));
 sg13g2_antennanp ANTENNA_472 (.A(net468));
 sg13g2_antennanp ANTENNA_473 (.A(net496));
 sg13g2_antennanp ANTENNA_474 (.A(net496));
 sg13g2_antennanp ANTENNA_475 (.A(net496));
 sg13g2_antennanp ANTENNA_476 (.A(net496));
 sg13g2_antennanp ANTENNA_477 (.A(net496));
 sg13g2_antennanp ANTENNA_478 (.A(net496));
 sg13g2_antennanp ANTENNA_479 (.A(net496));
 sg13g2_antennanp ANTENNA_480 (.A(net496));
 sg13g2_antennanp ANTENNA_481 (.A(net496));
 sg13g2_antennanp ANTENNA_482 (.A(net496));
 sg13g2_antennanp ANTENNA_483 (.A(net496));
 sg13g2_antennanp ANTENNA_484 (.A(net551));
 sg13g2_antennanp ANTENNA_485 (.A(net551));
 sg13g2_antennanp ANTENNA_486 (.A(net551));
 sg13g2_antennanp ANTENNA_487 (.A(net551));
 sg13g2_antennanp ANTENNA_488 (.A(net551));
 sg13g2_antennanp ANTENNA_489 (.A(net551));
 sg13g2_antennanp ANTENNA_490 (.A(net551));
 sg13g2_antennanp ANTENNA_491 (.A(net551));
 sg13g2_antennanp ANTENNA_492 (.A(net551));
 sg13g2_antennanp ANTENNA_493 (.A(net551));
 sg13g2_antennanp ANTENNA_494 (.A(net551));
 sg13g2_antennanp ANTENNA_495 (.A(net551));
 sg13g2_antennanp ANTENNA_496 (.A(net551));
 sg13g2_antennanp ANTENNA_497 (.A(net551));
 sg13g2_antennanp ANTENNA_498 (.A(net551));
 sg13g2_antennanp ANTENNA_499 (.A(net551));
 sg13g2_antennanp ANTENNA_500 (.A(net551));
 sg13g2_antennanp ANTENNA_501 (.A(net551));
 sg13g2_antennanp ANTENNA_502 (.A(net551));
 sg13g2_antennanp ANTENNA_503 (.A(net571));
 sg13g2_antennanp ANTENNA_504 (.A(net571));
 sg13g2_antennanp ANTENNA_505 (.A(net571));
 sg13g2_antennanp ANTENNA_506 (.A(net571));
 sg13g2_antennanp ANTENNA_507 (.A(net571));
 sg13g2_antennanp ANTENNA_508 (.A(net571));
 sg13g2_antennanp ANTENNA_509 (.A(net571));
 sg13g2_antennanp ANTENNA_510 (.A(net571));
 sg13g2_antennanp ANTENNA_511 (.A(net571));
 sg13g2_antennanp ANTENNA_512 (.A(net571));
 sg13g2_antennanp ANTENNA_513 (.A(net571));
 sg13g2_antennanp ANTENNA_514 (.A(net594));
 sg13g2_antennanp ANTENNA_515 (.A(net594));
 sg13g2_antennanp ANTENNA_516 (.A(net594));
 sg13g2_antennanp ANTENNA_517 (.A(net594));
 sg13g2_antennanp ANTENNA_518 (.A(net594));
 sg13g2_antennanp ANTENNA_519 (.A(net594));
 sg13g2_antennanp ANTENNA_520 (.A(net594));
 sg13g2_antennanp ANTENNA_521 (.A(net594));
 sg13g2_antennanp ANTENNA_522 (.A(net594));
 sg13g2_antennanp ANTENNA_523 (.A(net594));
 sg13g2_antennanp ANTENNA_524 (.A(net594));
 sg13g2_antennanp ANTENNA_525 (.A(net594));
 sg13g2_antennanp ANTENNA_526 (.A(net594));
 sg13g2_antennanp ANTENNA_527 (.A(net638));
 sg13g2_antennanp ANTENNA_528 (.A(net638));
 sg13g2_antennanp ANTENNA_529 (.A(net638));
 sg13g2_antennanp ANTENNA_530 (.A(net638));
 sg13g2_antennanp ANTENNA_531 (.A(net638));
 sg13g2_antennanp ANTENNA_532 (.A(net638));
 sg13g2_antennanp ANTENNA_533 (.A(net638));
 sg13g2_antennanp ANTENNA_534 (.A(net638));
 sg13g2_antennanp ANTENNA_535 (.A(net638));
 sg13g2_antennanp ANTENNA_536 (.A(net638));
 sg13g2_antennanp ANTENNA_537 (.A(net638));
 sg13g2_antennanp ANTENNA_538 (.A(net638));
 sg13g2_antennanp ANTENNA_539 (.A(net638));
 sg13g2_antennanp ANTENNA_540 (.A(net639));
 sg13g2_antennanp ANTENNA_541 (.A(net639));
 sg13g2_antennanp ANTENNA_542 (.A(net639));
 sg13g2_antennanp ANTENNA_543 (.A(net639));
 sg13g2_antennanp ANTENNA_544 (.A(net639));
 sg13g2_antennanp ANTENNA_545 (.A(net639));
 sg13g2_antennanp ANTENNA_546 (.A(net639));
 sg13g2_antennanp ANTENNA_547 (.A(net639));
 sg13g2_antennanp ANTENNA_548 (.A(net639));
 sg13g2_antennanp ANTENNA_549 (.A(net639));
 sg13g2_antennanp ANTENNA_550 (.A(net639));
 sg13g2_antennanp ANTENNA_551 (.A(net639));
 sg13g2_antennanp ANTENNA_552 (.A(net639));
 sg13g2_antennanp ANTENNA_553 (.A(net639));
 sg13g2_antennanp ANTENNA_554 (.A(net639));
 sg13g2_antennanp ANTENNA_555 (.A(net639));
 sg13g2_antennanp ANTENNA_556 (.A(net639));
 sg13g2_antennanp ANTENNA_557 (.A(net639));
 sg13g2_antennanp ANTENNA_558 (.A(net639));
 sg13g2_antennanp ANTENNA_559 (.A(net639));
 sg13g2_antennanp ANTENNA_560 (.A(net643));
 sg13g2_antennanp ANTENNA_561 (.A(net643));
 sg13g2_antennanp ANTENNA_562 (.A(net643));
 sg13g2_antennanp ANTENNA_563 (.A(net643));
 sg13g2_antennanp ANTENNA_564 (.A(net643));
 sg13g2_antennanp ANTENNA_565 (.A(net643));
 sg13g2_antennanp ANTENNA_566 (.A(net643));
 sg13g2_antennanp ANTENNA_567 (.A(net643));
 sg13g2_antennanp ANTENNA_568 (.A(net643));
 sg13g2_antennanp ANTENNA_569 (.A(net643));
 sg13g2_antennanp ANTENNA_570 (.A(net643));
 sg13g2_antennanp ANTENNA_571 (.A(net643));
 sg13g2_antennanp ANTENNA_572 (.A(net643));
 sg13g2_antennanp ANTENNA_573 (.A(net667));
 sg13g2_antennanp ANTENNA_574 (.A(net667));
 sg13g2_antennanp ANTENNA_575 (.A(net667));
 sg13g2_antennanp ANTENNA_576 (.A(net667));
 sg13g2_antennanp ANTENNA_577 (.A(net667));
 sg13g2_antennanp ANTENNA_578 (.A(net667));
 sg13g2_antennanp ANTENNA_579 (.A(net667));
 sg13g2_antennanp ANTENNA_580 (.A(net667));
 sg13g2_antennanp ANTENNA_581 (.A(net667));
 sg13g2_antennanp ANTENNA_582 (.A(net667));
 sg13g2_antennanp ANTENNA_583 (.A(net667));
 sg13g2_antennanp ANTENNA_584 (.A(net679));
 sg13g2_antennanp ANTENNA_585 (.A(net679));
 sg13g2_antennanp ANTENNA_586 (.A(net679));
 sg13g2_antennanp ANTENNA_587 (.A(net679));
 sg13g2_antennanp ANTENNA_588 (.A(net679));
 sg13g2_antennanp ANTENNA_589 (.A(net679));
 sg13g2_antennanp ANTENNA_590 (.A(net679));
 sg13g2_antennanp ANTENNA_591 (.A(net679));
 sg13g2_antennanp ANTENNA_592 (.A(net679));
 sg13g2_antennanp ANTENNA_593 (.A(net679));
 sg13g2_antennanp ANTENNA_594 (.A(net679));
 sg13g2_antennanp ANTENNA_595 (.A(net679));
 sg13g2_antennanp ANTENNA_596 (.A(net679));
 sg13g2_antennanp ANTENNA_597 (.A(net679));
 sg13g2_antennanp ANTENNA_598 (.A(net679));
 sg13g2_antennanp ANTENNA_599 (.A(net712));
 sg13g2_antennanp ANTENNA_600 (.A(net712));
 sg13g2_antennanp ANTENNA_601 (.A(net712));
 sg13g2_antennanp ANTENNA_602 (.A(net712));
 sg13g2_antennanp ANTENNA_603 (.A(net712));
 sg13g2_antennanp ANTENNA_604 (.A(net712));
 sg13g2_antennanp ANTENNA_605 (.A(net712));
 sg13g2_antennanp ANTENNA_606 (.A(net712));
 sg13g2_antennanp ANTENNA_607 (.A(net712));
 sg13g2_antennanp ANTENNA_608 (.A(net712));
 sg13g2_antennanp ANTENNA_609 (.A(net712));
 sg13g2_antennanp ANTENNA_610 (.A(net712));
 sg13g2_antennanp ANTENNA_611 (.A(net712));
 sg13g2_antennanp ANTENNA_612 (.A(net712));
 sg13g2_antennanp ANTENNA_613 (.A(net712));
 sg13g2_antennanp ANTENNA_614 (.A(net712));
 sg13g2_antennanp ANTENNA_615 (.A(net712));
 sg13g2_antennanp ANTENNA_616 (.A(net712));
 sg13g2_antennanp ANTENNA_617 (.A(net712));
 sg13g2_antennanp ANTENNA_618 (.A(net712));
 sg13g2_antennanp ANTENNA_619 (.A(net715));
 sg13g2_antennanp ANTENNA_620 (.A(net715));
 sg13g2_antennanp ANTENNA_621 (.A(net715));
 sg13g2_antennanp ANTENNA_622 (.A(net715));
 sg13g2_antennanp ANTENNA_623 (.A(net715));
 sg13g2_antennanp ANTENNA_624 (.A(net715));
 sg13g2_antennanp ANTENNA_625 (.A(net715));
 sg13g2_antennanp ANTENNA_626 (.A(net715));
 sg13g2_antennanp ANTENNA_627 (.A(net715));
 sg13g2_antennanp ANTENNA_628 (.A(net715));
 sg13g2_antennanp ANTENNA_629 (.A(net715));
 sg13g2_antennanp ANTENNA_630 (.A(net715));
 sg13g2_antennanp ANTENNA_631 (.A(net715));
 sg13g2_antennanp ANTENNA_632 (.A(net715));
 sg13g2_antennanp ANTENNA_633 (.A(net715));
 sg13g2_antennanp ANTENNA_634 (.A(net715));
 sg13g2_antennanp ANTENNA_635 (.A(net715));
 sg13g2_antennanp ANTENNA_636 (.A(net715));
 sg13g2_antennanp ANTENNA_637 (.A(net715));
 sg13g2_antennanp ANTENNA_638 (.A(net715));
 sg13g2_antennanp ANTENNA_639 (.A(net780));
 sg13g2_antennanp ANTENNA_640 (.A(net780));
 sg13g2_antennanp ANTENNA_641 (.A(net780));
 sg13g2_antennanp ANTENNA_642 (.A(net780));
 sg13g2_antennanp ANTENNA_643 (.A(net780));
 sg13g2_antennanp ANTENNA_644 (.A(net780));
 sg13g2_antennanp ANTENNA_645 (.A(net780));
 sg13g2_antennanp ANTENNA_646 (.A(net780));
 sg13g2_antennanp ANTENNA_647 (.A(net780));
 sg13g2_antennanp ANTENNA_648 (.A(net780));
 sg13g2_antennanp ANTENNA_649 (.A(net780));
 sg13g2_antennanp ANTENNA_650 (.A(net780));
 sg13g2_antennanp ANTENNA_651 (.A(net780));
 sg13g2_antennanp ANTENNA_652 (.A(net780));
 sg13g2_antennanp ANTENNA_653 (.A(net780));
 sg13g2_antennanp ANTENNA_654 (.A(net780));
 sg13g2_antennanp ANTENNA_655 (.A(net780));
 sg13g2_antennanp ANTENNA_656 (.A(net780));
 sg13g2_antennanp ANTENNA_657 (.A(net780));
 sg13g2_antennanp ANTENNA_658 (.A(net780));
 sg13g2_antennanp ANTENNA_659 (.A(net780));
 sg13g2_antennanp ANTENNA_660 (.A(net796));
 sg13g2_antennanp ANTENNA_661 (.A(net796));
 sg13g2_antennanp ANTENNA_662 (.A(net796));
 sg13g2_antennanp ANTENNA_663 (.A(net796));
 sg13g2_antennanp ANTENNA_664 (.A(net796));
 sg13g2_antennanp ANTENNA_665 (.A(net796));
 sg13g2_antennanp ANTENNA_666 (.A(net796));
 sg13g2_antennanp ANTENNA_667 (.A(net796));
 sg13g2_antennanp ANTENNA_668 (.A(net796));
 sg13g2_antennanp ANTENNA_669 (.A(net796));
 sg13g2_antennanp ANTENNA_670 (.A(net796));
 sg13g2_antennanp ANTENNA_671 (.A(net796));
 sg13g2_antennanp ANTENNA_672 (.A(net796));
 sg13g2_antennanp ANTENNA_673 (.A(net796));
 sg13g2_antennanp ANTENNA_674 (.A(net796));
 sg13g2_antennanp ANTENNA_675 (.A(net796));
 sg13g2_antennanp ANTENNA_676 (.A(net796));
 sg13g2_antennanp ANTENNA_677 (.A(net796));
 sg13g2_antennanp ANTENNA_678 (.A(net796));
 sg13g2_antennanp ANTENNA_679 (.A(net796));
 sg13g2_antennanp ANTENNA_680 (.A(net796));
 sg13g2_antennanp ANTENNA_681 (.A(net796));
 sg13g2_antennanp ANTENNA_682 (.A(net848));
 sg13g2_antennanp ANTENNA_683 (.A(net848));
 sg13g2_antennanp ANTENNA_684 (.A(net848));
 sg13g2_antennanp ANTENNA_685 (.A(net848));
 sg13g2_antennanp ANTENNA_686 (.A(net848));
 sg13g2_antennanp ANTENNA_687 (.A(net848));
 sg13g2_antennanp ANTENNA_688 (.A(net848));
 sg13g2_antennanp ANTENNA_689 (.A(net848));
 sg13g2_antennanp ANTENNA_690 (.A(net848));
 sg13g2_antennanp ANTENNA_691 (.A(net848));
 sg13g2_antennanp ANTENNA_692 (.A(net848));
 sg13g2_antennanp ANTENNA_693 (.A(net848));
 sg13g2_antennanp ANTENNA_694 (.A(net848));
 sg13g2_antennanp ANTENNA_695 (.A(net848));
 sg13g2_antennanp ANTENNA_696 (.A(net848));
 sg13g2_antennanp ANTENNA_697 (.A(net848));
 sg13g2_antennanp ANTENNA_698 (.A(net849));
 sg13g2_antennanp ANTENNA_699 (.A(net849));
 sg13g2_antennanp ANTENNA_700 (.A(net849));
 sg13g2_antennanp ANTENNA_701 (.A(net849));
 sg13g2_antennanp ANTENNA_702 (.A(net849));
 sg13g2_antennanp ANTENNA_703 (.A(net849));
 sg13g2_antennanp ANTENNA_704 (.A(net849));
 sg13g2_antennanp ANTENNA_705 (.A(net849));
 sg13g2_antennanp ANTENNA_706 (.A(net849));
 sg13g2_antennanp ANTENNA_707 (.A(net851));
 sg13g2_antennanp ANTENNA_708 (.A(net851));
 sg13g2_antennanp ANTENNA_709 (.A(net851));
 sg13g2_antennanp ANTENNA_710 (.A(net851));
 sg13g2_antennanp ANTENNA_711 (.A(net851));
 sg13g2_antennanp ANTENNA_712 (.A(net851));
 sg13g2_antennanp ANTENNA_713 (.A(net851));
 sg13g2_antennanp ANTENNA_714 (.A(net851));
 sg13g2_antennanp ANTENNA_715 (.A(net853));
 sg13g2_antennanp ANTENNA_716 (.A(net853));
 sg13g2_antennanp ANTENNA_717 (.A(net853));
 sg13g2_antennanp ANTENNA_718 (.A(net853));
 sg13g2_antennanp ANTENNA_719 (.A(net853));
 sg13g2_antennanp ANTENNA_720 (.A(net853));
 sg13g2_antennanp ANTENNA_721 (.A(net853));
 sg13g2_antennanp ANTENNA_722 (.A(net853));
 sg13g2_antennanp ANTENNA_723 (.A(net853));
 sg13g2_antennanp ANTENNA_724 (.A(net853));
 sg13g2_antennanp ANTENNA_725 (.A(net853));
 sg13g2_antennanp ANTENNA_726 (.A(net853));
 sg13g2_antennanp ANTENNA_727 (.A(net853));
 sg13g2_antennanp ANTENNA_728 (.A(net853));
 sg13g2_antennanp ANTENNA_729 (.A(net853));
 sg13g2_antennanp ANTENNA_730 (.A(net853));
 sg13g2_antennanp ANTENNA_731 (.A(net894));
 sg13g2_antennanp ANTENNA_732 (.A(net894));
 sg13g2_antennanp ANTENNA_733 (.A(net894));
 sg13g2_antennanp ANTENNA_734 (.A(net894));
 sg13g2_antennanp ANTENNA_735 (.A(net894));
 sg13g2_antennanp ANTENNA_736 (.A(net894));
 sg13g2_antennanp ANTENNA_737 (.A(net894));
 sg13g2_antennanp ANTENNA_738 (.A(net894));
 sg13g2_antennanp ANTENNA_739 (.A(net894));
 sg13g2_antennanp ANTENNA_740 (.A(net894));
 sg13g2_antennanp ANTENNA_741 (.A(net894));
 sg13g2_antennanp ANTENNA_742 (.A(net894));
 sg13g2_antennanp ANTENNA_743 (.A(net894));
 sg13g2_antennanp ANTENNA_744 (.A(net894));
 sg13g2_antennanp ANTENNA_745 (.A(net894));
 sg13g2_antennanp ANTENNA_746 (.A(net894));
 sg13g2_antennanp ANTENNA_747 (.A(net894));
 sg13g2_antennanp ANTENNA_748 (.A(net894));
 sg13g2_antennanp ANTENNA_749 (.A(net894));
 sg13g2_antennanp ANTENNA_750 (.A(net894));
 sg13g2_antennanp ANTENNA_751 (.A(net953));
 sg13g2_antennanp ANTENNA_752 (.A(net953));
 sg13g2_antennanp ANTENNA_753 (.A(net953));
 sg13g2_antennanp ANTENNA_754 (.A(net953));
 sg13g2_antennanp ANTENNA_755 (.A(net953));
 sg13g2_antennanp ANTENNA_756 (.A(net953));
 sg13g2_antennanp ANTENNA_757 (.A(net953));
 sg13g2_antennanp ANTENNA_758 (.A(net953));
 sg13g2_antennanp ANTENNA_759 (.A(net953));
 sg13g2_antennanp ANTENNA_760 (.A(net953));
 sg13g2_antennanp ANTENNA_761 (.A(net953));
 sg13g2_antennanp ANTENNA_762 (.A(net953));
 sg13g2_antennanp ANTENNA_763 (.A(net956));
 sg13g2_antennanp ANTENNA_764 (.A(net956));
 sg13g2_antennanp ANTENNA_765 (.A(net956));
 sg13g2_antennanp ANTENNA_766 (.A(net956));
 sg13g2_antennanp ANTENNA_767 (.A(net956));
 sg13g2_antennanp ANTENNA_768 (.A(net956));
 sg13g2_antennanp ANTENNA_769 (.A(net956));
 sg13g2_antennanp ANTENNA_770 (.A(net956));
 sg13g2_antennanp ANTENNA_771 (.A(net956));
 sg13g2_antennanp ANTENNA_772 (.A(net958));
 sg13g2_antennanp ANTENNA_773 (.A(net958));
 sg13g2_antennanp ANTENNA_774 (.A(net958));
 sg13g2_antennanp ANTENNA_775 (.A(net958));
 sg13g2_antennanp ANTENNA_776 (.A(net958));
 sg13g2_antennanp ANTENNA_777 (.A(net958));
 sg13g2_antennanp ANTENNA_778 (.A(net958));
 sg13g2_antennanp ANTENNA_779 (.A(net958));
 sg13g2_antennanp ANTENNA_780 (.A(net983));
 sg13g2_antennanp ANTENNA_781 (.A(net983));
 sg13g2_antennanp ANTENNA_782 (.A(net983));
 sg13g2_antennanp ANTENNA_783 (.A(net983));
 sg13g2_antennanp ANTENNA_784 (.A(net983));
 sg13g2_antennanp ANTENNA_785 (.A(net983));
 sg13g2_antennanp ANTENNA_786 (.A(net983));
 sg13g2_antennanp ANTENNA_787 (.A(net983));
 sg13g2_antennanp ANTENNA_788 (.A(net983));
 sg13g2_antennanp ANTENNA_789 (.A(net983));
 sg13g2_antennanp ANTENNA_790 (.A(net983));
 sg13g2_antennanp ANTENNA_791 (.A(net983));
 sg13g2_antennanp ANTENNA_792 (.A(net983));
 sg13g2_antennanp ANTENNA_793 (.A(net983));
 sg13g2_antennanp ANTENNA_794 (.A(net983));
 sg13g2_antennanp ANTENNA_795 (.A(net983));
 sg13g2_antennanp ANTENNA_796 (.A(net984));
 sg13g2_antennanp ANTENNA_797 (.A(net984));
 sg13g2_antennanp ANTENNA_798 (.A(net984));
 sg13g2_antennanp ANTENNA_799 (.A(net984));
 sg13g2_antennanp ANTENNA_800 (.A(net984));
 sg13g2_antennanp ANTENNA_801 (.A(net984));
 sg13g2_antennanp ANTENNA_802 (.A(net984));
 sg13g2_antennanp ANTENNA_803 (.A(net984));
 sg13g2_antennanp ANTENNA_804 (.A(net986));
 sg13g2_antennanp ANTENNA_805 (.A(net986));
 sg13g2_antennanp ANTENNA_806 (.A(net986));
 sg13g2_antennanp ANTENNA_807 (.A(net986));
 sg13g2_antennanp ANTENNA_808 (.A(net986));
 sg13g2_antennanp ANTENNA_809 (.A(net986));
 sg13g2_antennanp ANTENNA_810 (.A(net986));
 sg13g2_antennanp ANTENNA_811 (.A(net986));
 sg13g2_antennanp ANTENNA_812 (.A(net986));
 sg13g2_antennanp ANTENNA_813 (.A(net986));
 sg13g2_antennanp ANTENNA_814 (.A(net986));
 sg13g2_antennanp ANTENNA_815 (.A(net986));
 sg13g2_antennanp ANTENNA_816 (.A(net986));
 sg13g2_antennanp ANTENNA_817 (.A(net986));
 sg13g2_antennanp ANTENNA_818 (.A(net986));
 sg13g2_antennanp ANTENNA_819 (.A(net986));
 sg13g2_antennanp ANTENNA_820 (.A(net986));
 sg13g2_antennanp ANTENNA_821 (.A(net986));
 sg13g2_antennanp ANTENNA_822 (.A(net986));
 sg13g2_antennanp ANTENNA_823 (.A(net986));
 sg13g2_antennanp ANTENNA_824 (.A(net986));
 sg13g2_antennanp ANTENNA_825 (.A(net991));
 sg13g2_antennanp ANTENNA_826 (.A(net991));
 sg13g2_antennanp ANTENNA_827 (.A(net991));
 sg13g2_antennanp ANTENNA_828 (.A(net991));
 sg13g2_antennanp ANTENNA_829 (.A(net991));
 sg13g2_antennanp ANTENNA_830 (.A(net991));
 sg13g2_antennanp ANTENNA_831 (.A(net991));
 sg13g2_antennanp ANTENNA_832 (.A(net991));
 sg13g2_antennanp ANTENNA_833 (.A(net991));
 sg13g2_antennanp ANTENNA_834 (.A(net1038));
 sg13g2_antennanp ANTENNA_835 (.A(net1038));
 sg13g2_antennanp ANTENNA_836 (.A(net1038));
 sg13g2_antennanp ANTENNA_837 (.A(net1038));
 sg13g2_antennanp ANTENNA_838 (.A(net1038));
 sg13g2_antennanp ANTENNA_839 (.A(net1038));
 sg13g2_antennanp ANTENNA_840 (.A(net1038));
 sg13g2_antennanp ANTENNA_841 (.A(net1038));
 sg13g2_antennanp ANTENNA_842 (.A(net1038));
 sg13g2_antennanp ANTENNA_843 (.A(net1038));
 sg13g2_antennanp ANTENNA_844 (.A(net1038));
 sg13g2_antennanp ANTENNA_845 (.A(net1038));
 sg13g2_antennanp ANTENNA_846 (.A(net1038));
 sg13g2_antennanp ANTENNA_847 (.A(net1038));
 sg13g2_antennanp ANTENNA_848 (.A(net1038));
 sg13g2_antennanp ANTENNA_849 (.A(net1038));
 sg13g2_antennanp ANTENNA_850 (.A(net1038));
 sg13g2_antennanp ANTENNA_851 (.A(net1038));
 sg13g2_antennanp ANTENNA_852 (.A(net1038));
 sg13g2_antennanp ANTENNA_853 (.A(net1038));
 sg13g2_antennanp ANTENNA_854 (.A(net1038));
 sg13g2_antennanp ANTENNA_855 (.A(net1038));
 sg13g2_antennanp ANTENNA_856 (.A(net1038));
 sg13g2_antennanp ANTENNA_857 (.A(net1038));
 sg13g2_antennanp ANTENNA_858 (.A(net1038));
 sg13g2_antennanp ANTENNA_859 (.A(net1038));
 sg13g2_antennanp ANTENNA_860 (.A(net1038));
 sg13g2_antennanp ANTENNA_861 (.A(net1038));
 sg13g2_antennanp ANTENNA_862 (.A(net1038));
 sg13g2_antennanp ANTENNA_863 (.A(net1038));
 sg13g2_antennanp ANTENNA_864 (.A(net1056));
 sg13g2_antennanp ANTENNA_865 (.A(net1056));
 sg13g2_antennanp ANTENNA_866 (.A(net1056));
 sg13g2_antennanp ANTENNA_867 (.A(net1056));
 sg13g2_antennanp ANTENNA_868 (.A(net1056));
 sg13g2_antennanp ANTENNA_869 (.A(net1056));
 sg13g2_antennanp ANTENNA_870 (.A(net1056));
 sg13g2_antennanp ANTENNA_871 (.A(net1056));
 sg13g2_antennanp ANTENNA_872 (.A(net1056));
 sg13g2_antennanp ANTENNA_873 (.A(net1056));
 sg13g2_antennanp ANTENNA_874 (.A(net1056));
 sg13g2_antennanp ANTENNA_875 (.A(net1056));
 sg13g2_antennanp ANTENNA_876 (.A(_00237_));
 sg13g2_antennanp ANTENNA_877 (.A(_00789_));
 sg13g2_antennanp ANTENNA_878 (.A(_00798_));
 sg13g2_antennanp ANTENNA_879 (.A(_00930_));
 sg13g2_antennanp ANTENNA_880 (.A(_02788_));
 sg13g2_antennanp ANTENNA_881 (.A(_02788_));
 sg13g2_antennanp ANTENNA_882 (.A(_02788_));
 sg13g2_antennanp ANTENNA_883 (.A(_02788_));
 sg13g2_antennanp ANTENNA_884 (.A(_02788_));
 sg13g2_antennanp ANTENNA_885 (.A(_02788_));
 sg13g2_antennanp ANTENNA_886 (.A(_02788_));
 sg13g2_antennanp ANTENNA_887 (.A(_02788_));
 sg13g2_antennanp ANTENNA_888 (.A(_02788_));
 sg13g2_antennanp ANTENNA_889 (.A(_02797_));
 sg13g2_antennanp ANTENNA_890 (.A(_02797_));
 sg13g2_antennanp ANTENNA_891 (.A(_02797_));
 sg13g2_antennanp ANTENNA_892 (.A(_02797_));
 sg13g2_antennanp ANTENNA_893 (.A(_02797_));
 sg13g2_antennanp ANTENNA_894 (.A(_02797_));
 sg13g2_antennanp ANTENNA_895 (.A(_02797_));
 sg13g2_antennanp ANTENNA_896 (.A(_02797_));
 sg13g2_antennanp ANTENNA_897 (.A(_02797_));
 sg13g2_antennanp ANTENNA_898 (.A(_02801_));
 sg13g2_antennanp ANTENNA_899 (.A(_02801_));
 sg13g2_antennanp ANTENNA_900 (.A(_02801_));
 sg13g2_antennanp ANTENNA_901 (.A(_02801_));
 sg13g2_antennanp ANTENNA_902 (.A(_02801_));
 sg13g2_antennanp ANTENNA_903 (.A(_02801_));
 sg13g2_antennanp ANTENNA_904 (.A(_02801_));
 sg13g2_antennanp ANTENNA_905 (.A(_02801_));
 sg13g2_antennanp ANTENNA_906 (.A(_02801_));
 sg13g2_antennanp ANTENNA_907 (.A(_02805_));
 sg13g2_antennanp ANTENNA_908 (.A(_02805_));
 sg13g2_antennanp ANTENNA_909 (.A(_02805_));
 sg13g2_antennanp ANTENNA_910 (.A(_02805_));
 sg13g2_antennanp ANTENNA_911 (.A(_02805_));
 sg13g2_antennanp ANTENNA_912 (.A(_02805_));
 sg13g2_antennanp ANTENNA_913 (.A(_02805_));
 sg13g2_antennanp ANTENNA_914 (.A(_02805_));
 sg13g2_antennanp ANTENNA_915 (.A(_02805_));
 sg13g2_antennanp ANTENNA_916 (.A(_02908_));
 sg13g2_antennanp ANTENNA_917 (.A(_02908_));
 sg13g2_antennanp ANTENNA_918 (.A(_02908_));
 sg13g2_antennanp ANTENNA_919 (.A(_02908_));
 sg13g2_antennanp ANTENNA_920 (.A(_02908_));
 sg13g2_antennanp ANTENNA_921 (.A(_02908_));
 sg13g2_antennanp ANTENNA_922 (.A(_02917_));
 sg13g2_antennanp ANTENNA_923 (.A(_02917_));
 sg13g2_antennanp ANTENNA_924 (.A(_02917_));
 sg13g2_antennanp ANTENNA_925 (.A(_02917_));
 sg13g2_antennanp ANTENNA_926 (.A(_02918_));
 sg13g2_antennanp ANTENNA_927 (.A(_02918_));
 sg13g2_antennanp ANTENNA_928 (.A(_02918_));
 sg13g2_antennanp ANTENNA_929 (.A(_02919_));
 sg13g2_antennanp ANTENNA_930 (.A(_02919_));
 sg13g2_antennanp ANTENNA_931 (.A(_02919_));
 sg13g2_antennanp ANTENNA_932 (.A(_02919_));
 sg13g2_antennanp ANTENNA_933 (.A(_02920_));
 sg13g2_antennanp ANTENNA_934 (.A(_02920_));
 sg13g2_antennanp ANTENNA_935 (.A(_02920_));
 sg13g2_antennanp ANTENNA_936 (.A(_02920_));
 sg13g2_antennanp ANTENNA_937 (.A(_02920_));
 sg13g2_antennanp ANTENNA_938 (.A(_02920_));
 sg13g2_antennanp ANTENNA_939 (.A(_02920_));
 sg13g2_antennanp ANTENNA_940 (.A(_02920_));
 sg13g2_antennanp ANTENNA_941 (.A(_02920_));
 sg13g2_antennanp ANTENNA_942 (.A(_02920_));
 sg13g2_antennanp ANTENNA_943 (.A(_02922_));
 sg13g2_antennanp ANTENNA_944 (.A(_02922_));
 sg13g2_antennanp ANTENNA_945 (.A(_02922_));
 sg13g2_antennanp ANTENNA_946 (.A(_02927_));
 sg13g2_antennanp ANTENNA_947 (.A(_02927_));
 sg13g2_antennanp ANTENNA_948 (.A(_02927_));
 sg13g2_antennanp ANTENNA_949 (.A(_02927_));
 sg13g2_antennanp ANTENNA_950 (.A(_02927_));
 sg13g2_antennanp ANTENNA_951 (.A(_02927_));
 sg13g2_antennanp ANTENNA_952 (.A(_02927_));
 sg13g2_antennanp ANTENNA_953 (.A(_02927_));
 sg13g2_antennanp ANTENNA_954 (.A(_02927_));
 sg13g2_antennanp ANTENNA_955 (.A(_02927_));
 sg13g2_antennanp ANTENNA_956 (.A(_02936_));
 sg13g2_antennanp ANTENNA_957 (.A(_02936_));
 sg13g2_antennanp ANTENNA_958 (.A(_02936_));
 sg13g2_antennanp ANTENNA_959 (.A(_03293_));
 sg13g2_antennanp ANTENNA_960 (.A(_03323_));
 sg13g2_antennanp ANTENNA_961 (.A(_03324_));
 sg13g2_antennanp ANTENNA_962 (.A(_03329_));
 sg13g2_antennanp ANTENNA_963 (.A(_03397_));
 sg13g2_antennanp ANTENNA_964 (.A(_03397_));
 sg13g2_antennanp ANTENNA_965 (.A(_03397_));
 sg13g2_antennanp ANTENNA_966 (.A(_03397_));
 sg13g2_antennanp ANTENNA_967 (.A(_03697_));
 sg13g2_antennanp ANTENNA_968 (.A(_03697_));
 sg13g2_antennanp ANTENNA_969 (.A(_03697_));
 sg13g2_antennanp ANTENNA_970 (.A(_05114_));
 sg13g2_antennanp ANTENNA_971 (.A(_05142_));
 sg13g2_antennanp ANTENNA_972 (.A(_05173_));
 sg13g2_antennanp ANTENNA_973 (.A(_05204_));
 sg13g2_antennanp ANTENNA_974 (.A(_05236_));
 sg13g2_antennanp ANTENNA_975 (.A(_05248_));
 sg13g2_antennanp ANTENNA_976 (.A(_05255_));
 sg13g2_antennanp ANTENNA_977 (.A(_05407_));
 sg13g2_antennanp ANTENNA_978 (.A(_05412_));
 sg13g2_antennanp ANTENNA_979 (.A(_05477_));
 sg13g2_antennanp ANTENNA_980 (.A(_05556_));
 sg13g2_antennanp ANTENNA_981 (.A(_05681_));
 sg13g2_antennanp ANTENNA_982 (.A(_05695_));
 sg13g2_antennanp ANTENNA_983 (.A(_05708_));
 sg13g2_antennanp ANTENNA_984 (.A(_05735_));
 sg13g2_antennanp ANTENNA_985 (.A(_06655_));
 sg13g2_antennanp ANTENNA_986 (.A(_06655_));
 sg13g2_antennanp ANTENNA_987 (.A(_06655_));
 sg13g2_antennanp ANTENNA_988 (.A(_06655_));
 sg13g2_antennanp ANTENNA_989 (.A(_07439_));
 sg13g2_antennanp ANTENNA_990 (.A(_07476_));
 sg13g2_antennanp ANTENNA_991 (.A(_07476_));
 sg13g2_antennanp ANTENNA_992 (.A(_07476_));
 sg13g2_antennanp ANTENNA_993 (.A(_07476_));
 sg13g2_antennanp ANTENNA_994 (.A(_07476_));
 sg13g2_antennanp ANTENNA_995 (.A(_07476_));
 sg13g2_antennanp ANTENNA_996 (.A(_07476_));
 sg13g2_antennanp ANTENNA_997 (.A(_07476_));
 sg13g2_antennanp ANTENNA_998 (.A(_07476_));
 sg13g2_antennanp ANTENNA_999 (.A(_07476_));
 sg13g2_antennanp ANTENNA_1000 (.A(_07737_));
 sg13g2_antennanp ANTENNA_1001 (.A(_07737_));
 sg13g2_antennanp ANTENNA_1002 (.A(_07737_));
 sg13g2_antennanp ANTENNA_1003 (.A(_07737_));
 sg13g2_antennanp ANTENNA_1004 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1005 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1006 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1007 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1008 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1009 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1010 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1011 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1012 (.A(_08159_));
 sg13g2_antennanp ANTENNA_1013 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1014 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1015 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1016 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1017 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1018 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1019 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1020 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1021 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1022 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1023 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1024 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1025 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1026 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1027 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1028 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1029 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1030 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1031 (.A(_08476_));
 sg13g2_antennanp ANTENNA_1032 (.A(_08498_));
 sg13g2_antennanp ANTENNA_1033 (.A(_08498_));
 sg13g2_antennanp ANTENNA_1034 (.A(_08498_));
 sg13g2_antennanp ANTENNA_1035 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1036 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1037 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1038 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1039 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1040 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1041 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1042 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1043 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1044 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1045 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1046 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1047 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1048 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1049 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1050 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1051 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1052 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1053 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1054 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1055 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1056 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1057 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1058 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1059 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1060 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1061 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1062 (.A(_08583_));
 sg13g2_antennanp ANTENNA_1063 (.A(_08584_));
 sg13g2_antennanp ANTENNA_1064 (.A(_08584_));
 sg13g2_antennanp ANTENNA_1065 (.A(_08607_));
 sg13g2_antennanp ANTENNA_1066 (.A(_08607_));
 sg13g2_antennanp ANTENNA_1067 (.A(_08607_));
 sg13g2_antennanp ANTENNA_1068 (.A(_08627_));
 sg13g2_antennanp ANTENNA_1069 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1070 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1071 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1072 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1073 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1074 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1075 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1076 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1077 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1078 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1079 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1080 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1081 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1082 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1083 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1084 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1085 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1086 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1087 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1088 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1089 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1090 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1091 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1092 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1093 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1094 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1095 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1096 (.A(_09082_));
 sg13g2_antennanp ANTENNA_1097 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1098 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1099 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1100 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1101 (.A(_09095_));
 sg13g2_antennanp ANTENNA_1102 (.A(_09095_));
 sg13g2_antennanp ANTENNA_1103 (.A(_09102_));
 sg13g2_antennanp ANTENNA_1104 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1105 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1106 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1107 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1108 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1109 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1110 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1111 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1112 (.A(_09119_));
 sg13g2_antennanp ANTENNA_1113 (.A(_09123_));
 sg13g2_antennanp ANTENNA_1114 (.A(_09123_));
 sg13g2_antennanp ANTENNA_1115 (.A(_09123_));
 sg13g2_antennanp ANTENNA_1116 (.A(_09125_));
 sg13g2_antennanp ANTENNA_1117 (.A(_09125_));
 sg13g2_antennanp ANTENNA_1118 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1119 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1120 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1121 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1122 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1123 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1124 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1125 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1126 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1127 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1128 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1129 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1130 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1131 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1132 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1133 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1134 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1135 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1136 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1137 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1138 (.A(_09246_));
 sg13g2_antennanp ANTENNA_1139 (.A(_09248_));
 sg13g2_antennanp ANTENNA_1140 (.A(_09312_));
 sg13g2_antennanp ANTENNA_1141 (.A(_09315_));
 sg13g2_antennanp ANTENNA_1142 (.A(_09341_));
 sg13g2_antennanp ANTENNA_1143 (.A(_09443_));
 sg13g2_antennanp ANTENNA_1144 (.A(_09466_));
 sg13g2_antennanp ANTENNA_1145 (.A(_09492_));
 sg13g2_antennanp ANTENNA_1146 (.A(_09514_));
 sg13g2_antennanp ANTENNA_1147 (.A(_09536_));
 sg13g2_antennanp ANTENNA_1148 (.A(_09561_));
 sg13g2_antennanp ANTENNA_1149 (.A(_09585_));
 sg13g2_antennanp ANTENNA_1150 (.A(_09608_));
 sg13g2_antennanp ANTENNA_1151 (.A(_09608_));
 sg13g2_antennanp ANTENNA_1152 (.A(_09630_));
 sg13g2_antennanp ANTENNA_1153 (.A(_09759_));
 sg13g2_antennanp ANTENNA_1154 (.A(_09943_));
 sg13g2_antennanp ANTENNA_1155 (.A(_09943_));
 sg13g2_antennanp ANTENNA_1156 (.A(_09943_));
 sg13g2_antennanp ANTENNA_1157 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1158 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1159 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1160 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1161 (.A(_10078_));
 sg13g2_antennanp ANTENNA_1162 (.A(_10078_));
 sg13g2_antennanp ANTENNA_1163 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1164 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1165 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1166 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1167 (.A(_10758_));
 sg13g2_antennanp ANTENNA_1168 (.A(_10758_));
 sg13g2_antennanp ANTENNA_1169 (.A(_10758_));
 sg13g2_antennanp ANTENNA_1170 (.A(_10758_));
 sg13g2_antennanp ANTENNA_1171 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1172 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1173 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1174 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1175 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1176 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1177 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1178 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1179 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1180 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1181 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1182 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1183 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1184 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1185 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1186 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1187 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1188 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1189 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1190 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1191 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1192 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1193 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1194 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1195 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1196 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1197 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1198 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1199 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1200 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1201 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1202 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1203 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1204 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1205 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1206 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1207 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1208 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1209 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1210 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1211 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1212 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1213 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1214 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1215 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1216 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1217 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1218 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1219 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1220 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1221 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1222 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1223 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1224 (.A(clk));
 sg13g2_antennanp ANTENNA_1225 (.A(clk));
 sg13g2_antennanp ANTENNA_1226 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1227 (.A(net3));
 sg13g2_antennanp ANTENNA_1228 (.A(net3));
 sg13g2_antennanp ANTENNA_1229 (.A(net3));
 sg13g2_antennanp ANTENNA_1230 (.A(net19));
 sg13g2_antennanp ANTENNA_1231 (.A(net19));
 sg13g2_antennanp ANTENNA_1232 (.A(net151));
 sg13g2_antennanp ANTENNA_1233 (.A(net151));
 sg13g2_antennanp ANTENNA_1234 (.A(net151));
 sg13g2_antennanp ANTENNA_1235 (.A(net151));
 sg13g2_antennanp ANTENNA_1236 (.A(net151));
 sg13g2_antennanp ANTENNA_1237 (.A(net151));
 sg13g2_antennanp ANTENNA_1238 (.A(net151));
 sg13g2_antennanp ANTENNA_1239 (.A(net151));
 sg13g2_antennanp ANTENNA_1240 (.A(net151));
 sg13g2_antennanp ANTENNA_1241 (.A(net366));
 sg13g2_antennanp ANTENNA_1242 (.A(net366));
 sg13g2_antennanp ANTENNA_1243 (.A(net366));
 sg13g2_antennanp ANTENNA_1244 (.A(net366));
 sg13g2_antennanp ANTENNA_1245 (.A(net366));
 sg13g2_antennanp ANTENNA_1246 (.A(net366));
 sg13g2_antennanp ANTENNA_1247 (.A(net366));
 sg13g2_antennanp ANTENNA_1248 (.A(net366));
 sg13g2_antennanp ANTENNA_1249 (.A(net366));
 sg13g2_antennanp ANTENNA_1250 (.A(net366));
 sg13g2_antennanp ANTENNA_1251 (.A(net366));
 sg13g2_antennanp ANTENNA_1252 (.A(net366));
 sg13g2_antennanp ANTENNA_1253 (.A(net468));
 sg13g2_antennanp ANTENNA_1254 (.A(net468));
 sg13g2_antennanp ANTENNA_1255 (.A(net468));
 sg13g2_antennanp ANTENNA_1256 (.A(net468));
 sg13g2_antennanp ANTENNA_1257 (.A(net468));
 sg13g2_antennanp ANTENNA_1258 (.A(net468));
 sg13g2_antennanp ANTENNA_1259 (.A(net468));
 sg13g2_antennanp ANTENNA_1260 (.A(net468));
 sg13g2_antennanp ANTENNA_1261 (.A(net468));
 sg13g2_antennanp ANTENNA_1262 (.A(net594));
 sg13g2_antennanp ANTENNA_1263 (.A(net594));
 sg13g2_antennanp ANTENNA_1264 (.A(net594));
 sg13g2_antennanp ANTENNA_1265 (.A(net594));
 sg13g2_antennanp ANTENNA_1266 (.A(net594));
 sg13g2_antennanp ANTENNA_1267 (.A(net594));
 sg13g2_antennanp ANTENNA_1268 (.A(net594));
 sg13g2_antennanp ANTENNA_1269 (.A(net594));
 sg13g2_antennanp ANTENNA_1270 (.A(net638));
 sg13g2_antennanp ANTENNA_1271 (.A(net638));
 sg13g2_antennanp ANTENNA_1272 (.A(net638));
 sg13g2_antennanp ANTENNA_1273 (.A(net638));
 sg13g2_antennanp ANTENNA_1274 (.A(net638));
 sg13g2_antennanp ANTENNA_1275 (.A(net638));
 sg13g2_antennanp ANTENNA_1276 (.A(net638));
 sg13g2_antennanp ANTENNA_1277 (.A(net638));
 sg13g2_antennanp ANTENNA_1278 (.A(net638));
 sg13g2_antennanp ANTENNA_1279 (.A(net643));
 sg13g2_antennanp ANTENNA_1280 (.A(net643));
 sg13g2_antennanp ANTENNA_1281 (.A(net643));
 sg13g2_antennanp ANTENNA_1282 (.A(net643));
 sg13g2_antennanp ANTENNA_1283 (.A(net643));
 sg13g2_antennanp ANTENNA_1284 (.A(net643));
 sg13g2_antennanp ANTENNA_1285 (.A(net643));
 sg13g2_antennanp ANTENNA_1286 (.A(net643));
 sg13g2_antennanp ANTENNA_1287 (.A(net643));
 sg13g2_antennanp ANTENNA_1288 (.A(net643));
 sg13g2_antennanp ANTENNA_1289 (.A(net643));
 sg13g2_antennanp ANTENNA_1290 (.A(net643));
 sg13g2_antennanp ANTENNA_1291 (.A(net643));
 sg13g2_antennanp ANTENNA_1292 (.A(net643));
 sg13g2_antennanp ANTENNA_1293 (.A(net643));
 sg13g2_antennanp ANTENNA_1294 (.A(net643));
 sg13g2_antennanp ANTENNA_1295 (.A(net643));
 sg13g2_antennanp ANTENNA_1296 (.A(net643));
 sg13g2_antennanp ANTENNA_1297 (.A(net667));
 sg13g2_antennanp ANTENNA_1298 (.A(net667));
 sg13g2_antennanp ANTENNA_1299 (.A(net667));
 sg13g2_antennanp ANTENNA_1300 (.A(net667));
 sg13g2_antennanp ANTENNA_1301 (.A(net667));
 sg13g2_antennanp ANTENNA_1302 (.A(net667));
 sg13g2_antennanp ANTENNA_1303 (.A(net667));
 sg13g2_antennanp ANTENNA_1304 (.A(net667));
 sg13g2_antennanp ANTENNA_1305 (.A(net667));
 sg13g2_antennanp ANTENNA_1306 (.A(net667));
 sg13g2_antennanp ANTENNA_1307 (.A(net667));
 sg13g2_antennanp ANTENNA_1308 (.A(net667));
 sg13g2_antennanp ANTENNA_1309 (.A(net667));
 sg13g2_antennanp ANTENNA_1310 (.A(net667));
 sg13g2_antennanp ANTENNA_1311 (.A(net667));
 sg13g2_antennanp ANTENNA_1312 (.A(net667));
 sg13g2_antennanp ANTENNA_1313 (.A(net679));
 sg13g2_antennanp ANTENNA_1314 (.A(net679));
 sg13g2_antennanp ANTENNA_1315 (.A(net679));
 sg13g2_antennanp ANTENNA_1316 (.A(net679));
 sg13g2_antennanp ANTENNA_1317 (.A(net679));
 sg13g2_antennanp ANTENNA_1318 (.A(net679));
 sg13g2_antennanp ANTENNA_1319 (.A(net679));
 sg13g2_antennanp ANTENNA_1320 (.A(net679));
 sg13g2_antennanp ANTENNA_1321 (.A(net679));
 sg13g2_antennanp ANTENNA_1322 (.A(net679));
 sg13g2_antennanp ANTENNA_1323 (.A(net679));
 sg13g2_antennanp ANTENNA_1324 (.A(net679));
 sg13g2_antennanp ANTENNA_1325 (.A(net679));
 sg13g2_antennanp ANTENNA_1326 (.A(net679));
 sg13g2_antennanp ANTENNA_1327 (.A(net679));
 sg13g2_antennanp ANTENNA_1328 (.A(net780));
 sg13g2_antennanp ANTENNA_1329 (.A(net780));
 sg13g2_antennanp ANTENNA_1330 (.A(net780));
 sg13g2_antennanp ANTENNA_1331 (.A(net780));
 sg13g2_antennanp ANTENNA_1332 (.A(net780));
 sg13g2_antennanp ANTENNA_1333 (.A(net780));
 sg13g2_antennanp ANTENNA_1334 (.A(net780));
 sg13g2_antennanp ANTENNA_1335 (.A(net780));
 sg13g2_antennanp ANTENNA_1336 (.A(net780));
 sg13g2_antennanp ANTENNA_1337 (.A(net848));
 sg13g2_antennanp ANTENNA_1338 (.A(net848));
 sg13g2_antennanp ANTENNA_1339 (.A(net848));
 sg13g2_antennanp ANTENNA_1340 (.A(net848));
 sg13g2_antennanp ANTENNA_1341 (.A(net848));
 sg13g2_antennanp ANTENNA_1342 (.A(net848));
 sg13g2_antennanp ANTENNA_1343 (.A(net848));
 sg13g2_antennanp ANTENNA_1344 (.A(net848));
 sg13g2_antennanp ANTENNA_1345 (.A(net848));
 sg13g2_antennanp ANTENNA_1346 (.A(net851));
 sg13g2_antennanp ANTENNA_1347 (.A(net851));
 sg13g2_antennanp ANTENNA_1348 (.A(net851));
 sg13g2_antennanp ANTENNA_1349 (.A(net851));
 sg13g2_antennanp ANTENNA_1350 (.A(net851));
 sg13g2_antennanp ANTENNA_1351 (.A(net851));
 sg13g2_antennanp ANTENNA_1352 (.A(net851));
 sg13g2_antennanp ANTENNA_1353 (.A(net851));
 sg13g2_antennanp ANTENNA_1354 (.A(net853));
 sg13g2_antennanp ANTENNA_1355 (.A(net853));
 sg13g2_antennanp ANTENNA_1356 (.A(net853));
 sg13g2_antennanp ANTENNA_1357 (.A(net853));
 sg13g2_antennanp ANTENNA_1358 (.A(net853));
 sg13g2_antennanp ANTENNA_1359 (.A(net853));
 sg13g2_antennanp ANTENNA_1360 (.A(net853));
 sg13g2_antennanp ANTENNA_1361 (.A(net853));
 sg13g2_antennanp ANTENNA_1362 (.A(net853));
 sg13g2_antennanp ANTENNA_1363 (.A(net853));
 sg13g2_antennanp ANTENNA_1364 (.A(net853));
 sg13g2_antennanp ANTENNA_1365 (.A(net853));
 sg13g2_antennanp ANTENNA_1366 (.A(net853));
 sg13g2_antennanp ANTENNA_1367 (.A(net853));
 sg13g2_antennanp ANTENNA_1368 (.A(net853));
 sg13g2_antennanp ANTENNA_1369 (.A(net853));
 sg13g2_antennanp ANTENNA_1370 (.A(net853));
 sg13g2_antennanp ANTENNA_1371 (.A(net853));
 sg13g2_antennanp ANTENNA_1372 (.A(net853));
 sg13g2_antennanp ANTENNA_1373 (.A(net853));
 sg13g2_antennanp ANTENNA_1374 (.A(net853));
 sg13g2_antennanp ANTENNA_1375 (.A(net853));
 sg13g2_antennanp ANTENNA_1376 (.A(net894));
 sg13g2_antennanp ANTENNA_1377 (.A(net894));
 sg13g2_antennanp ANTENNA_1378 (.A(net894));
 sg13g2_antennanp ANTENNA_1379 (.A(net894));
 sg13g2_antennanp ANTENNA_1380 (.A(net894));
 sg13g2_antennanp ANTENNA_1381 (.A(net894));
 sg13g2_antennanp ANTENNA_1382 (.A(net894));
 sg13g2_antennanp ANTENNA_1383 (.A(net894));
 sg13g2_antennanp ANTENNA_1384 (.A(net894));
 sg13g2_antennanp ANTENNA_1385 (.A(net906));
 sg13g2_antennanp ANTENNA_1386 (.A(net906));
 sg13g2_antennanp ANTENNA_1387 (.A(net906));
 sg13g2_antennanp ANTENNA_1388 (.A(net906));
 sg13g2_antennanp ANTENNA_1389 (.A(net906));
 sg13g2_antennanp ANTENNA_1390 (.A(net906));
 sg13g2_antennanp ANTENNA_1391 (.A(net906));
 sg13g2_antennanp ANTENNA_1392 (.A(net906));
 sg13g2_antennanp ANTENNA_1393 (.A(net906));
 sg13g2_antennanp ANTENNA_1394 (.A(net956));
 sg13g2_antennanp ANTENNA_1395 (.A(net956));
 sg13g2_antennanp ANTENNA_1396 (.A(net956));
 sg13g2_antennanp ANTENNA_1397 (.A(net956));
 sg13g2_antennanp ANTENNA_1398 (.A(net956));
 sg13g2_antennanp ANTENNA_1399 (.A(net956));
 sg13g2_antennanp ANTENNA_1400 (.A(net956));
 sg13g2_antennanp ANTENNA_1401 (.A(net956));
 sg13g2_antennanp ANTENNA_1402 (.A(net956));
 sg13g2_antennanp ANTENNA_1403 (.A(net956));
 sg13g2_antennanp ANTENNA_1404 (.A(net956));
 sg13g2_antennanp ANTENNA_1405 (.A(net956));
 sg13g2_antennanp ANTENNA_1406 (.A(net956));
 sg13g2_antennanp ANTENNA_1407 (.A(net984));
 sg13g2_antennanp ANTENNA_1408 (.A(net984));
 sg13g2_antennanp ANTENNA_1409 (.A(net984));
 sg13g2_antennanp ANTENNA_1410 (.A(net984));
 sg13g2_antennanp ANTENNA_1411 (.A(net984));
 sg13g2_antennanp ANTENNA_1412 (.A(net984));
 sg13g2_antennanp ANTENNA_1413 (.A(net984));
 sg13g2_antennanp ANTENNA_1414 (.A(net984));
 sg13g2_antennanp ANTENNA_1415 (.A(net984));
 sg13g2_antennanp ANTENNA_1416 (.A(net984));
 sg13g2_antennanp ANTENNA_1417 (.A(net984));
 sg13g2_antennanp ANTENNA_1418 (.A(net984));
 sg13g2_antennanp ANTENNA_1419 (.A(net984));
 sg13g2_antennanp ANTENNA_1420 (.A(net984));
 sg13g2_antennanp ANTENNA_1421 (.A(net984));
 sg13g2_antennanp ANTENNA_1422 (.A(net984));
 sg13g2_antennanp ANTENNA_1423 (.A(net984));
 sg13g2_antennanp ANTENNA_1424 (.A(net984));
 sg13g2_antennanp ANTENNA_1425 (.A(net984));
 sg13g2_antennanp ANTENNA_1426 (.A(net984));
 sg13g2_antennanp ANTENNA_1427 (.A(net986));
 sg13g2_antennanp ANTENNA_1428 (.A(net986));
 sg13g2_antennanp ANTENNA_1429 (.A(net986));
 sg13g2_antennanp ANTENNA_1430 (.A(net986));
 sg13g2_antennanp ANTENNA_1431 (.A(net986));
 sg13g2_antennanp ANTENNA_1432 (.A(net986));
 sg13g2_antennanp ANTENNA_1433 (.A(net986));
 sg13g2_antennanp ANTENNA_1434 (.A(net986));
 sg13g2_antennanp ANTENNA_1435 (.A(net991));
 sg13g2_antennanp ANTENNA_1436 (.A(net991));
 sg13g2_antennanp ANTENNA_1437 (.A(net991));
 sg13g2_antennanp ANTENNA_1438 (.A(net991));
 sg13g2_antennanp ANTENNA_1439 (.A(net991));
 sg13g2_antennanp ANTENNA_1440 (.A(net991));
 sg13g2_antennanp ANTENNA_1441 (.A(net991));
 sg13g2_antennanp ANTENNA_1442 (.A(net991));
 sg13g2_antennanp ANTENNA_1443 (.A(net991));
 sg13g2_antennanp ANTENNA_1444 (.A(net1038));
 sg13g2_antennanp ANTENNA_1445 (.A(net1038));
 sg13g2_antennanp ANTENNA_1446 (.A(net1038));
 sg13g2_antennanp ANTENNA_1447 (.A(net1038));
 sg13g2_antennanp ANTENNA_1448 (.A(net1038));
 sg13g2_antennanp ANTENNA_1449 (.A(net1038));
 sg13g2_antennanp ANTENNA_1450 (.A(net1038));
 sg13g2_antennanp ANTENNA_1451 (.A(net1038));
 sg13g2_antennanp ANTENNA_1452 (.A(_00237_));
 sg13g2_antennanp ANTENNA_1453 (.A(_00789_));
 sg13g2_antennanp ANTENNA_1454 (.A(_00798_));
 sg13g2_antennanp ANTENNA_1455 (.A(_00930_));
 sg13g2_antennanp ANTENNA_1456 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1457 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1458 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1459 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1460 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1461 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1462 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1463 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1464 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1465 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1466 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1467 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1468 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1469 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1470 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1471 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1472 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1473 (.A(_02797_));
 sg13g2_antennanp ANTENNA_1474 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1475 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1476 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1477 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1478 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1479 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1480 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1481 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1482 (.A(_02801_));
 sg13g2_antennanp ANTENNA_1483 (.A(_02908_));
 sg13g2_antennanp ANTENNA_1484 (.A(_02908_));
 sg13g2_antennanp ANTENNA_1485 (.A(_02908_));
 sg13g2_antennanp ANTENNA_1486 (.A(_02908_));
 sg13g2_antennanp ANTENNA_1487 (.A(_02908_));
 sg13g2_antennanp ANTENNA_1488 (.A(_02908_));
 sg13g2_antennanp ANTENNA_1489 (.A(_02917_));
 sg13g2_antennanp ANTENNA_1490 (.A(_02917_));
 sg13g2_antennanp ANTENNA_1491 (.A(_02917_));
 sg13g2_antennanp ANTENNA_1492 (.A(_02917_));
 sg13g2_antennanp ANTENNA_1493 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1494 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1495 (.A(_02918_));
 sg13g2_antennanp ANTENNA_1496 (.A(_02919_));
 sg13g2_antennanp ANTENNA_1497 (.A(_02919_));
 sg13g2_antennanp ANTENNA_1498 (.A(_02919_));
 sg13g2_antennanp ANTENNA_1499 (.A(_02919_));
 sg13g2_antennanp ANTENNA_1500 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1501 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1502 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1503 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1504 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1505 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1506 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1507 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1508 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1509 (.A(_02920_));
 sg13g2_antennanp ANTENNA_1510 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1511 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1512 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1513 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1514 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1515 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1516 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1517 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1518 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1519 (.A(_02922_));
 sg13g2_antennanp ANTENNA_1520 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1521 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1522 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1523 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1524 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1525 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1526 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1527 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1528 (.A(_02927_));
 sg13g2_antennanp ANTENNA_1529 (.A(_02936_));
 sg13g2_antennanp ANTENNA_1530 (.A(_02936_));
 sg13g2_antennanp ANTENNA_1531 (.A(_02936_));
 sg13g2_antennanp ANTENNA_1532 (.A(_02936_));
 sg13g2_antennanp ANTENNA_1533 (.A(_03293_));
 sg13g2_antennanp ANTENNA_1534 (.A(_03323_));
 sg13g2_antennanp ANTENNA_1535 (.A(_03324_));
 sg13g2_antennanp ANTENNA_1536 (.A(_03329_));
 sg13g2_antennanp ANTENNA_1537 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1538 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1539 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1540 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1541 (.A(_03697_));
 sg13g2_antennanp ANTENNA_1542 (.A(_03697_));
 sg13g2_antennanp ANTENNA_1543 (.A(_03697_));
 sg13g2_antennanp ANTENNA_1544 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1545 (.A(_05114_));
 sg13g2_antennanp ANTENNA_1546 (.A(_05142_));
 sg13g2_antennanp ANTENNA_1547 (.A(_05173_));
 sg13g2_antennanp ANTENNA_1548 (.A(_05204_));
 sg13g2_antennanp ANTENNA_1549 (.A(_05236_));
 sg13g2_antennanp ANTENNA_1550 (.A(_05248_));
 sg13g2_antennanp ANTENNA_1551 (.A(_05255_));
 sg13g2_antennanp ANTENNA_1552 (.A(_05407_));
 sg13g2_antennanp ANTENNA_1553 (.A(_05412_));
 sg13g2_antennanp ANTENNA_1554 (.A(_05477_));
 sg13g2_antennanp ANTENNA_1555 (.A(_05556_));
 sg13g2_antennanp ANTENNA_1556 (.A(_05681_));
 sg13g2_antennanp ANTENNA_1557 (.A(_05695_));
 sg13g2_antennanp ANTENNA_1558 (.A(_05735_));
 sg13g2_antennanp ANTENNA_1559 (.A(_06655_));
 sg13g2_antennanp ANTENNA_1560 (.A(_06655_));
 sg13g2_antennanp ANTENNA_1561 (.A(_06655_));
 sg13g2_antennanp ANTENNA_1562 (.A(_06655_));
 sg13g2_antennanp ANTENNA_1563 (.A(_07439_));
 sg13g2_antennanp ANTENNA_1564 (.A(_08066_));
 sg13g2_antennanp ANTENNA_1565 (.A(_08066_));
 sg13g2_antennanp ANTENNA_1566 (.A(_08066_));
 sg13g2_antennanp ANTENNA_1567 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1568 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1569 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1570 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1571 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1572 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1573 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1574 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1575 (.A(_08401_));
 sg13g2_antennanp ANTENNA_1576 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1577 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1578 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1579 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1580 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1581 (.A(_08426_));
 sg13g2_antennanp ANTENNA_1582 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1583 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1584 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1585 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1586 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1587 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1588 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1589 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1590 (.A(_08450_));
 sg13g2_antennanp ANTENNA_1591 (.A(_08476_));
 sg13g2_antennanp ANTENNA_1592 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1593 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1594 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1595 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1596 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1597 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1598 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1599 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1600 (.A(_08522_));
 sg13g2_antennanp ANTENNA_1601 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1602 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1603 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1604 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1605 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1606 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1607 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1608 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1609 (.A(_08543_));
 sg13g2_antennanp ANTENNA_1610 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1611 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1612 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1613 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1614 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1615 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1616 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1617 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1618 (.A(_08564_));
 sg13g2_antennanp ANTENNA_1619 (.A(_08583_));
 sg13g2_antennanp ANTENNA_1620 (.A(_08607_));
 sg13g2_antennanp ANTENNA_1621 (.A(_08607_));
 sg13g2_antennanp ANTENNA_1622 (.A(_08607_));
 sg13g2_antennanp ANTENNA_1623 (.A(_08627_));
 sg13g2_antennanp ANTENNA_1624 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1625 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1626 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1627 (.A(_08650_));
 sg13g2_antennanp ANTENNA_1628 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1629 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1630 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1631 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1632 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1633 (.A(_08732_));
 sg13g2_antennanp ANTENNA_1634 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1635 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1636 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1637 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1638 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1639 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1640 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1641 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1642 (.A(_09014_));
 sg13g2_antennanp ANTENNA_1643 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1644 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1645 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1646 (.A(_09040_));
 sg13g2_antennanp ANTENNA_1647 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1648 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1649 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1650 (.A(_09094_));
 sg13g2_antennanp ANTENNA_1651 (.A(_09095_));
 sg13g2_antennanp ANTENNA_1652 (.A(_09095_));
 sg13g2_antennanp ANTENNA_1653 (.A(_09102_));
 sg13g2_antennanp ANTENNA_1654 (.A(_09123_));
 sg13g2_antennanp ANTENNA_1655 (.A(_09123_));
 sg13g2_antennanp ANTENNA_1656 (.A(_09123_));
 sg13g2_antennanp ANTENNA_1657 (.A(_09125_));
 sg13g2_antennanp ANTENNA_1658 (.A(_09125_));
 sg13g2_antennanp ANTENNA_1659 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1660 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1661 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1662 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1663 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1664 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1665 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1666 (.A(_09130_));
 sg13g2_antennanp ANTENNA_1667 (.A(_09246_));
 sg13g2_antennanp ANTENNA_1668 (.A(_09312_));
 sg13g2_antennanp ANTENNA_1669 (.A(_09312_));
 sg13g2_antennanp ANTENNA_1670 (.A(_09315_));
 sg13g2_antennanp ANTENNA_1671 (.A(_09315_));
 sg13g2_antennanp ANTENNA_1672 (.A(_09341_));
 sg13g2_antennanp ANTENNA_1673 (.A(_09443_));
 sg13g2_antennanp ANTENNA_1674 (.A(_09466_));
 sg13g2_antennanp ANTENNA_1675 (.A(_09492_));
 sg13g2_antennanp ANTENNA_1676 (.A(_09514_));
 sg13g2_antennanp ANTENNA_1677 (.A(_09536_));
 sg13g2_antennanp ANTENNA_1678 (.A(_09561_));
 sg13g2_antennanp ANTENNA_1679 (.A(_09585_));
 sg13g2_antennanp ANTENNA_1680 (.A(_09608_));
 sg13g2_antennanp ANTENNA_1681 (.A(_09630_));
 sg13g2_antennanp ANTENNA_1682 (.A(_09759_));
 sg13g2_antennanp ANTENNA_1683 (.A(_09759_));
 sg13g2_antennanp ANTENNA_1684 (.A(_09943_));
 sg13g2_antennanp ANTENNA_1685 (.A(_09943_));
 sg13g2_antennanp ANTENNA_1686 (.A(_09943_));
 sg13g2_antennanp ANTENNA_1687 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1688 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1689 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1690 (.A(_09944_));
 sg13g2_antennanp ANTENNA_1691 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1692 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1693 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1694 (.A(_10187_));
 sg13g2_antennanp ANTENNA_1695 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1696 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1697 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1698 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1699 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1700 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1701 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1702 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1703 (.A(_11761_));
 sg13g2_antennanp ANTENNA_1704 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1705 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1706 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1707 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1708 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1709 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1710 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1711 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1712 (.A(_11795_));
 sg13g2_antennanp ANTENNA_1713 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1714 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1715 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1716 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1717 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1718 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1719 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1720 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1721 (.A(_11812_));
 sg13g2_antennanp ANTENNA_1722 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1723 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1724 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1725 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1726 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1727 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1728 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1729 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1730 (.A(_11832_));
 sg13g2_antennanp ANTENNA_1731 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1732 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1733 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1734 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1735 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1736 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1737 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1738 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1739 (.A(_11925_));
 sg13g2_antennanp ANTENNA_1740 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1741 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1742 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1743 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1744 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1745 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1746 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1747 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1748 (.A(_11945_));
 sg13g2_antennanp ANTENNA_1749 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1750 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1751 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1752 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1753 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1754 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1755 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1756 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1757 (.A(_11974_));
 sg13g2_antennanp ANTENNA_1758 (.A(clk));
 sg13g2_antennanp ANTENNA_1759 (.A(clk));
 sg13g2_antennanp ANTENNA_1760 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1761 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1762 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1763 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1764 (.A(net3));
 sg13g2_antennanp ANTENNA_1765 (.A(net3));
 sg13g2_antennanp ANTENNA_1766 (.A(net3));
 sg13g2_antennanp ANTENNA_1767 (.A(net19));
 sg13g2_antennanp ANTENNA_1768 (.A(net19));
 sg13g2_antennanp ANTENNA_1769 (.A(net366));
 sg13g2_antennanp ANTENNA_1770 (.A(net366));
 sg13g2_antennanp ANTENNA_1771 (.A(net366));
 sg13g2_antennanp ANTENNA_1772 (.A(net366));
 sg13g2_antennanp ANTENNA_1773 (.A(net366));
 sg13g2_antennanp ANTENNA_1774 (.A(net366));
 sg13g2_antennanp ANTENNA_1775 (.A(net366));
 sg13g2_antennanp ANTENNA_1776 (.A(net366));
 sg13g2_antennanp ANTENNA_1777 (.A(net366));
 sg13g2_antennanp ANTENNA_1778 (.A(net366));
 sg13g2_antennanp ANTENNA_1779 (.A(net366));
 sg13g2_antennanp ANTENNA_1780 (.A(net366));
 sg13g2_antennanp ANTENNA_1781 (.A(net468));
 sg13g2_antennanp ANTENNA_1782 (.A(net468));
 sg13g2_antennanp ANTENNA_1783 (.A(net468));
 sg13g2_antennanp ANTENNA_1784 (.A(net468));
 sg13g2_antennanp ANTENNA_1785 (.A(net468));
 sg13g2_antennanp ANTENNA_1786 (.A(net468));
 sg13g2_antennanp ANTENNA_1787 (.A(net468));
 sg13g2_antennanp ANTENNA_1788 (.A(net468));
 sg13g2_antennanp ANTENNA_1789 (.A(net468));
 sg13g2_antennanp ANTENNA_1790 (.A(net551));
 sg13g2_antennanp ANTENNA_1791 (.A(net551));
 sg13g2_antennanp ANTENNA_1792 (.A(net551));
 sg13g2_antennanp ANTENNA_1793 (.A(net551));
 sg13g2_antennanp ANTENNA_1794 (.A(net551));
 sg13g2_antennanp ANTENNA_1795 (.A(net551));
 sg13g2_antennanp ANTENNA_1796 (.A(net551));
 sg13g2_antennanp ANTENNA_1797 (.A(net551));
 sg13g2_antennanp ANTENNA_1798 (.A(net551));
 sg13g2_antennanp ANTENNA_1799 (.A(net594));
 sg13g2_antennanp ANTENNA_1800 (.A(net594));
 sg13g2_antennanp ANTENNA_1801 (.A(net594));
 sg13g2_antennanp ANTENNA_1802 (.A(net594));
 sg13g2_antennanp ANTENNA_1803 (.A(net594));
 sg13g2_antennanp ANTENNA_1804 (.A(net594));
 sg13g2_antennanp ANTENNA_1805 (.A(net594));
 sg13g2_antennanp ANTENNA_1806 (.A(net594));
 sg13g2_antennanp ANTENNA_1807 (.A(net643));
 sg13g2_antennanp ANTENNA_1808 (.A(net643));
 sg13g2_antennanp ANTENNA_1809 (.A(net643));
 sg13g2_antennanp ANTENNA_1810 (.A(net643));
 sg13g2_antennanp ANTENNA_1811 (.A(net643));
 sg13g2_antennanp ANTENNA_1812 (.A(net643));
 sg13g2_antennanp ANTENNA_1813 (.A(net643));
 sg13g2_antennanp ANTENNA_1814 (.A(net643));
 sg13g2_antennanp ANTENNA_1815 (.A(net643));
 sg13g2_antennanp ANTENNA_1816 (.A(net643));
 sg13g2_antennanp ANTENNA_1817 (.A(net643));
 sg13g2_antennanp ANTENNA_1818 (.A(net643));
 sg13g2_antennanp ANTENNA_1819 (.A(net643));
 sg13g2_antennanp ANTENNA_1820 (.A(net643));
 sg13g2_antennanp ANTENNA_1821 (.A(net643));
 sg13g2_antennanp ANTENNA_1822 (.A(net643));
 sg13g2_antennanp ANTENNA_1823 (.A(net643));
 sg13g2_antennanp ANTENNA_1824 (.A(net643));
 sg13g2_antennanp ANTENNA_1825 (.A(net643));
 sg13g2_antennanp ANTENNA_1826 (.A(net643));
 sg13g2_antennanp ANTENNA_1827 (.A(net643));
 sg13g2_antennanp ANTENNA_1828 (.A(net643));
 sg13g2_antennanp ANTENNA_1829 (.A(net643));
 sg13g2_antennanp ANTENNA_1830 (.A(net643));
 sg13g2_antennanp ANTENNA_1831 (.A(net643));
 sg13g2_antennanp ANTENNA_1832 (.A(net643));
 sg13g2_antennanp ANTENNA_1833 (.A(net643));
 sg13g2_antennanp ANTENNA_1834 (.A(net643));
 sg13g2_antennanp ANTENNA_1835 (.A(net643));
 sg13g2_antennanp ANTENNA_1836 (.A(net643));
 sg13g2_antennanp ANTENNA_1837 (.A(net643));
 sg13g2_antennanp ANTENNA_1838 (.A(net643));
 sg13g2_antennanp ANTENNA_1839 (.A(net643));
 sg13g2_antennanp ANTENNA_1840 (.A(net643));
 sg13g2_antennanp ANTENNA_1841 (.A(net643));
 sg13g2_antennanp ANTENNA_1842 (.A(net643));
 sg13g2_antennanp ANTENNA_1843 (.A(net643));
 sg13g2_antennanp ANTENNA_1844 (.A(net643));
 sg13g2_antennanp ANTENNA_1845 (.A(net667));
 sg13g2_antennanp ANTENNA_1846 (.A(net667));
 sg13g2_antennanp ANTENNA_1847 (.A(net667));
 sg13g2_antennanp ANTENNA_1848 (.A(net667));
 sg13g2_antennanp ANTENNA_1849 (.A(net667));
 sg13g2_antennanp ANTENNA_1850 (.A(net667));
 sg13g2_antennanp ANTENNA_1851 (.A(net667));
 sg13g2_antennanp ANTENNA_1852 (.A(net667));
 sg13g2_antennanp ANTENNA_1853 (.A(net667));
 sg13g2_antennanp ANTENNA_1854 (.A(net667));
 sg13g2_antennanp ANTENNA_1855 (.A(net667));
 sg13g2_antennanp ANTENNA_1856 (.A(net667));
 sg13g2_antennanp ANTENNA_1857 (.A(net667));
 sg13g2_antennanp ANTENNA_1858 (.A(net667));
 sg13g2_antennanp ANTENNA_1859 (.A(net667));
 sg13g2_antennanp ANTENNA_1860 (.A(net679));
 sg13g2_antennanp ANTENNA_1861 (.A(net679));
 sg13g2_antennanp ANTENNA_1862 (.A(net679));
 sg13g2_antennanp ANTENNA_1863 (.A(net679));
 sg13g2_antennanp ANTENNA_1864 (.A(net679));
 sg13g2_antennanp ANTENNA_1865 (.A(net679));
 sg13g2_antennanp ANTENNA_1866 (.A(net679));
 sg13g2_antennanp ANTENNA_1867 (.A(net679));
 sg13g2_antennanp ANTENNA_1868 (.A(net679));
 sg13g2_antennanp ANTENNA_1869 (.A(net679));
 sg13g2_antennanp ANTENNA_1870 (.A(net679));
 sg13g2_antennanp ANTENNA_1871 (.A(net679));
 sg13g2_antennanp ANTENNA_1872 (.A(net679));
 sg13g2_antennanp ANTENNA_1873 (.A(net679));
 sg13g2_antennanp ANTENNA_1874 (.A(net679));
 sg13g2_antennanp ANTENNA_1875 (.A(net780));
 sg13g2_antennanp ANTENNA_1876 (.A(net780));
 sg13g2_antennanp ANTENNA_1877 (.A(net780));
 sg13g2_antennanp ANTENNA_1878 (.A(net780));
 sg13g2_antennanp ANTENNA_1879 (.A(net780));
 sg13g2_antennanp ANTENNA_1880 (.A(net780));
 sg13g2_antennanp ANTENNA_1881 (.A(net780));
 sg13g2_antennanp ANTENNA_1882 (.A(net780));
 sg13g2_antennanp ANTENNA_1883 (.A(net780));
 sg13g2_antennanp ANTENNA_1884 (.A(net848));
 sg13g2_antennanp ANTENNA_1885 (.A(net848));
 sg13g2_antennanp ANTENNA_1886 (.A(net848));
 sg13g2_antennanp ANTENNA_1887 (.A(net848));
 sg13g2_antennanp ANTENNA_1888 (.A(net848));
 sg13g2_antennanp ANTENNA_1889 (.A(net848));
 sg13g2_antennanp ANTENNA_1890 (.A(net848));
 sg13g2_antennanp ANTENNA_1891 (.A(net848));
 sg13g2_antennanp ANTENNA_1892 (.A(net848));
 sg13g2_antennanp ANTENNA_1893 (.A(net848));
 sg13g2_antennanp ANTENNA_1894 (.A(net848));
 sg13g2_antennanp ANTENNA_1895 (.A(net848));
 sg13g2_antennanp ANTENNA_1896 (.A(net848));
 sg13g2_antennanp ANTENNA_1897 (.A(net848));
 sg13g2_antennanp ANTENNA_1898 (.A(net848));
 sg13g2_antennanp ANTENNA_1899 (.A(net848));
 sg13g2_antennanp ANTENNA_1900 (.A(net853));
 sg13g2_antennanp ANTENNA_1901 (.A(net853));
 sg13g2_antennanp ANTENNA_1902 (.A(net853));
 sg13g2_antennanp ANTENNA_1903 (.A(net853));
 sg13g2_antennanp ANTENNA_1904 (.A(net853));
 sg13g2_antennanp ANTENNA_1905 (.A(net853));
 sg13g2_antennanp ANTENNA_1906 (.A(net853));
 sg13g2_antennanp ANTENNA_1907 (.A(net853));
 sg13g2_antennanp ANTENNA_1908 (.A(net853));
 sg13g2_antennanp ANTENNA_1909 (.A(net853));
 sg13g2_antennanp ANTENNA_1910 (.A(net853));
 sg13g2_antennanp ANTENNA_1911 (.A(net853));
 sg13g2_antennanp ANTENNA_1912 (.A(net853));
 sg13g2_antennanp ANTENNA_1913 (.A(net853));
 sg13g2_antennanp ANTENNA_1914 (.A(net853));
 sg13g2_antennanp ANTENNA_1915 (.A(net853));
 sg13g2_antennanp ANTENNA_1916 (.A(net853));
 sg13g2_antennanp ANTENNA_1917 (.A(net853));
 sg13g2_antennanp ANTENNA_1918 (.A(net853));
 sg13g2_antennanp ANTENNA_1919 (.A(net853));
 sg13g2_antennanp ANTENNA_1920 (.A(net853));
 sg13g2_antennanp ANTENNA_1921 (.A(net853));
 sg13g2_antennanp ANTENNA_1922 (.A(net894));
 sg13g2_antennanp ANTENNA_1923 (.A(net894));
 sg13g2_antennanp ANTENNA_1924 (.A(net894));
 sg13g2_antennanp ANTENNA_1925 (.A(net894));
 sg13g2_antennanp ANTENNA_1926 (.A(net894));
 sg13g2_antennanp ANTENNA_1927 (.A(net894));
 sg13g2_antennanp ANTENNA_1928 (.A(net894));
 sg13g2_antennanp ANTENNA_1929 (.A(net894));
 sg13g2_antennanp ANTENNA_1930 (.A(net894));
 sg13g2_antennanp ANTENNA_1931 (.A(net952));
 sg13g2_antennanp ANTENNA_1932 (.A(net952));
 sg13g2_antennanp ANTENNA_1933 (.A(net952));
 sg13g2_antennanp ANTENNA_1934 (.A(net952));
 sg13g2_antennanp ANTENNA_1935 (.A(net952));
 sg13g2_antennanp ANTENNA_1936 (.A(net952));
 sg13g2_antennanp ANTENNA_1937 (.A(net952));
 sg13g2_antennanp ANTENNA_1938 (.A(net952));
 sg13g2_antennanp ANTENNA_1939 (.A(net952));
 sg13g2_antennanp ANTENNA_1940 (.A(net952));
 sg13g2_antennanp ANTENNA_1941 (.A(net952));
 sg13g2_antennanp ANTENNA_1942 (.A(net952));
 sg13g2_antennanp ANTENNA_1943 (.A(net952));
 sg13g2_antennanp ANTENNA_1944 (.A(net952));
 sg13g2_antennanp ANTENNA_1945 (.A(net952));
 sg13g2_antennanp ANTENNA_1946 (.A(net952));
 sg13g2_antennanp ANTENNA_1947 (.A(net952));
 sg13g2_antennanp ANTENNA_1948 (.A(net952));
 sg13g2_antennanp ANTENNA_1949 (.A(net952));
 sg13g2_antennanp ANTENNA_1950 (.A(net952));
 sg13g2_antennanp ANTENNA_1951 (.A(net956));
 sg13g2_antennanp ANTENNA_1952 (.A(net956));
 sg13g2_antennanp ANTENNA_1953 (.A(net956));
 sg13g2_antennanp ANTENNA_1954 (.A(net956));
 sg13g2_antennanp ANTENNA_1955 (.A(net956));
 sg13g2_antennanp ANTENNA_1956 (.A(net956));
 sg13g2_antennanp ANTENNA_1957 (.A(net956));
 sg13g2_antennanp ANTENNA_1958 (.A(net956));
 sg13g2_antennanp ANTENNA_1959 (.A(net956));
 sg13g2_antennanp ANTENNA_1960 (.A(net958));
 sg13g2_antennanp ANTENNA_1961 (.A(net958));
 sg13g2_antennanp ANTENNA_1962 (.A(net958));
 sg13g2_antennanp ANTENNA_1963 (.A(net958));
 sg13g2_antennanp ANTENNA_1964 (.A(net958));
 sg13g2_antennanp ANTENNA_1965 (.A(net958));
 sg13g2_antennanp ANTENNA_1966 (.A(net958));
 sg13g2_antennanp ANTENNA_1967 (.A(net958));
 sg13g2_antennanp ANTENNA_1968 (.A(net986));
 sg13g2_antennanp ANTENNA_1969 (.A(net986));
 sg13g2_antennanp ANTENNA_1970 (.A(net986));
 sg13g2_antennanp ANTENNA_1971 (.A(net986));
 sg13g2_antennanp ANTENNA_1972 (.A(net986));
 sg13g2_antennanp ANTENNA_1973 (.A(net986));
 sg13g2_antennanp ANTENNA_1974 (.A(net986));
 sg13g2_antennanp ANTENNA_1975 (.A(net986));
 sg13g2_antennanp ANTENNA_1976 (.A(net986));
 sg13g2_antennanp ANTENNA_1977 (.A(net986));
 sg13g2_antennanp ANTENNA_1978 (.A(net986));
 sg13g2_antennanp ANTENNA_1979 (.A(net986));
 sg13g2_antennanp ANTENNA_1980 (.A(net986));
 sg13g2_antennanp ANTENNA_1981 (.A(net986));
 sg13g2_antennanp ANTENNA_1982 (.A(net986));
 sg13g2_antennanp ANTENNA_1983 (.A(net986));
 sg13g2_antennanp ANTENNA_1984 (.A(net991));
 sg13g2_antennanp ANTENNA_1985 (.A(net991));
 sg13g2_antennanp ANTENNA_1986 (.A(net991));
 sg13g2_antennanp ANTENNA_1987 (.A(net991));
 sg13g2_antennanp ANTENNA_1988 (.A(net991));
 sg13g2_antennanp ANTENNA_1989 (.A(net991));
 sg13g2_antennanp ANTENNA_1990 (.A(net991));
 sg13g2_antennanp ANTENNA_1991 (.A(net991));
 sg13g2_antennanp ANTENNA_1992 (.A(net991));
 sg13g2_antennanp ANTENNA_1993 (.A(_00237_));
 sg13g2_antennanp ANTENNA_1994 (.A(_00789_));
 sg13g2_antennanp ANTENNA_1995 (.A(_00798_));
 sg13g2_antennanp ANTENNA_1996 (.A(_00930_));
 sg13g2_antennanp ANTENNA_1997 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1998 (.A(_02788_));
 sg13g2_antennanp ANTENNA_1999 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2000 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2001 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2002 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2003 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2004 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2005 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2006 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2007 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2008 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2009 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2010 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2011 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2012 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2013 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2014 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2015 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2016 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2017 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2018 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2019 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2020 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2021 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2022 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2023 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2024 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2025 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2026 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2027 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2028 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2029 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2030 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2031 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2032 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2033 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2034 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2035 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2036 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2037 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2038 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2039 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2040 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2041 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2042 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2043 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2044 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2045 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2046 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2047 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2048 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2049 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2050 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2051 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2052 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2053 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2054 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2055 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2056 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2057 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2058 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2059 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2060 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2061 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2062 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2063 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2064 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2065 (.A(_03293_));
 sg13g2_antennanp ANTENNA_2066 (.A(_03317_));
 sg13g2_antennanp ANTENNA_2067 (.A(_03317_));
 sg13g2_antennanp ANTENNA_2068 (.A(_03323_));
 sg13g2_antennanp ANTENNA_2069 (.A(_03324_));
 sg13g2_antennanp ANTENNA_2070 (.A(_03329_));
 sg13g2_antennanp ANTENNA_2071 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2072 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2073 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2074 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2075 (.A(_03697_));
 sg13g2_antennanp ANTENNA_2076 (.A(_03697_));
 sg13g2_antennanp ANTENNA_2077 (.A(_03697_));
 sg13g2_antennanp ANTENNA_2078 (.A(_03697_));
 sg13g2_antennanp ANTENNA_2079 (.A(_03697_));
 sg13g2_antennanp ANTENNA_2080 (.A(_03697_));
 sg13g2_antennanp ANTENNA_2081 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2082 (.A(_05114_));
 sg13g2_antennanp ANTENNA_2083 (.A(_05142_));
 sg13g2_antennanp ANTENNA_2084 (.A(_05173_));
 sg13g2_antennanp ANTENNA_2085 (.A(_05204_));
 sg13g2_antennanp ANTENNA_2086 (.A(_05236_));
 sg13g2_antennanp ANTENNA_2087 (.A(_05248_));
 sg13g2_antennanp ANTENNA_2088 (.A(_05255_));
 sg13g2_antennanp ANTENNA_2089 (.A(_05407_));
 sg13g2_antennanp ANTENNA_2090 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2091 (.A(_05477_));
 sg13g2_antennanp ANTENNA_2092 (.A(_05556_));
 sg13g2_antennanp ANTENNA_2093 (.A(_05681_));
 sg13g2_antennanp ANTENNA_2094 (.A(_05695_));
 sg13g2_antennanp ANTENNA_2095 (.A(_05708_));
 sg13g2_antennanp ANTENNA_2096 (.A(_05735_));
 sg13g2_antennanp ANTENNA_2097 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2098 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2099 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2100 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2101 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2102 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2103 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2104 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2105 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2106 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2107 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2108 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2109 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2110 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2111 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2112 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2113 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2114 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2115 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2116 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2117 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2118 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2119 (.A(_08426_));
 sg13g2_antennanp ANTENNA_2120 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2121 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2122 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2123 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2124 (.A(_08476_));
 sg13g2_antennanp ANTENNA_2125 (.A(_08498_));
 sg13g2_antennanp ANTENNA_2126 (.A(_08498_));
 sg13g2_antennanp ANTENNA_2127 (.A(_08498_));
 sg13g2_antennanp ANTENNA_2128 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2129 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2130 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2131 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2132 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2133 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2134 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2135 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2136 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2137 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2138 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2139 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2140 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2141 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2142 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2143 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2144 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2145 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2146 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2147 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2148 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2149 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2150 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2151 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2152 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2153 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2154 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2155 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2156 (.A(_08583_));
 sg13g2_antennanp ANTENNA_2157 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2158 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2159 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2160 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2161 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2162 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2163 (.A(_08627_));
 sg13g2_antennanp ANTENNA_2164 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2165 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2166 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2167 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2168 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2169 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2170 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2171 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2172 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2173 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2174 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2175 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2176 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2177 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2178 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2179 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2180 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2181 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2182 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2183 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2184 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2185 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2186 (.A(_09102_));
 sg13g2_antennanp ANTENNA_2187 (.A(_09123_));
 sg13g2_antennanp ANTENNA_2188 (.A(_09123_));
 sg13g2_antennanp ANTENNA_2189 (.A(_09123_));
 sg13g2_antennanp ANTENNA_2190 (.A(_09125_));
 sg13g2_antennanp ANTENNA_2191 (.A(_09125_));
 sg13g2_antennanp ANTENNA_2192 (.A(_09246_));
 sg13g2_antennanp ANTENNA_2193 (.A(_09248_));
 sg13g2_antennanp ANTENNA_2194 (.A(_09312_));
 sg13g2_antennanp ANTENNA_2195 (.A(_09315_));
 sg13g2_antennanp ANTENNA_2196 (.A(_09341_));
 sg13g2_antennanp ANTENNA_2197 (.A(_09443_));
 sg13g2_antennanp ANTENNA_2198 (.A(_09466_));
 sg13g2_antennanp ANTENNA_2199 (.A(_09492_));
 sg13g2_antennanp ANTENNA_2200 (.A(_09514_));
 sg13g2_antennanp ANTENNA_2201 (.A(_09536_));
 sg13g2_antennanp ANTENNA_2202 (.A(_09561_));
 sg13g2_antennanp ANTENNA_2203 (.A(_09585_));
 sg13g2_antennanp ANTENNA_2204 (.A(_09608_));
 sg13g2_antennanp ANTENNA_2205 (.A(_09630_));
 sg13g2_antennanp ANTENNA_2206 (.A(_09759_));
 sg13g2_antennanp ANTENNA_2207 (.A(_09759_));
 sg13g2_antennanp ANTENNA_2208 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2209 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2210 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2211 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2212 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2213 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2214 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2215 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2216 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2217 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2218 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2219 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2220 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2221 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2222 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2223 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2224 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2225 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2226 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2227 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2228 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2229 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2230 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2231 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2232 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2233 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2234 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2235 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2236 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2237 (.A(_11807_));
 sg13g2_antennanp ANTENNA_2238 (.A(_11807_));
 sg13g2_antennanp ANTENNA_2239 (.A(_11807_));
 sg13g2_antennanp ANTENNA_2240 (.A(_11807_));
 sg13g2_antennanp ANTENNA_2241 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2242 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2243 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2244 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2245 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2246 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2247 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2248 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2249 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2250 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2251 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2252 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2253 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2254 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2255 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2256 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2257 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2258 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2259 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2260 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2261 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2262 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2263 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2264 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2265 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2266 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2267 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2268 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2269 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2270 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2271 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2272 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2273 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2274 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2275 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2276 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2277 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2278 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2279 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2280 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2281 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2282 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2283 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2284 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2285 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2286 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2287 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2288 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2289 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2290 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2291 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2292 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2293 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2294 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2295 (.A(clk));
 sg13g2_antennanp ANTENNA_2296 (.A(clk));
 sg13g2_antennanp ANTENNA_2297 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2298 (.A(net3));
 sg13g2_antennanp ANTENNA_2299 (.A(net3));
 sg13g2_antennanp ANTENNA_2300 (.A(net3));
 sg13g2_antennanp ANTENNA_2301 (.A(net19));
 sg13g2_antennanp ANTENNA_2302 (.A(net19));
 sg13g2_antennanp ANTENNA_2303 (.A(net151));
 sg13g2_antennanp ANTENNA_2304 (.A(net151));
 sg13g2_antennanp ANTENNA_2305 (.A(net151));
 sg13g2_antennanp ANTENNA_2306 (.A(net151));
 sg13g2_antennanp ANTENNA_2307 (.A(net151));
 sg13g2_antennanp ANTENNA_2308 (.A(net151));
 sg13g2_antennanp ANTENNA_2309 (.A(net151));
 sg13g2_antennanp ANTENNA_2310 (.A(net151));
 sg13g2_antennanp ANTENNA_2311 (.A(net151));
 sg13g2_antennanp ANTENNA_2312 (.A(net366));
 sg13g2_antennanp ANTENNA_2313 (.A(net366));
 sg13g2_antennanp ANTENNA_2314 (.A(net366));
 sg13g2_antennanp ANTENNA_2315 (.A(net366));
 sg13g2_antennanp ANTENNA_2316 (.A(net366));
 sg13g2_antennanp ANTENNA_2317 (.A(net366));
 sg13g2_antennanp ANTENNA_2318 (.A(net366));
 sg13g2_antennanp ANTENNA_2319 (.A(net366));
 sg13g2_antennanp ANTENNA_2320 (.A(net366));
 sg13g2_antennanp ANTENNA_2321 (.A(net366));
 sg13g2_antennanp ANTENNA_2322 (.A(net366));
 sg13g2_antennanp ANTENNA_2323 (.A(net366));
 sg13g2_antennanp ANTENNA_2324 (.A(net366));
 sg13g2_antennanp ANTENNA_2325 (.A(net366));
 sg13g2_antennanp ANTENNA_2326 (.A(net366));
 sg13g2_antennanp ANTENNA_2327 (.A(net366));
 sg13g2_antennanp ANTENNA_2328 (.A(net366));
 sg13g2_antennanp ANTENNA_2329 (.A(net366));
 sg13g2_antennanp ANTENNA_2330 (.A(net366));
 sg13g2_antennanp ANTENNA_2331 (.A(net366));
 sg13g2_antennanp ANTENNA_2332 (.A(net366));
 sg13g2_antennanp ANTENNA_2333 (.A(net468));
 sg13g2_antennanp ANTENNA_2334 (.A(net468));
 sg13g2_antennanp ANTENNA_2335 (.A(net468));
 sg13g2_antennanp ANTENNA_2336 (.A(net468));
 sg13g2_antennanp ANTENNA_2337 (.A(net468));
 sg13g2_antennanp ANTENNA_2338 (.A(net468));
 sg13g2_antennanp ANTENNA_2339 (.A(net468));
 sg13g2_antennanp ANTENNA_2340 (.A(net468));
 sg13g2_antennanp ANTENNA_2341 (.A(net468));
 sg13g2_antennanp ANTENNA_2342 (.A(net524));
 sg13g2_antennanp ANTENNA_2343 (.A(net524));
 sg13g2_antennanp ANTENNA_2344 (.A(net524));
 sg13g2_antennanp ANTENNA_2345 (.A(net524));
 sg13g2_antennanp ANTENNA_2346 (.A(net524));
 sg13g2_antennanp ANTENNA_2347 (.A(net524));
 sg13g2_antennanp ANTENNA_2348 (.A(net524));
 sg13g2_antennanp ANTENNA_2349 (.A(net524));
 sg13g2_antennanp ANTENNA_2350 (.A(net551));
 sg13g2_antennanp ANTENNA_2351 (.A(net551));
 sg13g2_antennanp ANTENNA_2352 (.A(net551));
 sg13g2_antennanp ANTENNA_2353 (.A(net551));
 sg13g2_antennanp ANTENNA_2354 (.A(net551));
 sg13g2_antennanp ANTENNA_2355 (.A(net551));
 sg13g2_antennanp ANTENNA_2356 (.A(net551));
 sg13g2_antennanp ANTENNA_2357 (.A(net551));
 sg13g2_antennanp ANTENNA_2358 (.A(net551));
 sg13g2_antennanp ANTENNA_2359 (.A(net594));
 sg13g2_antennanp ANTENNA_2360 (.A(net594));
 sg13g2_antennanp ANTENNA_2361 (.A(net594));
 sg13g2_antennanp ANTENNA_2362 (.A(net594));
 sg13g2_antennanp ANTENNA_2363 (.A(net594));
 sg13g2_antennanp ANTENNA_2364 (.A(net594));
 sg13g2_antennanp ANTENNA_2365 (.A(net594));
 sg13g2_antennanp ANTENNA_2366 (.A(net594));
 sg13g2_antennanp ANTENNA_2367 (.A(net638));
 sg13g2_antennanp ANTENNA_2368 (.A(net638));
 sg13g2_antennanp ANTENNA_2369 (.A(net638));
 sg13g2_antennanp ANTENNA_2370 (.A(net638));
 sg13g2_antennanp ANTENNA_2371 (.A(net638));
 sg13g2_antennanp ANTENNA_2372 (.A(net638));
 sg13g2_antennanp ANTENNA_2373 (.A(net638));
 sg13g2_antennanp ANTENNA_2374 (.A(net638));
 sg13g2_antennanp ANTENNA_2375 (.A(net638));
 sg13g2_antennanp ANTENNA_2376 (.A(net638));
 sg13g2_antennanp ANTENNA_2377 (.A(net638));
 sg13g2_antennanp ANTENNA_2378 (.A(net638));
 sg13g2_antennanp ANTENNA_2379 (.A(net638));
 sg13g2_antennanp ANTENNA_2380 (.A(net643));
 sg13g2_antennanp ANTENNA_2381 (.A(net643));
 sg13g2_antennanp ANTENNA_2382 (.A(net643));
 sg13g2_antennanp ANTENNA_2383 (.A(net643));
 sg13g2_antennanp ANTENNA_2384 (.A(net643));
 sg13g2_antennanp ANTENNA_2385 (.A(net643));
 sg13g2_antennanp ANTENNA_2386 (.A(net643));
 sg13g2_antennanp ANTENNA_2387 (.A(net643));
 sg13g2_antennanp ANTENNA_2388 (.A(net643));
 sg13g2_antennanp ANTENNA_2389 (.A(net643));
 sg13g2_antennanp ANTENNA_2390 (.A(net643));
 sg13g2_antennanp ANTENNA_2391 (.A(net643));
 sg13g2_antennanp ANTENNA_2392 (.A(net643));
 sg13g2_antennanp ANTENNA_2393 (.A(net643));
 sg13g2_antennanp ANTENNA_2394 (.A(net643));
 sg13g2_antennanp ANTENNA_2395 (.A(net643));
 sg13g2_antennanp ANTENNA_2396 (.A(net643));
 sg13g2_antennanp ANTENNA_2397 (.A(net643));
 sg13g2_antennanp ANTENNA_2398 (.A(net643));
 sg13g2_antennanp ANTENNA_2399 (.A(net643));
 sg13g2_antennanp ANTENNA_2400 (.A(net643));
 sg13g2_antennanp ANTENNA_2401 (.A(net643));
 sg13g2_antennanp ANTENNA_2402 (.A(net643));
 sg13g2_antennanp ANTENNA_2403 (.A(net643));
 sg13g2_antennanp ANTENNA_2404 (.A(net643));
 sg13g2_antennanp ANTENNA_2405 (.A(net667));
 sg13g2_antennanp ANTENNA_2406 (.A(net667));
 sg13g2_antennanp ANTENNA_2407 (.A(net667));
 sg13g2_antennanp ANTENNA_2408 (.A(net667));
 sg13g2_antennanp ANTENNA_2409 (.A(net667));
 sg13g2_antennanp ANTENNA_2410 (.A(net667));
 sg13g2_antennanp ANTENNA_2411 (.A(net667));
 sg13g2_antennanp ANTENNA_2412 (.A(net667));
 sg13g2_antennanp ANTENNA_2413 (.A(net667));
 sg13g2_antennanp ANTENNA_2414 (.A(net667));
 sg13g2_antennanp ANTENNA_2415 (.A(net667));
 sg13g2_antennanp ANTENNA_2416 (.A(net667));
 sg13g2_antennanp ANTENNA_2417 (.A(net667));
 sg13g2_antennanp ANTENNA_2418 (.A(net667));
 sg13g2_antennanp ANTENNA_2419 (.A(net667));
 sg13g2_antennanp ANTENNA_2420 (.A(net667));
 sg13g2_antennanp ANTENNA_2421 (.A(net667));
 sg13g2_antennanp ANTENNA_2422 (.A(net679));
 sg13g2_antennanp ANTENNA_2423 (.A(net679));
 sg13g2_antennanp ANTENNA_2424 (.A(net679));
 sg13g2_antennanp ANTENNA_2425 (.A(net679));
 sg13g2_antennanp ANTENNA_2426 (.A(net679));
 sg13g2_antennanp ANTENNA_2427 (.A(net679));
 sg13g2_antennanp ANTENNA_2428 (.A(net679));
 sg13g2_antennanp ANTENNA_2429 (.A(net679));
 sg13g2_antennanp ANTENNA_2430 (.A(net679));
 sg13g2_antennanp ANTENNA_2431 (.A(net848));
 sg13g2_antennanp ANTENNA_2432 (.A(net848));
 sg13g2_antennanp ANTENNA_2433 (.A(net848));
 sg13g2_antennanp ANTENNA_2434 (.A(net848));
 sg13g2_antennanp ANTENNA_2435 (.A(net848));
 sg13g2_antennanp ANTENNA_2436 (.A(net848));
 sg13g2_antennanp ANTENNA_2437 (.A(net848));
 sg13g2_antennanp ANTENNA_2438 (.A(net848));
 sg13g2_antennanp ANTENNA_2439 (.A(net848));
 sg13g2_antennanp ANTENNA_2440 (.A(net851));
 sg13g2_antennanp ANTENNA_2441 (.A(net851));
 sg13g2_antennanp ANTENNA_2442 (.A(net851));
 sg13g2_antennanp ANTENNA_2443 (.A(net851));
 sg13g2_antennanp ANTENNA_2444 (.A(net851));
 sg13g2_antennanp ANTENNA_2445 (.A(net851));
 sg13g2_antennanp ANTENNA_2446 (.A(net851));
 sg13g2_antennanp ANTENNA_2447 (.A(net851));
 sg13g2_antennanp ANTENNA_2448 (.A(net853));
 sg13g2_antennanp ANTENNA_2449 (.A(net853));
 sg13g2_antennanp ANTENNA_2450 (.A(net853));
 sg13g2_antennanp ANTENNA_2451 (.A(net853));
 sg13g2_antennanp ANTENNA_2452 (.A(net853));
 sg13g2_antennanp ANTENNA_2453 (.A(net853));
 sg13g2_antennanp ANTENNA_2454 (.A(net853));
 sg13g2_antennanp ANTENNA_2455 (.A(net853));
 sg13g2_antennanp ANTENNA_2456 (.A(net853));
 sg13g2_antennanp ANTENNA_2457 (.A(net853));
 sg13g2_antennanp ANTENNA_2458 (.A(net853));
 sg13g2_antennanp ANTENNA_2459 (.A(net853));
 sg13g2_antennanp ANTENNA_2460 (.A(net853));
 sg13g2_antennanp ANTENNA_2461 (.A(net853));
 sg13g2_antennanp ANTENNA_2462 (.A(net853));
 sg13g2_antennanp ANTENNA_2463 (.A(net853));
 sg13g2_antennanp ANTENNA_2464 (.A(net853));
 sg13g2_antennanp ANTENNA_2465 (.A(net853));
 sg13g2_antennanp ANTENNA_2466 (.A(net853));
 sg13g2_antennanp ANTENNA_2467 (.A(net853));
 sg13g2_antennanp ANTENNA_2468 (.A(net853));
 sg13g2_antennanp ANTENNA_2469 (.A(net853));
 sg13g2_antennanp ANTENNA_2470 (.A(net956));
 sg13g2_antennanp ANTENNA_2471 (.A(net956));
 sg13g2_antennanp ANTENNA_2472 (.A(net956));
 sg13g2_antennanp ANTENNA_2473 (.A(net956));
 sg13g2_antennanp ANTENNA_2474 (.A(net956));
 sg13g2_antennanp ANTENNA_2475 (.A(net956));
 sg13g2_antennanp ANTENNA_2476 (.A(net956));
 sg13g2_antennanp ANTENNA_2477 (.A(net956));
 sg13g2_antennanp ANTENNA_2478 (.A(net956));
 sg13g2_antennanp ANTENNA_2479 (.A(net958));
 sg13g2_antennanp ANTENNA_2480 (.A(net958));
 sg13g2_antennanp ANTENNA_2481 (.A(net958));
 sg13g2_antennanp ANTENNA_2482 (.A(net958));
 sg13g2_antennanp ANTENNA_2483 (.A(net958));
 sg13g2_antennanp ANTENNA_2484 (.A(net958));
 sg13g2_antennanp ANTENNA_2485 (.A(net958));
 sg13g2_antennanp ANTENNA_2486 (.A(net958));
 sg13g2_antennanp ANTENNA_2487 (.A(net958));
 sg13g2_antennanp ANTENNA_2488 (.A(net986));
 sg13g2_antennanp ANTENNA_2489 (.A(net986));
 sg13g2_antennanp ANTENNA_2490 (.A(net986));
 sg13g2_antennanp ANTENNA_2491 (.A(net986));
 sg13g2_antennanp ANTENNA_2492 (.A(net986));
 sg13g2_antennanp ANTENNA_2493 (.A(net986));
 sg13g2_antennanp ANTENNA_2494 (.A(net986));
 sg13g2_antennanp ANTENNA_2495 (.A(net986));
 sg13g2_antennanp ANTENNA_2496 (.A(net986));
 sg13g2_antennanp ANTENNA_2497 (.A(net986));
 sg13g2_antennanp ANTENNA_2498 (.A(net986));
 sg13g2_antennanp ANTENNA_2499 (.A(net986));
 sg13g2_antennanp ANTENNA_2500 (.A(net986));
 sg13g2_antennanp ANTENNA_2501 (.A(net986));
 sg13g2_antennanp ANTENNA_2502 (.A(net986));
 sg13g2_antennanp ANTENNA_2503 (.A(net986));
 sg13g2_antennanp ANTENNA_2504 (.A(net986));
 sg13g2_antennanp ANTENNA_2505 (.A(net986));
 sg13g2_antennanp ANTENNA_2506 (.A(net991));
 sg13g2_antennanp ANTENNA_2507 (.A(net991));
 sg13g2_antennanp ANTENNA_2508 (.A(net991));
 sg13g2_antennanp ANTENNA_2509 (.A(net991));
 sg13g2_antennanp ANTENNA_2510 (.A(net991));
 sg13g2_antennanp ANTENNA_2511 (.A(net991));
 sg13g2_antennanp ANTENNA_2512 (.A(net991));
 sg13g2_antennanp ANTENNA_2513 (.A(net991));
 sg13g2_antennanp ANTENNA_2514 (.A(net991));
 sg13g2_antennanp ANTENNA_2515 (.A(_00237_));
 sg13g2_antennanp ANTENNA_2516 (.A(_00789_));
 sg13g2_antennanp ANTENNA_2517 (.A(_00798_));
 sg13g2_antennanp ANTENNA_2518 (.A(_00930_));
 sg13g2_antennanp ANTENNA_2519 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2520 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2521 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2522 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2523 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2524 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2525 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2526 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2527 (.A(_02788_));
 sg13g2_antennanp ANTENNA_2528 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2529 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2530 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2531 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2532 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2533 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2534 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2535 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2536 (.A(_02797_));
 sg13g2_antennanp ANTENNA_2537 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2538 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2539 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2540 (.A(_02801_));
 sg13g2_antennanp ANTENNA_2541 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2542 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2543 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2544 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2545 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2546 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2547 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2548 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2549 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2550 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2551 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2552 (.A(_02908_));
 sg13g2_antennanp ANTENNA_2553 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2554 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2555 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2556 (.A(_02917_));
 sg13g2_antennanp ANTENNA_2557 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2558 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2559 (.A(_02918_));
 sg13g2_antennanp ANTENNA_2560 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2561 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2562 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2563 (.A(_02919_));
 sg13g2_antennanp ANTENNA_2564 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2565 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2566 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2567 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2568 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2569 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2570 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2571 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2572 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2573 (.A(_02920_));
 sg13g2_antennanp ANTENNA_2574 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2575 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2576 (.A(_02922_));
 sg13g2_antennanp ANTENNA_2577 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2578 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2579 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2580 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2581 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2582 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2583 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2584 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2585 (.A(_02927_));
 sg13g2_antennanp ANTENNA_2586 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2587 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2588 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2589 (.A(_02936_));
 sg13g2_antennanp ANTENNA_2590 (.A(_03293_));
 sg13g2_antennanp ANTENNA_2591 (.A(_03317_));
 sg13g2_antennanp ANTENNA_2592 (.A(_03317_));
 sg13g2_antennanp ANTENNA_2593 (.A(_03323_));
 sg13g2_antennanp ANTENNA_2594 (.A(_03324_));
 sg13g2_antennanp ANTENNA_2595 (.A(_03329_));
 sg13g2_antennanp ANTENNA_2596 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2597 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2598 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2599 (.A(_03397_));
 sg13g2_antennanp ANTENNA_2600 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2601 (.A(_05114_));
 sg13g2_antennanp ANTENNA_2602 (.A(_05142_));
 sg13g2_antennanp ANTENNA_2603 (.A(_05173_));
 sg13g2_antennanp ANTENNA_2604 (.A(_05204_));
 sg13g2_antennanp ANTENNA_2605 (.A(_05236_));
 sg13g2_antennanp ANTENNA_2606 (.A(_05248_));
 sg13g2_antennanp ANTENNA_2607 (.A(_05255_));
 sg13g2_antennanp ANTENNA_2608 (.A(_05407_));
 sg13g2_antennanp ANTENNA_2609 (.A(_05412_));
 sg13g2_antennanp ANTENNA_2610 (.A(_05477_));
 sg13g2_antennanp ANTENNA_2611 (.A(_05556_));
 sg13g2_antennanp ANTENNA_2612 (.A(_05681_));
 sg13g2_antennanp ANTENNA_2613 (.A(_05695_));
 sg13g2_antennanp ANTENNA_2614 (.A(_05708_));
 sg13g2_antennanp ANTENNA_2615 (.A(_05735_));
 sg13g2_antennanp ANTENNA_2616 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2617 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2618 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2619 (.A(_06655_));
 sg13g2_antennanp ANTENNA_2620 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2621 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2622 (.A(_07476_));
 sg13g2_antennanp ANTENNA_2623 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2624 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2625 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2626 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2627 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2628 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2629 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2630 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2631 (.A(_08401_));
 sg13g2_antennanp ANTENNA_2632 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2633 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2634 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2635 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2636 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2637 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2638 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2639 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2640 (.A(_08450_));
 sg13g2_antennanp ANTENNA_2641 (.A(_08476_));
 sg13g2_antennanp ANTENNA_2642 (.A(_08498_));
 sg13g2_antennanp ANTENNA_2643 (.A(_08498_));
 sg13g2_antennanp ANTENNA_2644 (.A(_08498_));
 sg13g2_antennanp ANTENNA_2645 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2646 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2647 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2648 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2649 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2650 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2651 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2652 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2653 (.A(_08522_));
 sg13g2_antennanp ANTENNA_2654 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2655 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2656 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2657 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2658 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2659 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2660 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2661 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2662 (.A(_08543_));
 sg13g2_antennanp ANTENNA_2663 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2664 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2665 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2666 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2667 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2668 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2669 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2670 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2671 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2672 (.A(_08564_));
 sg13g2_antennanp ANTENNA_2673 (.A(_08583_));
 sg13g2_antennanp ANTENNA_2674 (.A(_08583_));
 sg13g2_antennanp ANTENNA_2675 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2676 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2677 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2678 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2679 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2680 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2681 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2682 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2683 (.A(_08607_));
 sg13g2_antennanp ANTENNA_2684 (.A(_08627_));
 sg13g2_antennanp ANTENNA_2685 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2686 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2687 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2688 (.A(_08650_));
 sg13g2_antennanp ANTENNA_2689 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2690 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2691 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2692 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2693 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2694 (.A(_08732_));
 sg13g2_antennanp ANTENNA_2695 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2696 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2697 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2698 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2699 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2700 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2701 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2702 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2703 (.A(_09014_));
 sg13g2_antennanp ANTENNA_2704 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2705 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2706 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2707 (.A(_09040_));
 sg13g2_antennanp ANTENNA_2708 (.A(_09102_));
 sg13g2_antennanp ANTENNA_2709 (.A(_09119_));
 sg13g2_antennanp ANTENNA_2710 (.A(_09119_));
 sg13g2_antennanp ANTENNA_2711 (.A(_09119_));
 sg13g2_antennanp ANTENNA_2712 (.A(_09123_));
 sg13g2_antennanp ANTENNA_2713 (.A(_09123_));
 sg13g2_antennanp ANTENNA_2714 (.A(_09123_));
 sg13g2_antennanp ANTENNA_2715 (.A(_09125_));
 sg13g2_antennanp ANTENNA_2716 (.A(_09125_));
 sg13g2_antennanp ANTENNA_2717 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2718 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2719 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2720 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2721 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2722 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2723 (.A(_09130_));
 sg13g2_antennanp ANTENNA_2724 (.A(_09248_));
 sg13g2_antennanp ANTENNA_2725 (.A(_09312_));
 sg13g2_antennanp ANTENNA_2726 (.A(_09315_));
 sg13g2_antennanp ANTENNA_2727 (.A(_09341_));
 sg13g2_antennanp ANTENNA_2728 (.A(_09443_));
 sg13g2_antennanp ANTENNA_2729 (.A(_09466_));
 sg13g2_antennanp ANTENNA_2730 (.A(_09492_));
 sg13g2_antennanp ANTENNA_2731 (.A(_09514_));
 sg13g2_antennanp ANTENNA_2732 (.A(_09514_));
 sg13g2_antennanp ANTENNA_2733 (.A(_09536_));
 sg13g2_antennanp ANTENNA_2734 (.A(_09561_));
 sg13g2_antennanp ANTENNA_2735 (.A(_09585_));
 sg13g2_antennanp ANTENNA_2736 (.A(_09608_));
 sg13g2_antennanp ANTENNA_2737 (.A(_09630_));
 sg13g2_antennanp ANTENNA_2738 (.A(_09630_));
 sg13g2_antennanp ANTENNA_2739 (.A(_09759_));
 sg13g2_antennanp ANTENNA_2740 (.A(_09759_));
 sg13g2_antennanp ANTENNA_2741 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2742 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2743 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2744 (.A(_09943_));
 sg13g2_antennanp ANTENNA_2745 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2746 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2747 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2748 (.A(_09944_));
 sg13g2_antennanp ANTENNA_2749 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2750 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2751 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2752 (.A(_10187_));
 sg13g2_antennanp ANTENNA_2753 (.A(_11070_));
 sg13g2_antennanp ANTENNA_2754 (.A(_11070_));
 sg13g2_antennanp ANTENNA_2755 (.A(_11070_));
 sg13g2_antennanp ANTENNA_2756 (.A(_11070_));
 sg13g2_antennanp ANTENNA_2757 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2758 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2759 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2760 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2761 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2762 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2763 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2764 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2765 (.A(_11761_));
 sg13g2_antennanp ANTENNA_2766 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2767 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2768 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2769 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2770 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2771 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2772 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2773 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2774 (.A(_11795_));
 sg13g2_antennanp ANTENNA_2775 (.A(_11807_));
 sg13g2_antennanp ANTENNA_2776 (.A(_11807_));
 sg13g2_antennanp ANTENNA_2777 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2778 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2779 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2780 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2781 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2782 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2783 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2784 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2785 (.A(_11812_));
 sg13g2_antennanp ANTENNA_2786 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2787 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2788 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2789 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2790 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2791 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2792 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2793 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2794 (.A(_11832_));
 sg13g2_antennanp ANTENNA_2795 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2796 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2797 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2798 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2799 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2800 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2801 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2802 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2803 (.A(_11925_));
 sg13g2_antennanp ANTENNA_2804 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2805 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2806 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2807 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2808 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2809 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2810 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2811 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2812 (.A(_11938_));
 sg13g2_antennanp ANTENNA_2813 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2814 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2815 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2816 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2817 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2818 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2819 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2820 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2821 (.A(_11945_));
 sg13g2_antennanp ANTENNA_2822 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2823 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2824 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2825 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2826 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2827 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2828 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2829 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2830 (.A(_11974_));
 sg13g2_antennanp ANTENNA_2831 (.A(clk));
 sg13g2_antennanp ANTENNA_2832 (.A(clk));
 sg13g2_antennanp ANTENNA_2833 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2834 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2835 (.A(net3));
 sg13g2_antennanp ANTENNA_2836 (.A(net3));
 sg13g2_antennanp ANTENNA_2837 (.A(net3));
 sg13g2_antennanp ANTENNA_2838 (.A(net19));
 sg13g2_antennanp ANTENNA_2839 (.A(net19));
 sg13g2_antennanp ANTENNA_2840 (.A(net151));
 sg13g2_antennanp ANTENNA_2841 (.A(net151));
 sg13g2_antennanp ANTENNA_2842 (.A(net151));
 sg13g2_antennanp ANTENNA_2843 (.A(net151));
 sg13g2_antennanp ANTENNA_2844 (.A(net151));
 sg13g2_antennanp ANTENNA_2845 (.A(net151));
 sg13g2_antennanp ANTENNA_2846 (.A(net151));
 sg13g2_antennanp ANTENNA_2847 (.A(net151));
 sg13g2_antennanp ANTENNA_2848 (.A(net151));
 sg13g2_antennanp ANTENNA_2849 (.A(net366));
 sg13g2_antennanp ANTENNA_2850 (.A(net366));
 sg13g2_antennanp ANTENNA_2851 (.A(net366));
 sg13g2_antennanp ANTENNA_2852 (.A(net366));
 sg13g2_antennanp ANTENNA_2853 (.A(net366));
 sg13g2_antennanp ANTENNA_2854 (.A(net366));
 sg13g2_antennanp ANTENNA_2855 (.A(net366));
 sg13g2_antennanp ANTENNA_2856 (.A(net366));
 sg13g2_antennanp ANTENNA_2857 (.A(net366));
 sg13g2_antennanp ANTENNA_2858 (.A(net366));
 sg13g2_antennanp ANTENNA_2859 (.A(net366));
 sg13g2_antennanp ANTENNA_2860 (.A(net366));
 sg13g2_antennanp ANTENNA_2861 (.A(net366));
 sg13g2_antennanp ANTENNA_2862 (.A(net366));
 sg13g2_antennanp ANTENNA_2863 (.A(net366));
 sg13g2_antennanp ANTENNA_2864 (.A(net366));
 sg13g2_antennanp ANTENNA_2865 (.A(net366));
 sg13g2_antennanp ANTENNA_2866 (.A(net366));
 sg13g2_antennanp ANTENNA_2867 (.A(net366));
 sg13g2_antennanp ANTENNA_2868 (.A(net366));
 sg13g2_antennanp ANTENNA_2869 (.A(net366));
 sg13g2_antennanp ANTENNA_2870 (.A(net366));
 sg13g2_antennanp ANTENNA_2871 (.A(net366));
 sg13g2_antennanp ANTENNA_2872 (.A(net366));
 sg13g2_antennanp ANTENNA_2873 (.A(net366));
 sg13g2_antennanp ANTENNA_2874 (.A(net366));
 sg13g2_antennanp ANTENNA_2875 (.A(net366));
 sg13g2_antennanp ANTENNA_2876 (.A(net366));
 sg13g2_antennanp ANTENNA_2877 (.A(net366));
 sg13g2_antennanp ANTENNA_2878 (.A(net366));
 sg13g2_antennanp ANTENNA_2879 (.A(net366));
 sg13g2_antennanp ANTENNA_2880 (.A(net366));
 sg13g2_antennanp ANTENNA_2881 (.A(net366));
 sg13g2_antennanp ANTENNA_2882 (.A(net366));
 sg13g2_antennanp ANTENNA_2883 (.A(net468));
 sg13g2_antennanp ANTENNA_2884 (.A(net468));
 sg13g2_antennanp ANTENNA_2885 (.A(net468));
 sg13g2_antennanp ANTENNA_2886 (.A(net468));
 sg13g2_antennanp ANTENNA_2887 (.A(net468));
 sg13g2_antennanp ANTENNA_2888 (.A(net468));
 sg13g2_antennanp ANTENNA_2889 (.A(net468));
 sg13g2_antennanp ANTENNA_2890 (.A(net468));
 sg13g2_antennanp ANTENNA_2891 (.A(net468));
 sg13g2_antennanp ANTENNA_2892 (.A(net643));
 sg13g2_antennanp ANTENNA_2893 (.A(net643));
 sg13g2_antennanp ANTENNA_2894 (.A(net643));
 sg13g2_antennanp ANTENNA_2895 (.A(net643));
 sg13g2_antennanp ANTENNA_2896 (.A(net643));
 sg13g2_antennanp ANTENNA_2897 (.A(net643));
 sg13g2_antennanp ANTENNA_2898 (.A(net643));
 sg13g2_antennanp ANTENNA_2899 (.A(net643));
 sg13g2_antennanp ANTENNA_2900 (.A(net643));
 sg13g2_antennanp ANTENNA_2901 (.A(net643));
 sg13g2_antennanp ANTENNA_2902 (.A(net643));
 sg13g2_antennanp ANTENNA_2903 (.A(net643));
 sg13g2_antennanp ANTENNA_2904 (.A(net643));
 sg13g2_antennanp ANTENNA_2905 (.A(net643));
 sg13g2_antennanp ANTENNA_2906 (.A(net643));
 sg13g2_antennanp ANTENNA_2907 (.A(net643));
 sg13g2_antennanp ANTENNA_2908 (.A(net643));
 sg13g2_antennanp ANTENNA_2909 (.A(net643));
 sg13g2_antennanp ANTENNA_2910 (.A(net643));
 sg13g2_antennanp ANTENNA_2911 (.A(net643));
 sg13g2_antennanp ANTENNA_2912 (.A(net643));
 sg13g2_antennanp ANTENNA_2913 (.A(net643));
 sg13g2_antennanp ANTENNA_2914 (.A(net643));
 sg13g2_antennanp ANTENNA_2915 (.A(net643));
 sg13g2_antennanp ANTENNA_2916 (.A(net643));
 sg13g2_antennanp ANTENNA_2917 (.A(net643));
 sg13g2_antennanp ANTENNA_2918 (.A(net643));
 sg13g2_antennanp ANTENNA_2919 (.A(net643));
 sg13g2_antennanp ANTENNA_2920 (.A(net643));
 sg13g2_antennanp ANTENNA_2921 (.A(net643));
 sg13g2_antennanp ANTENNA_2922 (.A(net643));
 sg13g2_antennanp ANTENNA_2923 (.A(net643));
 sg13g2_antennanp ANTENNA_2924 (.A(net643));
 sg13g2_antennanp ANTENNA_2925 (.A(net643));
 sg13g2_antennanp ANTENNA_2926 (.A(net667));
 sg13g2_antennanp ANTENNA_2927 (.A(net667));
 sg13g2_antennanp ANTENNA_2928 (.A(net667));
 sg13g2_antennanp ANTENNA_2929 (.A(net667));
 sg13g2_antennanp ANTENNA_2930 (.A(net667));
 sg13g2_antennanp ANTENNA_2931 (.A(net667));
 sg13g2_antennanp ANTENNA_2932 (.A(net667));
 sg13g2_antennanp ANTENNA_2933 (.A(net667));
 sg13g2_antennanp ANTENNA_2934 (.A(net667));
 sg13g2_antennanp ANTENNA_2935 (.A(net667));
 sg13g2_antennanp ANTENNA_2936 (.A(net667));
 sg13g2_antennanp ANTENNA_2937 (.A(net667));
 sg13g2_antennanp ANTENNA_2938 (.A(net667));
 sg13g2_antennanp ANTENNA_2939 (.A(net667));
 sg13g2_antennanp ANTENNA_2940 (.A(net667));
 sg13g2_antennanp ANTENNA_2941 (.A(net679));
 sg13g2_antennanp ANTENNA_2942 (.A(net679));
 sg13g2_antennanp ANTENNA_2943 (.A(net679));
 sg13g2_antennanp ANTENNA_2944 (.A(net679));
 sg13g2_antennanp ANTENNA_2945 (.A(net679));
 sg13g2_antennanp ANTENNA_2946 (.A(net679));
 sg13g2_antennanp ANTENNA_2947 (.A(net679));
 sg13g2_antennanp ANTENNA_2948 (.A(net679));
 sg13g2_antennanp ANTENNA_2949 (.A(net679));
 sg13g2_antennanp ANTENNA_2950 (.A(net796));
 sg13g2_antennanp ANTENNA_2951 (.A(net796));
 sg13g2_antennanp ANTENNA_2952 (.A(net796));
 sg13g2_antennanp ANTENNA_2953 (.A(net796));
 sg13g2_antennanp ANTENNA_2954 (.A(net796));
 sg13g2_antennanp ANTENNA_2955 (.A(net796));
 sg13g2_antennanp ANTENNA_2956 (.A(net796));
 sg13g2_antennanp ANTENNA_2957 (.A(net796));
 sg13g2_antennanp ANTENNA_2958 (.A(net848));
 sg13g2_antennanp ANTENNA_2959 (.A(net848));
 sg13g2_antennanp ANTENNA_2960 (.A(net848));
 sg13g2_antennanp ANTENNA_2961 (.A(net848));
 sg13g2_antennanp ANTENNA_2962 (.A(net848));
 sg13g2_antennanp ANTENNA_2963 (.A(net848));
 sg13g2_antennanp ANTENNA_2964 (.A(net848));
 sg13g2_antennanp ANTENNA_2965 (.A(net848));
 sg13g2_antennanp ANTENNA_2966 (.A(net848));
 sg13g2_antennanp ANTENNA_2967 (.A(net853));
 sg13g2_antennanp ANTENNA_2968 (.A(net853));
 sg13g2_antennanp ANTENNA_2969 (.A(net853));
 sg13g2_antennanp ANTENNA_2970 (.A(net853));
 sg13g2_antennanp ANTENNA_2971 (.A(net853));
 sg13g2_antennanp ANTENNA_2972 (.A(net853));
 sg13g2_antennanp ANTENNA_2973 (.A(net853));
 sg13g2_antennanp ANTENNA_2974 (.A(net853));
 sg13g2_antennanp ANTENNA_2975 (.A(net853));
 sg13g2_antennanp ANTENNA_2976 (.A(net853));
 sg13g2_antennanp ANTENNA_2977 (.A(net853));
 sg13g2_antennanp ANTENNA_2978 (.A(net853));
 sg13g2_antennanp ANTENNA_2979 (.A(net853));
 sg13g2_antennanp ANTENNA_2980 (.A(net853));
 sg13g2_antennanp ANTENNA_2981 (.A(net853));
 sg13g2_antennanp ANTENNA_2982 (.A(net853));
 sg13g2_antennanp ANTENNA_2983 (.A(net853));
 sg13g2_antennanp ANTENNA_2984 (.A(net853));
 sg13g2_antennanp ANTENNA_2985 (.A(net853));
 sg13g2_antennanp ANTENNA_2986 (.A(net853));
 sg13g2_antennanp ANTENNA_2987 (.A(net853));
 sg13g2_antennanp ANTENNA_2988 (.A(net853));
 sg13g2_antennanp ANTENNA_2989 (.A(net956));
 sg13g2_antennanp ANTENNA_2990 (.A(net956));
 sg13g2_antennanp ANTENNA_2991 (.A(net956));
 sg13g2_antennanp ANTENNA_2992 (.A(net956));
 sg13g2_antennanp ANTENNA_2993 (.A(net956));
 sg13g2_antennanp ANTENNA_2994 (.A(net956));
 sg13g2_antennanp ANTENNA_2995 (.A(net956));
 sg13g2_antennanp ANTENNA_2996 (.A(net956));
 sg13g2_antennanp ANTENNA_2997 (.A(net956));
 sg13g2_antennanp ANTENNA_2998 (.A(net958));
 sg13g2_antennanp ANTENNA_2999 (.A(net958));
 sg13g2_antennanp ANTENNA_3000 (.A(net958));
 sg13g2_antennanp ANTENNA_3001 (.A(net958));
 sg13g2_antennanp ANTENNA_3002 (.A(net958));
 sg13g2_antennanp ANTENNA_3003 (.A(net958));
 sg13g2_antennanp ANTENNA_3004 (.A(net958));
 sg13g2_antennanp ANTENNA_3005 (.A(net958));
 sg13g2_antennanp ANTENNA_3006 (.A(net986));
 sg13g2_antennanp ANTENNA_3007 (.A(net986));
 sg13g2_antennanp ANTENNA_3008 (.A(net986));
 sg13g2_antennanp ANTENNA_3009 (.A(net986));
 sg13g2_antennanp ANTENNA_3010 (.A(net986));
 sg13g2_antennanp ANTENNA_3011 (.A(net986));
 sg13g2_antennanp ANTENNA_3012 (.A(net986));
 sg13g2_antennanp ANTENNA_3013 (.A(net986));
 sg13g2_antennanp ANTENNA_3014 (.A(net991));
 sg13g2_antennanp ANTENNA_3015 (.A(net991));
 sg13g2_antennanp ANTENNA_3016 (.A(net991));
 sg13g2_antennanp ANTENNA_3017 (.A(net991));
 sg13g2_antennanp ANTENNA_3018 (.A(net991));
 sg13g2_antennanp ANTENNA_3019 (.A(net991));
 sg13g2_antennanp ANTENNA_3020 (.A(net991));
 sg13g2_antennanp ANTENNA_3021 (.A(net991));
 sg13g2_antennanp ANTENNA_3022 (.A(net991));
 sg13g2_antennanp ANTENNA_3023 (.A(net1038));
 sg13g2_antennanp ANTENNA_3024 (.A(net1038));
 sg13g2_antennanp ANTENNA_3025 (.A(net1038));
 sg13g2_antennanp ANTENNA_3026 (.A(net1038));
 sg13g2_antennanp ANTENNA_3027 (.A(net1038));
 sg13g2_antennanp ANTENNA_3028 (.A(net1038));
 sg13g2_antennanp ANTENNA_3029 (.A(net1038));
 sg13g2_antennanp ANTENNA_3030 (.A(net1038));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_fill_1 FILLER_0_70 ();
 sg13g2_fill_2 FILLER_0_97 ();
 sg13g2_decap_4 FILLER_0_103 ();
 sg13g2_fill_2 FILLER_0_107 ();
 sg13g2_decap_4 FILLER_0_113 ();
 sg13g2_fill_2 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_4 FILLER_0_130 ();
 sg13g2_fill_2 FILLER_0_134 ();
 sg13g2_fill_2 FILLER_0_146 ();
 sg13g2_fill_1 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_153 ();
 sg13g2_fill_2 FILLER_0_160 ();
 sg13g2_fill_1 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_167 ();
 sg13g2_decap_8 FILLER_0_174 ();
 sg13g2_decap_8 FILLER_0_181 ();
 sg13g2_fill_1 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_4 FILLER_0_214 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_decap_4 FILLER_0_223 ();
 sg13g2_fill_2 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_fill_2 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_fill_2 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_4 FILLER_0_307 ();
 sg13g2_fill_2 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_4 FILLER_0_385 ();
 sg13g2_fill_2 FILLER_0_389 ();
 sg13g2_decap_4 FILLER_0_395 ();
 sg13g2_fill_2 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_4 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_fill_1 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_454 ();
 sg13g2_decap_8 FILLER_0_461 ();
 sg13g2_decap_4 FILLER_0_482 ();
 sg13g2_fill_2 FILLER_0_489 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_524 ();
 sg13g2_decap_8 FILLER_0_531 ();
 sg13g2_decap_8 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_545 ();
 sg13g2_decap_8 FILLER_0_552 ();
 sg13g2_decap_8 FILLER_0_559 ();
 sg13g2_fill_1 FILLER_0_566 ();
 sg13g2_decap_8 FILLER_0_571 ();
 sg13g2_decap_8 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_fill_1 FILLER_0_678 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_fill_1 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_fill_2 FILLER_0_757 ();
 sg13g2_fill_1 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_fill_2 FILLER_0_777 ();
 sg13g2_fill_1 FILLER_0_779 ();
 sg13g2_fill_1 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_fill_2 FILLER_0_802 ();
 sg13g2_decap_4 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_844 ();
 sg13g2_decap_8 FILLER_0_851 ();
 sg13g2_decap_8 FILLER_0_858 ();
 sg13g2_fill_1 FILLER_0_865 ();
 sg13g2_decap_8 FILLER_0_870 ();
 sg13g2_decap_8 FILLER_0_877 ();
 sg13g2_decap_4 FILLER_0_884 ();
 sg13g2_fill_1 FILLER_0_888 ();
 sg13g2_fill_2 FILLER_0_928 ();
 sg13g2_fill_1 FILLER_0_930 ();
 sg13g2_decap_8 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_971 ();
 sg13g2_fill_2 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_fill_2 FILLER_0_1013 ();
 sg13g2_decap_4 FILLER_0_1055 ();
 sg13g2_fill_1 FILLER_0_1059 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_fill_1 FILLER_0_1071 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1100 ();
 sg13g2_decap_8 FILLER_0_1107 ();
 sg13g2_decap_8 FILLER_0_1114 ();
 sg13g2_decap_8 FILLER_0_1121 ();
 sg13g2_decap_8 FILLER_0_1128 ();
 sg13g2_decap_8 FILLER_0_1135 ();
 sg13g2_decap_4 FILLER_0_1142 ();
 sg13g2_fill_2 FILLER_0_1146 ();
 sg13g2_fill_1 FILLER_0_1152 ();
 sg13g2_fill_2 FILLER_0_1162 ();
 sg13g2_fill_2 FILLER_0_1168 ();
 sg13g2_fill_1 FILLER_0_1174 ();
 sg13g2_fill_1 FILLER_0_1180 ();
 sg13g2_decap_8 FILLER_0_1185 ();
 sg13g2_decap_8 FILLER_0_1192 ();
 sg13g2_decap_8 FILLER_0_1199 ();
 sg13g2_decap_8 FILLER_0_1206 ();
 sg13g2_decap_8 FILLER_0_1213 ();
 sg13g2_decap_8 FILLER_0_1220 ();
 sg13g2_decap_4 FILLER_0_1227 ();
 sg13g2_fill_2 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1241 ();
 sg13g2_fill_2 FILLER_0_1248 ();
 sg13g2_decap_8 FILLER_0_1254 ();
 sg13g2_decap_8 FILLER_0_1261 ();
 sg13g2_decap_8 FILLER_0_1268 ();
 sg13g2_decap_8 FILLER_0_1275 ();
 sg13g2_decap_8 FILLER_0_1282 ();
 sg13g2_decap_8 FILLER_0_1319 ();
 sg13g2_decap_4 FILLER_0_1326 ();
 sg13g2_fill_2 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_fill_2 FILLER_0_1372 ();
 sg13g2_fill_1 FILLER_0_1374 ();
 sg13g2_fill_1 FILLER_0_1388 ();
 sg13g2_decap_4 FILLER_0_1403 ();
 sg13g2_fill_2 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1439 ();
 sg13g2_decap_8 FILLER_0_1446 ();
 sg13g2_decap_8 FILLER_0_1453 ();
 sg13g2_fill_2 FILLER_0_1460 ();
 sg13g2_fill_1 FILLER_0_1462 ();
 sg13g2_decap_8 FILLER_0_1481 ();
 sg13g2_decap_8 FILLER_0_1488 ();
 sg13g2_decap_8 FILLER_0_1495 ();
 sg13g2_decap_8 FILLER_0_1502 ();
 sg13g2_decap_4 FILLER_0_1509 ();
 sg13g2_fill_2 FILLER_0_1513 ();
 sg13g2_decap_8 FILLER_0_1545 ();
 sg13g2_decap_8 FILLER_0_1552 ();
 sg13g2_decap_8 FILLER_0_1559 ();
 sg13g2_fill_2 FILLER_0_1566 ();
 sg13g2_decap_8 FILLER_0_1572 ();
 sg13g2_decap_8 FILLER_0_1579 ();
 sg13g2_decap_8 FILLER_0_1586 ();
 sg13g2_decap_8 FILLER_0_1610 ();
 sg13g2_decap_8 FILLER_0_1617 ();
 sg13g2_decap_8 FILLER_0_1624 ();
 sg13g2_decap_8 FILLER_0_1631 ();
 sg13g2_fill_1 FILLER_0_1638 ();
 sg13g2_decap_8 FILLER_0_1665 ();
 sg13g2_decap_4 FILLER_0_1672 ();
 sg13g2_fill_1 FILLER_0_1676 ();
 sg13g2_decap_8 FILLER_0_1703 ();
 sg13g2_fill_1 FILLER_0_1710 ();
 sg13g2_fill_2 FILLER_0_1719 ();
 sg13g2_decap_8 FILLER_0_1734 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_4 FILLER_0_1762 ();
 sg13g2_fill_2 FILLER_0_1766 ();
 sg13g2_decap_8 FILLER_0_1794 ();
 sg13g2_fill_1 FILLER_0_1801 ();
 sg13g2_decap_8 FILLER_0_1816 ();
 sg13g2_decap_8 FILLER_0_1823 ();
 sg13g2_decap_8 FILLER_0_1830 ();
 sg13g2_decap_8 FILLER_0_1837 ();
 sg13g2_decap_4 FILLER_0_1858 ();
 sg13g2_fill_2 FILLER_0_1862 ();
 sg13g2_decap_8 FILLER_0_1874 ();
 sg13g2_decap_8 FILLER_0_1881 ();
 sg13g2_decap_8 FILLER_0_1888 ();
 sg13g2_decap_8 FILLER_0_1895 ();
 sg13g2_decap_8 FILLER_0_1902 ();
 sg13g2_decap_4 FILLER_0_1909 ();
 sg13g2_fill_2 FILLER_0_1913 ();
 sg13g2_decap_8 FILLER_0_1929 ();
 sg13g2_decap_8 FILLER_0_1936 ();
 sg13g2_fill_1 FILLER_0_1943 ();
 sg13g2_decap_8 FILLER_0_1948 ();
 sg13g2_decap_4 FILLER_0_1955 ();
 sg13g2_fill_1 FILLER_0_1959 ();
 sg13g2_fill_1 FILLER_0_1964 ();
 sg13g2_decap_8 FILLER_0_1969 ();
 sg13g2_decap_8 FILLER_0_1976 ();
 sg13g2_decap_4 FILLER_0_1983 ();
 sg13g2_decap_8 FILLER_0_2013 ();
 sg13g2_decap_8 FILLER_0_2020 ();
 sg13g2_decap_8 FILLER_0_2027 ();
 sg13g2_fill_2 FILLER_0_2034 ();
 sg13g2_decap_8 FILLER_0_2046 ();
 sg13g2_decap_8 FILLER_0_2074 ();
 sg13g2_decap_8 FILLER_0_2081 ();
 sg13g2_decap_8 FILLER_0_2088 ();
 sg13g2_decap_8 FILLER_0_2095 ();
 sg13g2_decap_8 FILLER_0_2132 ();
 sg13g2_decap_8 FILLER_0_2139 ();
 sg13g2_decap_8 FILLER_0_2146 ();
 sg13g2_decap_4 FILLER_0_2153 ();
 sg13g2_fill_2 FILLER_0_2157 ();
 sg13g2_decap_8 FILLER_0_2185 ();
 sg13g2_decap_4 FILLER_0_2192 ();
 sg13g2_decap_8 FILLER_0_2226 ();
 sg13g2_decap_8 FILLER_0_2233 ();
 sg13g2_decap_8 FILLER_0_2240 ();
 sg13g2_decap_8 FILLER_0_2251 ();
 sg13g2_decap_8 FILLER_0_2258 ();
 sg13g2_decap_4 FILLER_0_2265 ();
 sg13g2_fill_2 FILLER_0_2269 ();
 sg13g2_decap_4 FILLER_0_2281 ();
 sg13g2_fill_2 FILLER_0_2289 ();
 sg13g2_decap_8 FILLER_0_2301 ();
 sg13g2_decap_8 FILLER_0_2308 ();
 sg13g2_decap_8 FILLER_0_2315 ();
 sg13g2_decap_8 FILLER_0_2322 ();
 sg13g2_decap_8 FILLER_0_2349 ();
 sg13g2_decap_8 FILLER_0_2356 ();
 sg13g2_decap_8 FILLER_0_2363 ();
 sg13g2_decap_8 FILLER_0_2370 ();
 sg13g2_decap_8 FILLER_0_2377 ();
 sg13g2_decap_8 FILLER_0_2384 ();
 sg13g2_decap_8 FILLER_0_2391 ();
 sg13g2_decap_8 FILLER_0_2398 ();
 sg13g2_decap_8 FILLER_0_2405 ();
 sg13g2_decap_8 FILLER_0_2412 ();
 sg13g2_decap_8 FILLER_0_2419 ();
 sg13g2_decap_8 FILLER_0_2426 ();
 sg13g2_decap_8 FILLER_0_2433 ();
 sg13g2_decap_8 FILLER_0_2440 ();
 sg13g2_decap_8 FILLER_0_2447 ();
 sg13g2_decap_8 FILLER_0_2454 ();
 sg13g2_decap_8 FILLER_0_2461 ();
 sg13g2_decap_8 FILLER_0_2468 ();
 sg13g2_decap_8 FILLER_0_2475 ();
 sg13g2_decap_8 FILLER_0_2482 ();
 sg13g2_decap_8 FILLER_0_2489 ();
 sg13g2_decap_8 FILLER_0_2496 ();
 sg13g2_decap_8 FILLER_0_2503 ();
 sg13g2_decap_8 FILLER_0_2510 ();
 sg13g2_decap_8 FILLER_0_2517 ();
 sg13g2_decap_8 FILLER_0_2524 ();
 sg13g2_decap_8 FILLER_0_2531 ();
 sg13g2_decap_8 FILLER_0_2538 ();
 sg13g2_decap_8 FILLER_0_2545 ();
 sg13g2_decap_8 FILLER_0_2552 ();
 sg13g2_decap_8 FILLER_0_2559 ();
 sg13g2_decap_8 FILLER_0_2566 ();
 sg13g2_decap_8 FILLER_0_2573 ();
 sg13g2_decap_8 FILLER_0_2580 ();
 sg13g2_decap_8 FILLER_0_2587 ();
 sg13g2_decap_8 FILLER_0_2594 ();
 sg13g2_decap_8 FILLER_0_2601 ();
 sg13g2_decap_8 FILLER_0_2608 ();
 sg13g2_decap_8 FILLER_0_2615 ();
 sg13g2_decap_8 FILLER_0_2622 ();
 sg13g2_decap_8 FILLER_0_2629 ();
 sg13g2_decap_8 FILLER_0_2636 ();
 sg13g2_decap_8 FILLER_0_2643 ();
 sg13g2_decap_8 FILLER_0_2650 ();
 sg13g2_decap_8 FILLER_0_2657 ();
 sg13g2_decap_4 FILLER_0_2664 ();
 sg13g2_fill_2 FILLER_0_2668 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_fill_2 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_148 ();
 sg13g2_fill_2 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_210 ();
 sg13g2_fill_1 FILLER_1_263 ();
 sg13g2_fill_1 FILLER_1_320 ();
 sg13g2_fill_1 FILLER_1_325 ();
 sg13g2_fill_1 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_fill_2 FILLER_1_420 ();
 sg13g2_fill_1 FILLER_1_422 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_4 FILLER_1_511 ();
 sg13g2_fill_2 FILLER_1_515 ();
 sg13g2_decap_8 FILLER_1_543 ();
 sg13g2_fill_2 FILLER_1_550 ();
 sg13g2_fill_1 FILLER_1_552 ();
 sg13g2_fill_2 FILLER_1_594 ();
 sg13g2_fill_2 FILLER_1_604 ();
 sg13g2_fill_1 FILLER_1_606 ();
 sg13g2_decap_4 FILLER_1_611 ();
 sg13g2_fill_1 FILLER_1_615 ();
 sg13g2_decap_8 FILLER_1_620 ();
 sg13g2_decap_4 FILLER_1_627 ();
 sg13g2_fill_1 FILLER_1_631 ();
 sg13g2_fill_2 FILLER_1_661 ();
 sg13g2_decap_8 FILLER_1_703 ();
 sg13g2_fill_1 FILLER_1_710 ();
 sg13g2_fill_2 FILLER_1_737 ();
 sg13g2_fill_1 FILLER_1_739 ();
 sg13g2_decap_8 FILLER_1_766 ();
 sg13g2_fill_1 FILLER_1_799 ();
 sg13g2_decap_4 FILLER_1_840 ();
 sg13g2_fill_2 FILLER_1_932 ();
 sg13g2_decap_4 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_1014 ();
 sg13g2_fill_2 FILLER_1_1051 ();
 sg13g2_fill_2 FILLER_1_1079 ();
 sg13g2_fill_1 FILLER_1_1081 ();
 sg13g2_fill_1 FILLER_1_1108 ();
 sg13g2_fill_2 FILLER_1_1135 ();
 sg13g2_fill_1 FILLER_1_1137 ();
 sg13g2_fill_2 FILLER_1_1199 ();
 sg13g2_decap_8 FILLER_1_1205 ();
 sg13g2_fill_2 FILLER_1_1212 ();
 sg13g2_fill_2 FILLER_1_1223 ();
 sg13g2_fill_1 FILLER_1_1230 ();
 sg13g2_fill_2 FILLER_1_1261 ();
 sg13g2_decap_8 FILLER_1_1361 ();
 sg13g2_decap_8 FILLER_1_1368 ();
 sg13g2_fill_2 FILLER_1_1375 ();
 sg13g2_fill_1 FILLER_1_1377 ();
 sg13g2_fill_2 FILLER_1_1404 ();
 sg13g2_decap_4 FILLER_1_1420 ();
 sg13g2_fill_2 FILLER_1_1424 ();
 sg13g2_decap_8 FILLER_1_1452 ();
 sg13g2_decap_8 FILLER_1_1459 ();
 sg13g2_fill_2 FILLER_1_1466 ();
 sg13g2_fill_1 FILLER_1_1468 ();
 sg13g2_decap_4 FILLER_1_1495 ();
 sg13g2_decap_4 FILLER_1_1520 ();
 sg13g2_decap_8 FILLER_1_1528 ();
 sg13g2_decap_8 FILLER_1_1535 ();
 sg13g2_fill_1 FILLER_1_1542 ();
 sg13g2_fill_1 FILLER_1_1577 ();
 sg13g2_decap_4 FILLER_1_1612 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_decap_4 FILLER_1_1631 ();
 sg13g2_decap_8 FILLER_1_1695 ();
 sg13g2_decap_4 FILLER_1_1702 ();
 sg13g2_fill_2 FILLER_1_1706 ();
 sg13g2_fill_1 FILLER_1_1800 ();
 sg13g2_decap_8 FILLER_1_1827 ();
 sg13g2_fill_1 FILLER_1_1834 ();
 sg13g2_fill_1 FILLER_1_1861 ();
 sg13g2_fill_1 FILLER_1_1866 ();
 sg13g2_fill_1 FILLER_1_1943 ();
 sg13g2_fill_1 FILLER_1_1948 ();
 sg13g2_fill_2 FILLER_1_1979 ();
 sg13g2_decap_4 FILLER_1_1991 ();
 sg13g2_decap_4 FILLER_1_1999 ();
 sg13g2_fill_2 FILLER_1_2003 ();
 sg13g2_decap_4 FILLER_1_2015 ();
 sg13g2_decap_4 FILLER_1_2033 ();
 sg13g2_fill_1 FILLER_1_2037 ();
 sg13g2_fill_1 FILLER_1_2110 ();
 sg13g2_decap_8 FILLER_1_2132 ();
 sg13g2_decap_4 FILLER_1_2139 ();
 sg13g2_fill_1 FILLER_1_2143 ();
 sg13g2_decap_4 FILLER_1_2164 ();
 sg13g2_fill_1 FILLER_1_2168 ();
 sg13g2_decap_8 FILLER_1_2194 ();
 sg13g2_fill_1 FILLER_1_2221 ();
 sg13g2_fill_2 FILLER_1_2239 ();
 sg13g2_decap_8 FILLER_1_2267 ();
 sg13g2_fill_2 FILLER_1_2274 ();
 sg13g2_fill_1 FILLER_1_2326 ();
 sg13g2_decap_8 FILLER_1_2357 ();
 sg13g2_decap_8 FILLER_1_2364 ();
 sg13g2_fill_1 FILLER_1_2371 ();
 sg13g2_decap_8 FILLER_1_2408 ();
 sg13g2_decap_8 FILLER_1_2415 ();
 sg13g2_decap_8 FILLER_1_2422 ();
 sg13g2_decap_8 FILLER_1_2429 ();
 sg13g2_decap_8 FILLER_1_2436 ();
 sg13g2_decap_8 FILLER_1_2443 ();
 sg13g2_decap_8 FILLER_1_2450 ();
 sg13g2_decap_8 FILLER_1_2457 ();
 sg13g2_decap_8 FILLER_1_2464 ();
 sg13g2_decap_8 FILLER_1_2471 ();
 sg13g2_decap_8 FILLER_1_2478 ();
 sg13g2_decap_8 FILLER_1_2485 ();
 sg13g2_decap_8 FILLER_1_2492 ();
 sg13g2_decap_8 FILLER_1_2499 ();
 sg13g2_decap_8 FILLER_1_2506 ();
 sg13g2_decap_8 FILLER_1_2513 ();
 sg13g2_decap_8 FILLER_1_2520 ();
 sg13g2_decap_8 FILLER_1_2527 ();
 sg13g2_decap_8 FILLER_1_2534 ();
 sg13g2_decap_8 FILLER_1_2541 ();
 sg13g2_decap_8 FILLER_1_2548 ();
 sg13g2_decap_8 FILLER_1_2555 ();
 sg13g2_decap_8 FILLER_1_2562 ();
 sg13g2_decap_8 FILLER_1_2569 ();
 sg13g2_decap_8 FILLER_1_2576 ();
 sg13g2_decap_8 FILLER_1_2583 ();
 sg13g2_decap_8 FILLER_1_2590 ();
 sg13g2_decap_8 FILLER_1_2597 ();
 sg13g2_decap_8 FILLER_1_2604 ();
 sg13g2_decap_8 FILLER_1_2611 ();
 sg13g2_decap_8 FILLER_1_2618 ();
 sg13g2_decap_8 FILLER_1_2625 ();
 sg13g2_decap_8 FILLER_1_2632 ();
 sg13g2_decap_8 FILLER_1_2639 ();
 sg13g2_decap_8 FILLER_1_2646 ();
 sg13g2_decap_8 FILLER_1_2653 ();
 sg13g2_decap_8 FILLER_1_2660 ();
 sg13g2_fill_2 FILLER_1_2667 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_decap_4 FILLER_2_84 ();
 sg13g2_fill_1 FILLER_2_148 ();
 sg13g2_fill_1 FILLER_2_175 ();
 sg13g2_fill_1 FILLER_2_212 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_fill_1 FILLER_2_301 ();
 sg13g2_fill_2 FILLER_2_328 ();
 sg13g2_fill_2 FILLER_2_335 ();
 sg13g2_fill_1 FILLER_2_337 ();
 sg13g2_fill_1 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_412 ();
 sg13g2_fill_1 FILLER_2_414 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_fill_2 FILLER_2_439 ();
 sg13g2_fill_1 FILLER_2_441 ();
 sg13g2_fill_1 FILLER_2_507 ();
 sg13g2_fill_1 FILLER_2_548 ();
 sg13g2_decap_8 FILLER_2_646 ();
 sg13g2_fill_2 FILLER_2_653 ();
 sg13g2_fill_1 FILLER_2_689 ();
 sg13g2_fill_1 FILLER_2_700 ();
 sg13g2_fill_2 FILLER_2_721 ();
 sg13g2_fill_1 FILLER_2_723 ();
 sg13g2_decap_8 FILLER_2_727 ();
 sg13g2_decap_4 FILLER_2_734 ();
 sg13g2_fill_2 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_975 ();
 sg13g2_decap_8 FILLER_2_982 ();
 sg13g2_fill_2 FILLER_2_999 ();
 sg13g2_fill_1 FILLER_2_1001 ();
 sg13g2_fill_2 FILLER_2_1033 ();
 sg13g2_fill_1 FILLER_2_1094 ();
 sg13g2_fill_1 FILLER_2_1121 ();
 sg13g2_fill_2 FILLER_2_1148 ();
 sg13g2_fill_2 FILLER_2_1250 ();
 sg13g2_fill_1 FILLER_2_1252 ();
 sg13g2_fill_1 FILLER_2_1278 ();
 sg13g2_fill_2 FILLER_2_1306 ();
 sg13g2_fill_2 FILLER_2_1334 ();
 sg13g2_decap_8 FILLER_2_1366 ();
 sg13g2_fill_1 FILLER_2_1373 ();
 sg13g2_fill_2 FILLER_2_1436 ();
 sg13g2_decap_8 FILLER_2_1442 ();
 sg13g2_fill_2 FILLER_2_1449 ();
 sg13g2_decap_4 FILLER_2_1569 ();
 sg13g2_fill_2 FILLER_2_1649 ();
 sg13g2_fill_1 FILLER_2_1659 ();
 sg13g2_fill_1 FILLER_2_1664 ();
 sg13g2_fill_1 FILLER_2_1695 ();
 sg13g2_decap_8 FILLER_2_1700 ();
 sg13g2_fill_1 FILLER_2_1745 ();
 sg13g2_decap_8 FILLER_2_1750 ();
 sg13g2_decap_4 FILLER_2_1757 ();
 sg13g2_fill_1 FILLER_2_1801 ();
 sg13g2_fill_1 FILLER_2_1828 ();
 sg13g2_fill_2 FILLER_2_1881 ();
 sg13g2_fill_1 FILLER_2_1992 ();
 sg13g2_fill_1 FILLER_2_2019 ();
 sg13g2_fill_1 FILLER_2_2046 ();
 sg13g2_fill_1 FILLER_2_2073 ();
 sg13g2_decap_4 FILLER_2_2108 ();
 sg13g2_fill_2 FILLER_2_2138 ();
 sg13g2_fill_1 FILLER_2_2170 ();
 sg13g2_fill_1 FILLER_2_2197 ();
 sg13g2_fill_1 FILLER_2_2224 ();
 sg13g2_fill_1 FILLER_2_2313 ();
 sg13g2_decap_8 FILLER_2_2406 ();
 sg13g2_decap_8 FILLER_2_2413 ();
 sg13g2_decap_8 FILLER_2_2420 ();
 sg13g2_decap_8 FILLER_2_2427 ();
 sg13g2_decap_8 FILLER_2_2434 ();
 sg13g2_decap_8 FILLER_2_2441 ();
 sg13g2_decap_8 FILLER_2_2448 ();
 sg13g2_decap_8 FILLER_2_2455 ();
 sg13g2_decap_8 FILLER_2_2462 ();
 sg13g2_decap_8 FILLER_2_2469 ();
 sg13g2_decap_8 FILLER_2_2476 ();
 sg13g2_decap_8 FILLER_2_2483 ();
 sg13g2_decap_8 FILLER_2_2490 ();
 sg13g2_decap_8 FILLER_2_2497 ();
 sg13g2_decap_8 FILLER_2_2504 ();
 sg13g2_decap_8 FILLER_2_2511 ();
 sg13g2_decap_8 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2525 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_8 FILLER_2_2539 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_4 FILLER_2_2665 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_128 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_fill_2 FILLER_3_174 ();
 sg13g2_fill_2 FILLER_3_193 ();
 sg13g2_fill_1 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_fill_1 FILLER_3_224 ();
 sg13g2_fill_2 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_293 ();
 sg13g2_fill_2 FILLER_3_300 ();
 sg13g2_decap_8 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_314 ();
 sg13g2_decap_4 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_325 ();
 sg13g2_fill_1 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_fill_1 FILLER_3_355 ();
 sg13g2_fill_2 FILLER_3_370 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_fill_2 FILLER_3_405 ();
 sg13g2_fill_1 FILLER_3_433 ();
 sg13g2_fill_1 FILLER_3_439 ();
 sg13g2_fill_2 FILLER_3_445 ();
 sg13g2_fill_2 FILLER_3_451 ();
 sg13g2_fill_2 FILLER_3_458 ();
 sg13g2_fill_1 FILLER_3_490 ();
 sg13g2_fill_2 FILLER_3_525 ();
 sg13g2_fill_1 FILLER_3_527 ();
 sg13g2_fill_1 FILLER_3_532 ();
 sg13g2_fill_2 FILLER_3_537 ();
 sg13g2_fill_1 FILLER_3_539 ();
 sg13g2_fill_2 FILLER_3_566 ();
 sg13g2_fill_2 FILLER_3_615 ();
 sg13g2_fill_1 FILLER_3_657 ();
 sg13g2_fill_1 FILLER_3_662 ();
 sg13g2_fill_1 FILLER_3_689 ();
 sg13g2_fill_2 FILLER_3_711 ();
 sg13g2_fill_1 FILLER_3_723 ();
 sg13g2_fill_2 FILLER_3_745 ();
 sg13g2_decap_4 FILLER_3_811 ();
 sg13g2_fill_2 FILLER_3_818 ();
 sg13g2_fill_2 FILLER_3_851 ();
 sg13g2_fill_1 FILLER_3_853 ();
 sg13g2_fill_2 FILLER_3_884 ();
 sg13g2_fill_1 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_901 ();
 sg13g2_decap_8 FILLER_3_908 ();
 sg13g2_decap_8 FILLER_3_918 ();
 sg13g2_fill_1 FILLER_3_935 ();
 sg13g2_fill_1 FILLER_3_939 ();
 sg13g2_fill_2 FILLER_3_954 ();
 sg13g2_fill_1 FILLER_3_982 ();
 sg13g2_fill_2 FILLER_3_1009 ();
 sg13g2_fill_2 FILLER_3_1015 ();
 sg13g2_decap_4 FILLER_3_1043 ();
 sg13g2_fill_1 FILLER_3_1072 ();
 sg13g2_fill_1 FILLER_3_1094 ();
 sg13g2_fill_1 FILLER_3_1115 ();
 sg13g2_decap_8 FILLER_3_1120 ();
 sg13g2_fill_2 FILLER_3_1127 ();
 sg13g2_decap_4 FILLER_3_1137 ();
 sg13g2_fill_2 FILLER_3_1145 ();
 sg13g2_fill_2 FILLER_3_1204 ();
 sg13g2_fill_1 FILLER_3_1206 ();
 sg13g2_fill_2 FILLER_3_1267 ();
 sg13g2_fill_1 FILLER_3_1269 ();
 sg13g2_decap_4 FILLER_3_1296 ();
 sg13g2_fill_1 FILLER_3_1300 ();
 sg13g2_fill_1 FILLER_3_1305 ();
 sg13g2_decap_8 FILLER_3_1314 ();
 sg13g2_fill_2 FILLER_3_1321 ();
 sg13g2_fill_1 FILLER_3_1333 ();
 sg13g2_fill_2 FILLER_3_1348 ();
 sg13g2_decap_8 FILLER_3_1354 ();
 sg13g2_decap_8 FILLER_3_1361 ();
 sg13g2_fill_1 FILLER_3_1368 ();
 sg13g2_fill_2 FILLER_3_1492 ();
 sg13g2_fill_1 FILLER_3_1494 ();
 sg13g2_decap_8 FILLER_3_1544 ();
 sg13g2_fill_1 FILLER_3_1551 ();
 sg13g2_fill_2 FILLER_3_1593 ();
 sg13g2_fill_1 FILLER_3_1595 ();
 sg13g2_fill_1 FILLER_3_1609 ();
 sg13g2_fill_2 FILLER_3_1636 ();
 sg13g2_fill_2 FILLER_3_1644 ();
 sg13g2_fill_1 FILLER_3_1646 ();
 sg13g2_decap_4 FILLER_3_1653 ();
 sg13g2_fill_2 FILLER_3_1657 ();
 sg13g2_decap_8 FILLER_3_1671 ();
 sg13g2_decap_8 FILLER_3_1678 ();
 sg13g2_fill_1 FILLER_3_1685 ();
 sg13g2_decap_8 FILLER_3_1750 ();
 sg13g2_decap_8 FILLER_3_1757 ();
 sg13g2_fill_2 FILLER_3_1764 ();
 sg13g2_fill_2 FILLER_3_1780 ();
 sg13g2_decap_8 FILLER_3_1792 ();
 sg13g2_decap_4 FILLER_3_1799 ();
 sg13g2_decap_8 FILLER_3_1817 ();
 sg13g2_fill_1 FILLER_3_1824 ();
 sg13g2_decap_4 FILLER_3_1852 ();
 sg13g2_decap_8 FILLER_3_1881 ();
 sg13g2_fill_1 FILLER_3_1888 ();
 sg13g2_decap_8 FILLER_3_1936 ();
 sg13g2_fill_1 FILLER_3_1943 ();
 sg13g2_fill_2 FILLER_3_1983 ();
 sg13g2_decap_4 FILLER_3_2007 ();
 sg13g2_decap_8 FILLER_3_2032 ();
 sg13g2_fill_2 FILLER_3_2053 ();
 sg13g2_fill_2 FILLER_3_2059 ();
 sg13g2_fill_1 FILLER_3_2061 ();
 sg13g2_fill_2 FILLER_3_2088 ();
 sg13g2_fill_1 FILLER_3_2090 ();
 sg13g2_fill_2 FILLER_3_2101 ();
 sg13g2_fill_1 FILLER_3_2103 ();
 sg13g2_fill_2 FILLER_3_2114 ();
 sg13g2_fill_2 FILLER_3_2146 ();
 sg13g2_fill_1 FILLER_3_2148 ();
 sg13g2_decap_4 FILLER_3_2153 ();
 sg13g2_fill_2 FILLER_3_2157 ();
 sg13g2_fill_2 FILLER_3_2195 ();
 sg13g2_fill_1 FILLER_3_2197 ();
 sg13g2_fill_1 FILLER_3_2234 ();
 sg13g2_fill_2 FILLER_3_2294 ();
 sg13g2_fill_1 FILLER_3_2296 ();
 sg13g2_fill_1 FILLER_3_2323 ();
 sg13g2_fill_1 FILLER_3_2334 ();
 sg13g2_fill_1 FILLER_3_2339 ();
 sg13g2_fill_1 FILLER_3_2366 ();
 sg13g2_decap_8 FILLER_3_2411 ();
 sg13g2_decap_8 FILLER_3_2418 ();
 sg13g2_decap_8 FILLER_3_2425 ();
 sg13g2_decap_8 FILLER_3_2432 ();
 sg13g2_decap_8 FILLER_3_2439 ();
 sg13g2_decap_8 FILLER_3_2446 ();
 sg13g2_decap_8 FILLER_3_2453 ();
 sg13g2_decap_8 FILLER_3_2460 ();
 sg13g2_decap_8 FILLER_3_2467 ();
 sg13g2_decap_8 FILLER_3_2474 ();
 sg13g2_decap_8 FILLER_3_2481 ();
 sg13g2_decap_8 FILLER_3_2488 ();
 sg13g2_decap_8 FILLER_3_2495 ();
 sg13g2_decap_8 FILLER_3_2502 ();
 sg13g2_decap_8 FILLER_3_2509 ();
 sg13g2_decap_8 FILLER_3_2516 ();
 sg13g2_decap_8 FILLER_3_2523 ();
 sg13g2_decap_8 FILLER_3_2530 ();
 sg13g2_decap_8 FILLER_3_2537 ();
 sg13g2_decap_8 FILLER_3_2544 ();
 sg13g2_decap_8 FILLER_3_2551 ();
 sg13g2_decap_8 FILLER_3_2558 ();
 sg13g2_decap_8 FILLER_3_2565 ();
 sg13g2_decap_8 FILLER_3_2572 ();
 sg13g2_decap_8 FILLER_3_2579 ();
 sg13g2_decap_8 FILLER_3_2586 ();
 sg13g2_decap_8 FILLER_3_2593 ();
 sg13g2_decap_8 FILLER_3_2600 ();
 sg13g2_decap_8 FILLER_3_2607 ();
 sg13g2_decap_8 FILLER_3_2614 ();
 sg13g2_decap_8 FILLER_3_2621 ();
 sg13g2_decap_8 FILLER_3_2628 ();
 sg13g2_decap_8 FILLER_3_2635 ();
 sg13g2_decap_8 FILLER_3_2642 ();
 sg13g2_decap_8 FILLER_3_2649 ();
 sg13g2_decap_8 FILLER_3_2656 ();
 sg13g2_decap_8 FILLER_3_2663 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_fill_2 FILLER_4_39 ();
 sg13g2_fill_1 FILLER_4_72 ();
 sg13g2_fill_1 FILLER_4_77 ();
 sg13g2_fill_1 FILLER_4_82 ();
 sg13g2_decap_4 FILLER_4_88 ();
 sg13g2_fill_2 FILLER_4_92 ();
 sg13g2_decap_4 FILLER_4_104 ();
 sg13g2_fill_1 FILLER_4_108 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_150 ();
 sg13g2_fill_2 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_202 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_decap_4 FILLER_4_249 ();
 sg13g2_fill_2 FILLER_4_253 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_290 ();
 sg13g2_fill_1 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_fill_2 FILLER_4_325 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_decap_4 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_fill_2 FILLER_4_397 ();
 sg13g2_decap_8 FILLER_4_407 ();
 sg13g2_decap_4 FILLER_4_418 ();
 sg13g2_fill_2 FILLER_4_482 ();
 sg13g2_fill_1 FILLER_4_489 ();
 sg13g2_decap_8 FILLER_4_509 ();
 sg13g2_decap_8 FILLER_4_516 ();
 sg13g2_decap_8 FILLER_4_523 ();
 sg13g2_fill_2 FILLER_4_530 ();
 sg13g2_fill_1 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_555 ();
 sg13g2_fill_1 FILLER_4_562 ();
 sg13g2_decap_4 FILLER_4_571 ();
 sg13g2_fill_1 FILLER_4_575 ();
 sg13g2_fill_1 FILLER_4_613 ();
 sg13g2_fill_2 FILLER_4_628 ();
 sg13g2_fill_2 FILLER_4_634 ();
 sg13g2_fill_2 FILLER_4_662 ();
 sg13g2_fill_1 FILLER_4_664 ();
 sg13g2_fill_1 FILLER_4_691 ();
 sg13g2_fill_2 FILLER_4_718 ();
 sg13g2_fill_1 FILLER_4_720 ();
 sg13g2_decap_4 FILLER_4_725 ();
 sg13g2_fill_2 FILLER_4_729 ();
 sg13g2_fill_1 FILLER_4_768 ();
 sg13g2_decap_8 FILLER_4_773 ();
 sg13g2_decap_4 FILLER_4_780 ();
 sg13g2_fill_1 FILLER_4_784 ();
 sg13g2_decap_4 FILLER_4_811 ();
 sg13g2_fill_1 FILLER_4_836 ();
 sg13g2_decap_4 FILLER_4_841 ();
 sg13g2_decap_4 FILLER_4_885 ();
 sg13g2_fill_1 FILLER_4_889 ();
 sg13g2_decap_4 FILLER_4_900 ();
 sg13g2_fill_2 FILLER_4_908 ();
 sg13g2_fill_1 FILLER_4_914 ();
 sg13g2_fill_1 FILLER_4_974 ();
 sg13g2_fill_2 FILLER_4_985 ();
 sg13g2_fill_1 FILLER_4_987 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_fill_2 FILLER_4_1025 ();
 sg13g2_decap_4 FILLER_4_1037 ();
 sg13g2_fill_2 FILLER_4_1041 ();
 sg13g2_decap_8 FILLER_4_1047 ();
 sg13g2_decap_8 FILLER_4_1054 ();
 sg13g2_decap_8 FILLER_4_1061 ();
 sg13g2_fill_2 FILLER_4_1068 ();
 sg13g2_fill_2 FILLER_4_1091 ();
 sg13g2_fill_1 FILLER_4_1093 ();
 sg13g2_fill_1 FILLER_4_1102 ();
 sg13g2_fill_2 FILLER_4_1107 ();
 sg13g2_fill_2 FILLER_4_1119 ();
 sg13g2_fill_1 FILLER_4_1121 ();
 sg13g2_decap_8 FILLER_4_1152 ();
 sg13g2_fill_1 FILLER_4_1163 ();
 sg13g2_fill_2 FILLER_4_1168 ();
 sg13g2_fill_2 FILLER_4_1178 ();
 sg13g2_decap_8 FILLER_4_1184 ();
 sg13g2_decap_8 FILLER_4_1191 ();
 sg13g2_decap_8 FILLER_4_1198 ();
 sg13g2_decap_4 FILLER_4_1205 ();
 sg13g2_fill_1 FILLER_4_1213 ();
 sg13g2_fill_2 FILLER_4_1218 ();
 sg13g2_fill_2 FILLER_4_1224 ();
 sg13g2_fill_2 FILLER_4_1230 ();
 sg13g2_fill_2 FILLER_4_1236 ();
 sg13g2_fill_2 FILLER_4_1310 ();
 sg13g2_decap_8 FILLER_4_1322 ();
 sg13g2_decap_4 FILLER_4_1339 ();
 sg13g2_decap_8 FILLER_4_1347 ();
 sg13g2_decap_8 FILLER_4_1354 ();
 sg13g2_fill_2 FILLER_4_1361 ();
 sg13g2_decap_4 FILLER_4_1418 ();
 sg13g2_fill_1 FILLER_4_1422 ();
 sg13g2_decap_8 FILLER_4_1433 ();
 sg13g2_decap_8 FILLER_4_1440 ();
 sg13g2_fill_2 FILLER_4_1447 ();
 sg13g2_fill_2 FILLER_4_1459 ();
 sg13g2_fill_1 FILLER_4_1461 ();
 sg13g2_decap_4 FILLER_4_1466 ();
 sg13g2_fill_1 FILLER_4_1470 ();
 sg13g2_fill_1 FILLER_4_1511 ();
 sg13g2_fill_2 FILLER_4_1522 ();
 sg13g2_fill_1 FILLER_4_1524 ();
 sg13g2_fill_1 FILLER_4_1535 ();
 sg13g2_decap_8 FILLER_4_1540 ();
 sg13g2_decap_8 FILLER_4_1547 ();
 sg13g2_decap_4 FILLER_4_1554 ();
 sg13g2_fill_2 FILLER_4_1558 ();
 sg13g2_fill_2 FILLER_4_1596 ();
 sg13g2_decap_8 FILLER_4_1620 ();
 sg13g2_decap_4 FILLER_4_1627 ();
 sg13g2_fill_1 FILLER_4_1631 ();
 sg13g2_decap_8 FILLER_4_1637 ();
 sg13g2_fill_2 FILLER_4_1644 ();
 sg13g2_fill_1 FILLER_4_1646 ();
 sg13g2_fill_1 FILLER_4_1652 ();
 sg13g2_decap_4 FILLER_4_1658 ();
 sg13g2_fill_1 FILLER_4_1662 ();
 sg13g2_fill_2 FILLER_4_1668 ();
 sg13g2_fill_1 FILLER_4_1670 ();
 sg13g2_decap_8 FILLER_4_1675 ();
 sg13g2_fill_2 FILLER_4_1687 ();
 sg13g2_fill_1 FILLER_4_1689 ();
 sg13g2_decap_4 FILLER_4_1696 ();
 sg13g2_fill_2 FILLER_4_1718 ();
 sg13g2_fill_1 FILLER_4_1720 ();
 sg13g2_fill_2 FILLER_4_1727 ();
 sg13g2_decap_8 FILLER_4_1755 ();
 sg13g2_decap_8 FILLER_4_1762 ();
 sg13g2_decap_8 FILLER_4_1769 ();
 sg13g2_decap_8 FILLER_4_1776 ();
 sg13g2_fill_2 FILLER_4_1783 ();
 sg13g2_decap_8 FILLER_4_1817 ();
 sg13g2_decap_8 FILLER_4_1824 ();
 sg13g2_decap_8 FILLER_4_1831 ();
 sg13g2_decap_8 FILLER_4_1838 ();
 sg13g2_fill_1 FILLER_4_1845 ();
 sg13g2_fill_2 FILLER_4_1856 ();
 sg13g2_decap_8 FILLER_4_1868 ();
 sg13g2_decap_8 FILLER_4_1875 ();
 sg13g2_decap_8 FILLER_4_1882 ();
 sg13g2_decap_8 FILLER_4_1889 ();
 sg13g2_fill_2 FILLER_4_1896 ();
 sg13g2_decap_8 FILLER_4_1902 ();
 sg13g2_decap_8 FILLER_4_1909 ();
 sg13g2_decap_4 FILLER_4_1937 ();
 sg13g2_fill_1 FILLER_4_1945 ();
 sg13g2_fill_1 FILLER_4_1966 ();
 sg13g2_fill_1 FILLER_4_1971 ();
 sg13g2_fill_1 FILLER_4_1998 ();
 sg13g2_fill_1 FILLER_4_2009 ();
 sg13g2_decap_8 FILLER_4_2036 ();
 sg13g2_fill_2 FILLER_4_2043 ();
 sg13g2_fill_2 FILLER_4_2102 ();
 sg13g2_fill_1 FILLER_4_2104 ();
 sg13g2_fill_1 FILLER_4_2128 ();
 sg13g2_decap_8 FILLER_4_2146 ();
 sg13g2_decap_8 FILLER_4_2153 ();
 sg13g2_fill_2 FILLER_4_2160 ();
 sg13g2_fill_1 FILLER_4_2162 ();
 sg13g2_fill_2 FILLER_4_2173 ();
 sg13g2_decap_8 FILLER_4_2179 ();
 sg13g2_decap_8 FILLER_4_2186 ();
 sg13g2_decap_8 FILLER_4_2193 ();
 sg13g2_decap_4 FILLER_4_2200 ();
 sg13g2_fill_2 FILLER_4_2208 ();
 sg13g2_decap_8 FILLER_4_2235 ();
 sg13g2_fill_2 FILLER_4_2242 ();
 sg13g2_fill_1 FILLER_4_2244 ();
 sg13g2_decap_4 FILLER_4_2255 ();
 sg13g2_fill_2 FILLER_4_2263 ();
 sg13g2_fill_2 FILLER_4_2268 ();
 sg13g2_fill_1 FILLER_4_2270 ();
 sg13g2_decap_8 FILLER_4_2275 ();
 sg13g2_decap_4 FILLER_4_2282 ();
 sg13g2_fill_2 FILLER_4_2286 ();
 sg13g2_fill_2 FILLER_4_2309 ();
 sg13g2_decap_8 FILLER_4_2315 ();
 sg13g2_decap_4 FILLER_4_2322 ();
 sg13g2_fill_1 FILLER_4_2326 ();
 sg13g2_decap_8 FILLER_4_2413 ();
 sg13g2_decap_8 FILLER_4_2420 ();
 sg13g2_decap_8 FILLER_4_2427 ();
 sg13g2_decap_8 FILLER_4_2434 ();
 sg13g2_decap_8 FILLER_4_2441 ();
 sg13g2_decap_8 FILLER_4_2448 ();
 sg13g2_decap_8 FILLER_4_2455 ();
 sg13g2_decap_8 FILLER_4_2462 ();
 sg13g2_decap_8 FILLER_4_2469 ();
 sg13g2_decap_8 FILLER_4_2476 ();
 sg13g2_decap_8 FILLER_4_2483 ();
 sg13g2_decap_8 FILLER_4_2490 ();
 sg13g2_decap_8 FILLER_4_2497 ();
 sg13g2_decap_8 FILLER_4_2504 ();
 sg13g2_decap_8 FILLER_4_2511 ();
 sg13g2_decap_8 FILLER_4_2518 ();
 sg13g2_decap_8 FILLER_4_2525 ();
 sg13g2_decap_8 FILLER_4_2532 ();
 sg13g2_decap_8 FILLER_4_2539 ();
 sg13g2_decap_8 FILLER_4_2546 ();
 sg13g2_decap_8 FILLER_4_2553 ();
 sg13g2_decap_8 FILLER_4_2560 ();
 sg13g2_decap_8 FILLER_4_2567 ();
 sg13g2_decap_8 FILLER_4_2574 ();
 sg13g2_decap_8 FILLER_4_2581 ();
 sg13g2_decap_8 FILLER_4_2588 ();
 sg13g2_decap_8 FILLER_4_2595 ();
 sg13g2_decap_8 FILLER_4_2602 ();
 sg13g2_decap_8 FILLER_4_2609 ();
 sg13g2_decap_8 FILLER_4_2616 ();
 sg13g2_decap_8 FILLER_4_2623 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_8 FILLER_4_2644 ();
 sg13g2_decap_8 FILLER_4_2651 ();
 sg13g2_decap_8 FILLER_4_2658 ();
 sg13g2_decap_4 FILLER_4_2665 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_13 ();
 sg13g2_fill_1 FILLER_5_52 ();
 sg13g2_fill_2 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_fill_2 FILLER_5_100 ();
 sg13g2_fill_1 FILLER_5_143 ();
 sg13g2_fill_1 FILLER_5_170 ();
 sg13g2_decap_8 FILLER_5_211 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_decap_4 FILLER_5_246 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_2 FILLER_5_278 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_fill_2 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_288 ();
 sg13g2_fill_1 FILLER_5_299 ();
 sg13g2_fill_2 FILLER_5_330 ();
 sg13g2_fill_2 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_4 FILLER_5_393 ();
 sg13g2_fill_2 FILLER_5_397 ();
 sg13g2_fill_1 FILLER_5_403 ();
 sg13g2_decap_4 FILLER_5_413 ();
 sg13g2_fill_2 FILLER_5_417 ();
 sg13g2_fill_1 FILLER_5_432 ();
 sg13g2_decap_4 FILLER_5_516 ();
 sg13g2_fill_1 FILLER_5_520 ();
 sg13g2_fill_2 FILLER_5_563 ();
 sg13g2_decap_8 FILLER_5_569 ();
 sg13g2_decap_8 FILLER_5_576 ();
 sg13g2_fill_1 FILLER_5_583 ();
 sg13g2_fill_1 FILLER_5_590 ();
 sg13g2_fill_1 FILLER_5_603 ();
 sg13g2_decap_4 FILLER_5_640 ();
 sg13g2_fill_1 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_649 ();
 sg13g2_decap_8 FILLER_5_656 ();
 sg13g2_fill_2 FILLER_5_663 ();
 sg13g2_decap_4 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_fill_2 FILLER_5_704 ();
 sg13g2_fill_1 FILLER_5_706 ();
 sg13g2_decap_8 FILLER_5_717 ();
 sg13g2_fill_1 FILLER_5_764 ();
 sg13g2_decap_8 FILLER_5_775 ();
 sg13g2_decap_8 FILLER_5_782 ();
 sg13g2_fill_2 FILLER_5_789 ();
 sg13g2_decap_4 FILLER_5_821 ();
 sg13g2_fill_2 FILLER_5_825 ();
 sg13g2_fill_1 FILLER_5_853 ();
 sg13g2_fill_1 FILLER_5_864 ();
 sg13g2_fill_1 FILLER_5_869 ();
 sg13g2_decap_4 FILLER_5_896 ();
 sg13g2_fill_2 FILLER_5_936 ();
 sg13g2_decap_8 FILLER_5_941 ();
 sg13g2_decap_8 FILLER_5_969 ();
 sg13g2_decap_8 FILLER_5_976 ();
 sg13g2_decap_4 FILLER_5_983 ();
 sg13g2_fill_1 FILLER_5_987 ();
 sg13g2_decap_8 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1013 ();
 sg13g2_decap_4 FILLER_5_1020 ();
 sg13g2_fill_2 FILLER_5_1024 ();
 sg13g2_decap_8 FILLER_5_1062 ();
 sg13g2_decap_8 FILLER_5_1069 ();
 sg13g2_decap_4 FILLER_5_1076 ();
 sg13g2_fill_1 FILLER_5_1090 ();
 sg13g2_decap_4 FILLER_5_1168 ();
 sg13g2_fill_1 FILLER_5_1172 ();
 sg13g2_fill_1 FILLER_5_1177 ();
 sg13g2_fill_1 FILLER_5_1183 ();
 sg13g2_fill_2 FILLER_5_1214 ();
 sg13g2_fill_1 FILLER_5_1216 ();
 sg13g2_decap_4 FILLER_5_1247 ();
 sg13g2_fill_1 FILLER_5_1251 ();
 sg13g2_fill_1 FILLER_5_1269 ();
 sg13g2_decap_4 FILLER_5_1304 ();
 sg13g2_fill_2 FILLER_5_1308 ();
 sg13g2_fill_2 FILLER_5_1362 ();
 sg13g2_fill_1 FILLER_5_1364 ();
 sg13g2_decap_8 FILLER_5_1395 ();
 sg13g2_decap_8 FILLER_5_1424 ();
 sg13g2_decap_8 FILLER_5_1431 ();
 sg13g2_decap_8 FILLER_5_1438 ();
 sg13g2_decap_8 FILLER_5_1445 ();
 sg13g2_decap_4 FILLER_5_1452 ();
 sg13g2_fill_1 FILLER_5_1456 ();
 sg13g2_fill_2 FILLER_5_1467 ();
 sg13g2_decap_4 FILLER_5_1490 ();
 sg13g2_fill_1 FILLER_5_1494 ();
 sg13g2_decap_8 FILLER_5_1535 ();
 sg13g2_decap_8 FILLER_5_1542 ();
 sg13g2_decap_8 FILLER_5_1549 ();
 sg13g2_decap_8 FILLER_5_1556 ();
 sg13g2_fill_2 FILLER_5_1563 ();
 sg13g2_fill_1 FILLER_5_1565 ();
 sg13g2_decap_4 FILLER_5_1574 ();
 sg13g2_decap_8 FILLER_5_1629 ();
 sg13g2_fill_2 FILLER_5_1636 ();
 sg13g2_fill_1 FILLER_5_1638 ();
 sg13g2_fill_2 FILLER_5_1644 ();
 sg13g2_fill_1 FILLER_5_1651 ();
 sg13g2_fill_2 FILLER_5_1662 ();
 sg13g2_fill_1 FILLER_5_1695 ();
 sg13g2_fill_2 FILLER_5_1700 ();
 sg13g2_decap_8 FILLER_5_1751 ();
 sg13g2_fill_1 FILLER_5_1762 ();
 sg13g2_decap_4 FILLER_5_1776 ();
 sg13g2_fill_1 FILLER_5_1794 ();
 sg13g2_decap_4 FILLER_5_1821 ();
 sg13g2_fill_2 FILLER_5_1825 ();
 sg13g2_decap_8 FILLER_5_1889 ();
 sg13g2_decap_4 FILLER_5_1896 ();
 sg13g2_fill_1 FILLER_5_1900 ();
 sg13g2_fill_2 FILLER_5_1911 ();
 sg13g2_fill_1 FILLER_5_1913 ();
 sg13g2_decap_4 FILLER_5_1940 ();
 sg13g2_fill_2 FILLER_5_1944 ();
 sg13g2_fill_1 FILLER_5_1956 ();
 sg13g2_fill_1 FILLER_5_1961 ();
 sg13g2_fill_2 FILLER_5_1966 ();
 sg13g2_fill_1 FILLER_5_1968 ();
 sg13g2_decap_4 FILLER_5_1973 ();
 sg13g2_fill_2 FILLER_5_1977 ();
 sg13g2_decap_8 FILLER_5_1987 ();
 sg13g2_decap_4 FILLER_5_1994 ();
 sg13g2_fill_1 FILLER_5_1998 ();
 sg13g2_fill_2 FILLER_5_2007 ();
 sg13g2_fill_1 FILLER_5_2009 ();
 sg13g2_fill_1 FILLER_5_2032 ();
 sg13g2_decap_4 FILLER_5_2037 ();
 sg13g2_fill_2 FILLER_5_2041 ();
 sg13g2_decap_8 FILLER_5_2108 ();
 sg13g2_fill_2 FILLER_5_2115 ();
 sg13g2_decap_8 FILLER_5_2127 ();
 sg13g2_decap_4 FILLER_5_2134 ();
 sg13g2_fill_1 FILLER_5_2138 ();
 sg13g2_fill_2 FILLER_5_2165 ();
 sg13g2_decap_4 FILLER_5_2171 ();
 sg13g2_fill_1 FILLER_5_2175 ();
 sg13g2_fill_2 FILLER_5_2216 ();
 sg13g2_fill_1 FILLER_5_2218 ();
 sg13g2_decap_8 FILLER_5_2229 ();
 sg13g2_fill_2 FILLER_5_2236 ();
 sg13g2_fill_1 FILLER_5_2238 ();
 sg13g2_decap_8 FILLER_5_2284 ();
 sg13g2_fill_1 FILLER_5_2291 ();
 sg13g2_decap_4 FILLER_5_2296 ();
 sg13g2_decap_8 FILLER_5_2327 ();
 sg13g2_decap_8 FILLER_5_2334 ();
 sg13g2_decap_4 FILLER_5_2341 ();
 sg13g2_decap_8 FILLER_5_2366 ();
 sg13g2_decap_8 FILLER_5_2373 ();
 sg13g2_decap_8 FILLER_5_2393 ();
 sg13g2_decap_8 FILLER_5_2400 ();
 sg13g2_decap_8 FILLER_5_2407 ();
 sg13g2_decap_8 FILLER_5_2414 ();
 sg13g2_decap_8 FILLER_5_2421 ();
 sg13g2_decap_8 FILLER_5_2428 ();
 sg13g2_decap_8 FILLER_5_2435 ();
 sg13g2_decap_8 FILLER_5_2442 ();
 sg13g2_decap_8 FILLER_5_2449 ();
 sg13g2_decap_8 FILLER_5_2456 ();
 sg13g2_decap_8 FILLER_5_2463 ();
 sg13g2_decap_8 FILLER_5_2470 ();
 sg13g2_decap_8 FILLER_5_2477 ();
 sg13g2_decap_8 FILLER_5_2484 ();
 sg13g2_decap_8 FILLER_5_2491 ();
 sg13g2_decap_8 FILLER_5_2498 ();
 sg13g2_decap_8 FILLER_5_2505 ();
 sg13g2_decap_8 FILLER_5_2512 ();
 sg13g2_decap_8 FILLER_5_2519 ();
 sg13g2_decap_8 FILLER_5_2526 ();
 sg13g2_decap_8 FILLER_5_2533 ();
 sg13g2_decap_8 FILLER_5_2540 ();
 sg13g2_decap_8 FILLER_5_2547 ();
 sg13g2_decap_8 FILLER_5_2554 ();
 sg13g2_decap_8 FILLER_5_2561 ();
 sg13g2_decap_8 FILLER_5_2568 ();
 sg13g2_decap_8 FILLER_5_2575 ();
 sg13g2_decap_8 FILLER_5_2582 ();
 sg13g2_decap_8 FILLER_5_2589 ();
 sg13g2_decap_8 FILLER_5_2596 ();
 sg13g2_decap_8 FILLER_5_2603 ();
 sg13g2_decap_8 FILLER_5_2610 ();
 sg13g2_decap_8 FILLER_5_2617 ();
 sg13g2_decap_8 FILLER_5_2624 ();
 sg13g2_decap_8 FILLER_5_2631 ();
 sg13g2_decap_8 FILLER_5_2638 ();
 sg13g2_decap_8 FILLER_5_2645 ();
 sg13g2_decap_8 FILLER_5_2652 ();
 sg13g2_decap_8 FILLER_5_2659 ();
 sg13g2_decap_4 FILLER_5_2666 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_12 ();
 sg13g2_fill_2 FILLER_6_44 ();
 sg13g2_fill_1 FILLER_6_50 ();
 sg13g2_fill_2 FILLER_6_89 ();
 sg13g2_decap_4 FILLER_6_95 ();
 sg13g2_fill_2 FILLER_6_170 ();
 sg13g2_fill_1 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_4 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_246 ();
 sg13g2_fill_2 FILLER_6_296 ();
 sg13g2_fill_2 FILLER_6_307 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_2 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_fill_2 FILLER_6_390 ();
 sg13g2_fill_1 FILLER_6_392 ();
 sg13g2_fill_2 FILLER_6_397 ();
 sg13g2_fill_2 FILLER_6_403 ();
 sg13g2_fill_1 FILLER_6_405 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_439 ();
 sg13g2_fill_2 FILLER_6_451 ();
 sg13g2_fill_1 FILLER_6_471 ();
 sg13g2_fill_1 FILLER_6_477 ();
 sg13g2_fill_1 FILLER_6_495 ();
 sg13g2_fill_2 FILLER_6_512 ();
 sg13g2_fill_1 FILLER_6_546 ();
 sg13g2_fill_1 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_fill_2 FILLER_6_722 ();
 sg13g2_fill_2 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_fill_1 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_790 ();
 sg13g2_decap_4 FILLER_6_797 ();
 sg13g2_fill_2 FILLER_6_809 ();
 sg13g2_fill_1 FILLER_6_811 ();
 sg13g2_decap_4 FILLER_6_822 ();
 sg13g2_fill_1 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_8 FILLER_6_858 ();
 sg13g2_fill_2 FILLER_6_865 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_fill_1 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_959 ();
 sg13g2_decap_8 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_decap_8 FILLER_6_987 ();
 sg13g2_decap_8 FILLER_6_994 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_decap_8 FILLER_6_1008 ();
 sg13g2_decap_8 FILLER_6_1015 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1029 ();
 sg13g2_fill_2 FILLER_6_1036 ();
 sg13g2_fill_1 FILLER_6_1038 ();
 sg13g2_decap_8 FILLER_6_1065 ();
 sg13g2_decap_8 FILLER_6_1072 ();
 sg13g2_fill_1 FILLER_6_1079 ();
 sg13g2_fill_2 FILLER_6_1132 ();
 sg13g2_fill_1 FILLER_6_1160 ();
 sg13g2_fill_2 FILLER_6_1166 ();
 sg13g2_fill_2 FILLER_6_1194 ();
 sg13g2_fill_1 FILLER_6_1196 ();
 sg13g2_fill_2 FILLER_6_1202 ();
 sg13g2_fill_1 FILLER_6_1239 ();
 sg13g2_fill_2 FILLER_6_1283 ();
 sg13g2_decap_4 FILLER_6_1294 ();
 sg13g2_fill_1 FILLER_6_1298 ();
 sg13g2_fill_1 FILLER_6_1311 ();
 sg13g2_fill_1 FILLER_6_1316 ();
 sg13g2_fill_2 FILLER_6_1321 ();
 sg13g2_fill_1 FILLER_6_1323 ();
 sg13g2_decap_4 FILLER_6_1355 ();
 sg13g2_fill_1 FILLER_6_1359 ();
 sg13g2_decap_8 FILLER_6_1368 ();
 sg13g2_decap_8 FILLER_6_1375 ();
 sg13g2_fill_2 FILLER_6_1386 ();
 sg13g2_fill_2 FILLER_6_1409 ();
 sg13g2_fill_1 FILLER_6_1415 ();
 sg13g2_fill_1 FILLER_6_1420 ();
 sg13g2_fill_2 FILLER_6_1447 ();
 sg13g2_decap_8 FILLER_6_1483 ();
 sg13g2_decap_4 FILLER_6_1490 ();
 sg13g2_decap_8 FILLER_6_1533 ();
 sg13g2_decap_4 FILLER_6_1540 ();
 sg13g2_fill_1 FILLER_6_1544 ();
 sg13g2_decap_4 FILLER_6_1581 ();
 sg13g2_fill_1 FILLER_6_1585 ();
 sg13g2_fill_1 FILLER_6_1595 ();
 sg13g2_fill_2 FILLER_6_1601 ();
 sg13g2_fill_1 FILLER_6_1603 ();
 sg13g2_fill_2 FILLER_6_1639 ();
 sg13g2_fill_1 FILLER_6_1641 ();
 sg13g2_decap_4 FILLER_6_1647 ();
 sg13g2_fill_1 FILLER_6_1651 ();
 sg13g2_fill_2 FILLER_6_1657 ();
 sg13g2_fill_2 FILLER_6_1669 ();
 sg13g2_fill_1 FILLER_6_1671 ();
 sg13g2_fill_1 FILLER_6_1698 ();
 sg13g2_fill_1 FILLER_6_1703 ();
 sg13g2_fill_2 FILLER_6_1720 ();
 sg13g2_fill_1 FILLER_6_1722 ();
 sg13g2_fill_2 FILLER_6_1757 ();
 sg13g2_fill_2 FILLER_6_1764 ();
 sg13g2_fill_2 FILLER_6_1792 ();
 sg13g2_fill_2 FILLER_6_1825 ();
 sg13g2_fill_2 FILLER_6_1863 ();
 sg13g2_fill_1 FILLER_6_1865 ();
 sg13g2_fill_2 FILLER_6_1870 ();
 sg13g2_fill_1 FILLER_6_1872 ();
 sg13g2_decap_4 FILLER_6_1975 ();
 sg13g2_fill_2 FILLER_6_1979 ();
 sg13g2_fill_1 FILLER_6_2022 ();
 sg13g2_fill_2 FILLER_6_2078 ();
 sg13g2_fill_2 FILLER_6_2130 ();
 sg13g2_fill_1 FILLER_6_2132 ();
 sg13g2_fill_2 FILLER_6_2137 ();
 sg13g2_fill_2 FILLER_6_2160 ();
 sg13g2_fill_1 FILLER_6_2162 ();
 sg13g2_decap_8 FILLER_6_2167 ();
 sg13g2_fill_2 FILLER_6_2174 ();
 sg13g2_fill_2 FILLER_6_2185 ();
 sg13g2_fill_1 FILLER_6_2221 ();
 sg13g2_fill_1 FILLER_6_2264 ();
 sg13g2_fill_2 FILLER_6_2269 ();
 sg13g2_fill_2 FILLER_6_2274 ();
 sg13g2_fill_2 FILLER_6_2338 ();
 sg13g2_fill_2 FILLER_6_2350 ();
 sg13g2_fill_2 FILLER_6_2356 ();
 sg13g2_fill_1 FILLER_6_2358 ();
 sg13g2_fill_2 FILLER_6_2385 ();
 sg13g2_fill_1 FILLER_6_2387 ();
 sg13g2_fill_2 FILLER_6_2398 ();
 sg13g2_decap_4 FILLER_6_2410 ();
 sg13g2_decap_8 FILLER_6_2418 ();
 sg13g2_decap_8 FILLER_6_2425 ();
 sg13g2_decap_8 FILLER_6_2432 ();
 sg13g2_decap_8 FILLER_6_2439 ();
 sg13g2_decap_8 FILLER_6_2446 ();
 sg13g2_decap_8 FILLER_6_2453 ();
 sg13g2_decap_8 FILLER_6_2460 ();
 sg13g2_decap_8 FILLER_6_2467 ();
 sg13g2_decap_8 FILLER_6_2474 ();
 sg13g2_decap_8 FILLER_6_2481 ();
 sg13g2_decap_8 FILLER_6_2488 ();
 sg13g2_decap_8 FILLER_6_2495 ();
 sg13g2_decap_8 FILLER_6_2502 ();
 sg13g2_decap_8 FILLER_6_2509 ();
 sg13g2_decap_8 FILLER_6_2516 ();
 sg13g2_decap_8 FILLER_6_2523 ();
 sg13g2_decap_8 FILLER_6_2530 ();
 sg13g2_decap_8 FILLER_6_2537 ();
 sg13g2_decap_8 FILLER_6_2544 ();
 sg13g2_decap_8 FILLER_6_2551 ();
 sg13g2_decap_8 FILLER_6_2558 ();
 sg13g2_decap_8 FILLER_6_2565 ();
 sg13g2_decap_8 FILLER_6_2572 ();
 sg13g2_decap_8 FILLER_6_2579 ();
 sg13g2_decap_8 FILLER_6_2586 ();
 sg13g2_decap_8 FILLER_6_2593 ();
 sg13g2_decap_8 FILLER_6_2600 ();
 sg13g2_decap_8 FILLER_6_2607 ();
 sg13g2_decap_8 FILLER_6_2614 ();
 sg13g2_decap_8 FILLER_6_2621 ();
 sg13g2_decap_8 FILLER_6_2628 ();
 sg13g2_decap_8 FILLER_6_2635 ();
 sg13g2_decap_8 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2656 ();
 sg13g2_decap_8 FILLER_6_2663 ();
 sg13g2_fill_1 FILLER_7_32 ();
 sg13g2_fill_1 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_45 ();
 sg13g2_fill_1 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_66 ();
 sg13g2_fill_1 FILLER_7_93 ();
 sg13g2_fill_1 FILLER_7_99 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_fill_2 FILLER_7_191 ();
 sg13g2_fill_1 FILLER_7_243 ();
 sg13g2_fill_2 FILLER_7_254 ();
 sg13g2_fill_2 FILLER_7_260 ();
 sg13g2_fill_1 FILLER_7_262 ();
 sg13g2_fill_2 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_decap_4 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_285 ();
 sg13g2_decap_4 FILLER_7_296 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_7_355 ();
 sg13g2_fill_1 FILLER_7_416 ();
 sg13g2_fill_1 FILLER_7_437 ();
 sg13g2_fill_2 FILLER_7_442 ();
 sg13g2_fill_2 FILLER_7_467 ();
 sg13g2_fill_2 FILLER_7_474 ();
 sg13g2_fill_1 FILLER_7_496 ();
 sg13g2_fill_2 FILLER_7_505 ();
 sg13g2_fill_1 FILLER_7_507 ();
 sg13g2_fill_2 FILLER_7_522 ();
 sg13g2_fill_1 FILLER_7_524 ();
 sg13g2_decap_4 FILLER_7_537 ();
 sg13g2_decap_8 FILLER_7_547 ();
 sg13g2_fill_2 FILLER_7_554 ();
 sg13g2_decap_4 FILLER_7_561 ();
 sg13g2_decap_4 FILLER_7_571 ();
 sg13g2_decap_8 FILLER_7_624 ();
 sg13g2_fill_2 FILLER_7_631 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_fill_2 FILLER_7_686 ();
 sg13g2_fill_2 FILLER_7_706 ();
 sg13g2_fill_1 FILLER_7_708 ();
 sg13g2_decap_4 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_fill_2 FILLER_7_791 ();
 sg13g2_decap_4 FILLER_7_850 ();
 sg13g2_fill_2 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_887 ();
 sg13g2_fill_1 FILLER_7_894 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_4 FILLER_7_910 ();
 sg13g2_fill_2 FILLER_7_967 ();
 sg13g2_fill_1 FILLER_7_969 ();
 sg13g2_fill_2 FILLER_7_996 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_fill_1 FILLER_7_1039 ();
 sg13g2_fill_2 FILLER_7_1044 ();
 sg13g2_fill_2 FILLER_7_1085 ();
 sg13g2_fill_1 FILLER_7_1087 ();
 sg13g2_fill_2 FILLER_7_1114 ();
 sg13g2_fill_1 FILLER_7_1116 ();
 sg13g2_fill_1 FILLER_7_1164 ();
 sg13g2_fill_2 FILLER_7_1170 ();
 sg13g2_fill_1 FILLER_7_1172 ();
 sg13g2_fill_1 FILLER_7_1178 ();
 sg13g2_fill_1 FILLER_7_1225 ();
 sg13g2_fill_2 FILLER_7_1230 ();
 sg13g2_fill_2 FILLER_7_1237 ();
 sg13g2_fill_1 FILLER_7_1239 ();
 sg13g2_decap_4 FILLER_7_1266 ();
 sg13g2_fill_2 FILLER_7_1275 ();
 sg13g2_fill_1 FILLER_7_1277 ();
 sg13g2_fill_1 FILLER_7_1282 ();
 sg13g2_fill_2 FILLER_7_1304 ();
 sg13g2_fill_2 FILLER_7_1310 ();
 sg13g2_fill_1 FILLER_7_1312 ();
 sg13g2_fill_1 FILLER_7_1365 ();
 sg13g2_fill_2 FILLER_7_1428 ();
 sg13g2_fill_1 FILLER_7_1430 ();
 sg13g2_decap_8 FILLER_7_1441 ();
 sg13g2_fill_2 FILLER_7_1448 ();
 sg13g2_fill_1 FILLER_7_1512 ();
 sg13g2_fill_2 FILLER_7_1517 ();
 sg13g2_fill_1 FILLER_7_1545 ();
 sg13g2_decap_4 FILLER_7_1587 ();
 sg13g2_fill_2 FILLER_7_1591 ();
 sg13g2_fill_2 FILLER_7_1649 ();
 sg13g2_fill_2 FILLER_7_1656 ();
 sg13g2_fill_1 FILLER_7_1658 ();
 sg13g2_fill_1 FILLER_7_1663 ();
 sg13g2_fill_2 FILLER_7_1669 ();
 sg13g2_fill_1 FILLER_7_1675 ();
 sg13g2_fill_1 FILLER_7_1686 ();
 sg13g2_fill_1 FILLER_7_1696 ();
 sg13g2_decap_4 FILLER_7_1763 ();
 sg13g2_fill_2 FILLER_7_1767 ();
 sg13g2_decap_4 FILLER_7_1777 ();
 sg13g2_fill_1 FILLER_7_1781 ();
 sg13g2_fill_1 FILLER_7_1786 ();
 sg13g2_decap_8 FILLER_7_1797 ();
 sg13g2_fill_1 FILLER_7_1804 ();
 sg13g2_fill_1 FILLER_7_1815 ();
 sg13g2_fill_2 FILLER_7_1823 ();
 sg13g2_fill_2 FILLER_7_1872 ();
 sg13g2_fill_2 FILLER_7_1885 ();
 sg13g2_fill_1 FILLER_7_1913 ();
 sg13g2_fill_2 FILLER_7_1975 ();
 sg13g2_decap_8 FILLER_7_1987 ();
 sg13g2_fill_1 FILLER_7_2020 ();
 sg13g2_decap_4 FILLER_7_2057 ();
 sg13g2_fill_2 FILLER_7_2097 ();
 sg13g2_fill_1 FILLER_7_2099 ();
 sg13g2_decap_8 FILLER_7_2230 ();
 sg13g2_fill_2 FILLER_7_2263 ();
 sg13g2_fill_2 FILLER_7_2399 ();
 sg13g2_fill_1 FILLER_7_2427 ();
 sg13g2_decap_8 FILLER_7_2432 ();
 sg13g2_decap_8 FILLER_7_2439 ();
 sg13g2_decap_8 FILLER_7_2446 ();
 sg13g2_decap_8 FILLER_7_2453 ();
 sg13g2_decap_8 FILLER_7_2460 ();
 sg13g2_decap_8 FILLER_7_2467 ();
 sg13g2_decap_8 FILLER_7_2474 ();
 sg13g2_decap_8 FILLER_7_2481 ();
 sg13g2_decap_8 FILLER_7_2488 ();
 sg13g2_decap_8 FILLER_7_2495 ();
 sg13g2_decap_8 FILLER_7_2502 ();
 sg13g2_decap_8 FILLER_7_2509 ();
 sg13g2_decap_8 FILLER_7_2516 ();
 sg13g2_decap_8 FILLER_7_2523 ();
 sg13g2_decap_8 FILLER_7_2530 ();
 sg13g2_decap_8 FILLER_7_2537 ();
 sg13g2_decap_8 FILLER_7_2544 ();
 sg13g2_decap_8 FILLER_7_2551 ();
 sg13g2_decap_8 FILLER_7_2558 ();
 sg13g2_decap_8 FILLER_7_2565 ();
 sg13g2_decap_8 FILLER_7_2572 ();
 sg13g2_decap_8 FILLER_7_2579 ();
 sg13g2_decap_8 FILLER_7_2586 ();
 sg13g2_decap_8 FILLER_7_2593 ();
 sg13g2_decap_8 FILLER_7_2600 ();
 sg13g2_decap_8 FILLER_7_2607 ();
 sg13g2_decap_8 FILLER_7_2614 ();
 sg13g2_decap_8 FILLER_7_2621 ();
 sg13g2_decap_8 FILLER_7_2628 ();
 sg13g2_decap_8 FILLER_7_2635 ();
 sg13g2_decap_8 FILLER_7_2642 ();
 sg13g2_decap_8 FILLER_7_2649 ();
 sg13g2_decap_8 FILLER_7_2656 ();
 sg13g2_decap_8 FILLER_7_2663 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_13 ();
 sg13g2_fill_2 FILLER_8_20 ();
 sg13g2_fill_1 FILLER_8_27 ();
 sg13g2_decap_4 FILLER_8_32 ();
 sg13g2_fill_1 FILLER_8_36 ();
 sg13g2_fill_2 FILLER_8_41 ();
 sg13g2_decap_8 FILLER_8_51 ();
 sg13g2_fill_2 FILLER_8_58 ();
 sg13g2_fill_1 FILLER_8_60 ();
 sg13g2_fill_1 FILLER_8_83 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_4 FILLER_8_105 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_fill_1 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_171 ();
 sg13g2_fill_2 FILLER_8_181 ();
 sg13g2_fill_2 FILLER_8_230 ();
 sg13g2_decap_4 FILLER_8_262 ();
 sg13g2_decap_4 FILLER_8_270 ();
 sg13g2_decap_4 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_decap_4 FILLER_8_341 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_368 ();
 sg13g2_fill_1 FILLER_8_370 ();
 sg13g2_fill_2 FILLER_8_377 ();
 sg13g2_fill_1 FILLER_8_379 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_fill_1 FILLER_8_420 ();
 sg13g2_fill_1 FILLER_8_426 ();
 sg13g2_fill_1 FILLER_8_443 ();
 sg13g2_fill_1 FILLER_8_468 ();
 sg13g2_decap_4 FILLER_8_480 ();
 sg13g2_fill_1 FILLER_8_499 ();
 sg13g2_fill_1 FILLER_8_526 ();
 sg13g2_fill_1 FILLER_8_531 ();
 sg13g2_fill_2 FILLER_8_558 ();
 sg13g2_fill_1 FILLER_8_574 ();
 sg13g2_decap_4 FILLER_8_583 ();
 sg13g2_fill_1 FILLER_8_587 ();
 sg13g2_fill_1 FILLER_8_599 ();
 sg13g2_decap_8 FILLER_8_636 ();
 sg13g2_decap_4 FILLER_8_643 ();
 sg13g2_fill_1 FILLER_8_647 ();
 sg13g2_decap_8 FILLER_8_652 ();
 sg13g2_decap_8 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_666 ();
 sg13g2_fill_2 FILLER_8_699 ();
 sg13g2_fill_2 FILLER_8_727 ();
 sg13g2_fill_2 FILLER_8_733 ();
 sg13g2_fill_1 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_762 ();
 sg13g2_fill_2 FILLER_8_769 ();
 sg13g2_decap_4 FILLER_8_781 ();
 sg13g2_fill_2 FILLER_8_785 ();
 sg13g2_decap_8 FILLER_8_827 ();
 sg13g2_decap_8 FILLER_8_834 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_8_908 ();
 sg13g2_decap_4 FILLER_8_915 ();
 sg13g2_fill_1 FILLER_8_919 ();
 sg13g2_fill_1 FILLER_8_1007 ();
 sg13g2_fill_1 FILLER_8_1012 ();
 sg13g2_decap_4 FILLER_8_1039 ();
 sg13g2_fill_2 FILLER_8_1043 ();
 sg13g2_fill_2 FILLER_8_1055 ();
 sg13g2_fill_2 FILLER_8_1061 ();
 sg13g2_decap_8 FILLER_8_1098 ();
 sg13g2_fill_2 FILLER_8_1105 ();
 sg13g2_fill_2 FILLER_8_1141 ();
 sg13g2_fill_2 FILLER_8_1155 ();
 sg13g2_fill_1 FILLER_8_1187 ();
 sg13g2_fill_1 FILLER_8_1222 ();
 sg13g2_fill_1 FILLER_8_1228 ();
 sg13g2_fill_1 FILLER_8_1233 ();
 sg13g2_decap_4 FILLER_8_1276 ();
 sg13g2_decap_8 FILLER_8_1316 ();
 sg13g2_fill_2 FILLER_8_1323 ();
 sg13g2_decap_8 FILLER_8_1334 ();
 sg13g2_decap_8 FILLER_8_1341 ();
 sg13g2_decap_4 FILLER_8_1348 ();
 sg13g2_fill_2 FILLER_8_1386 ();
 sg13g2_fill_2 FILLER_8_1401 ();
 sg13g2_fill_1 FILLER_8_1403 ();
 sg13g2_fill_1 FILLER_8_1429 ();
 sg13g2_fill_2 FILLER_8_1507 ();
 sg13g2_fill_2 FILLER_8_1519 ();
 sg13g2_fill_1 FILLER_8_1521 ();
 sg13g2_fill_2 FILLER_8_1548 ();
 sg13g2_fill_1 FILLER_8_1550 ();
 sg13g2_fill_1 FILLER_8_1592 ();
 sg13g2_fill_1 FILLER_8_1608 ();
 sg13g2_fill_2 FILLER_8_1620 ();
 sg13g2_fill_2 FILLER_8_1659 ();
 sg13g2_fill_2 FILLER_8_1665 ();
 sg13g2_fill_1 FILLER_8_1667 ();
 sg13g2_fill_1 FILLER_8_1687 ();
 sg13g2_fill_2 FILLER_8_1714 ();
 sg13g2_fill_1 FILLER_8_1721 ();
 sg13g2_fill_1 FILLER_8_1728 ();
 sg13g2_decap_4 FILLER_8_1761 ();
 sg13g2_fill_1 FILLER_8_1765 ();
 sg13g2_decap_8 FILLER_8_1770 ();
 sg13g2_decap_4 FILLER_8_1781 ();
 sg13g2_fill_2 FILLER_8_1785 ();
 sg13g2_decap_8 FILLER_8_1824 ();
 sg13g2_fill_2 FILLER_8_1831 ();
 sg13g2_decap_4 FILLER_8_1837 ();
 sg13g2_decap_4 FILLER_8_1845 ();
 sg13g2_fill_1 FILLER_8_1849 ();
 sg13g2_decap_8 FILLER_8_1854 ();
 sg13g2_decap_8 FILLER_8_1861 ();
 sg13g2_decap_4 FILLER_8_1868 ();
 sg13g2_fill_2 FILLER_8_1872 ();
 sg13g2_fill_2 FILLER_8_1879 ();
 sg13g2_fill_1 FILLER_8_1881 ();
 sg13g2_decap_8 FILLER_8_1886 ();
 sg13g2_decap_4 FILLER_8_1893 ();
 sg13g2_fill_2 FILLER_8_1907 ();
 sg13g2_fill_1 FILLER_8_1909 ();
 sg13g2_decap_8 FILLER_8_1914 ();
 sg13g2_fill_2 FILLER_8_1921 ();
 sg13g2_decap_4 FILLER_8_1927 ();
 sg13g2_fill_2 FILLER_8_1931 ();
 sg13g2_fill_2 FILLER_8_1937 ();
 sg13g2_fill_1 FILLER_8_1939 ();
 sg13g2_fill_1 FILLER_8_1974 ();
 sg13g2_fill_2 FILLER_8_2001 ();
 sg13g2_fill_2 FILLER_8_2035 ();
 sg13g2_decap_4 FILLER_8_2084 ();
 sg13g2_fill_1 FILLER_8_2088 ();
 sg13g2_fill_1 FILLER_8_2114 ();
 sg13g2_decap_4 FILLER_8_2119 ();
 sg13g2_fill_2 FILLER_8_2123 ();
 sg13g2_fill_1 FILLER_8_2135 ();
 sg13g2_fill_2 FILLER_8_2146 ();
 sg13g2_fill_1 FILLER_8_2148 ();
 sg13g2_fill_2 FILLER_8_2188 ();
 sg13g2_decap_8 FILLER_8_2236 ();
 sg13g2_fill_2 FILLER_8_2243 ();
 sg13g2_fill_2 FILLER_8_2278 ();
 sg13g2_fill_1 FILLER_8_2354 ();
 sg13g2_decap_4 FILLER_8_2369 ();
 sg13g2_fill_1 FILLER_8_2373 ();
 sg13g2_decap_8 FILLER_8_2434 ();
 sg13g2_decap_8 FILLER_8_2441 ();
 sg13g2_decap_8 FILLER_8_2448 ();
 sg13g2_decap_8 FILLER_8_2455 ();
 sg13g2_decap_8 FILLER_8_2462 ();
 sg13g2_decap_8 FILLER_8_2469 ();
 sg13g2_decap_8 FILLER_8_2476 ();
 sg13g2_decap_8 FILLER_8_2483 ();
 sg13g2_decap_8 FILLER_8_2490 ();
 sg13g2_decap_8 FILLER_8_2497 ();
 sg13g2_decap_8 FILLER_8_2504 ();
 sg13g2_decap_8 FILLER_8_2511 ();
 sg13g2_decap_8 FILLER_8_2518 ();
 sg13g2_decap_8 FILLER_8_2525 ();
 sg13g2_decap_8 FILLER_8_2532 ();
 sg13g2_decap_8 FILLER_8_2539 ();
 sg13g2_decap_8 FILLER_8_2546 ();
 sg13g2_decap_8 FILLER_8_2553 ();
 sg13g2_decap_8 FILLER_8_2560 ();
 sg13g2_decap_8 FILLER_8_2567 ();
 sg13g2_decap_8 FILLER_8_2574 ();
 sg13g2_decap_8 FILLER_8_2581 ();
 sg13g2_decap_8 FILLER_8_2588 ();
 sg13g2_decap_8 FILLER_8_2595 ();
 sg13g2_decap_8 FILLER_8_2602 ();
 sg13g2_decap_8 FILLER_8_2609 ();
 sg13g2_decap_8 FILLER_8_2616 ();
 sg13g2_decap_8 FILLER_8_2623 ();
 sg13g2_decap_8 FILLER_8_2630 ();
 sg13g2_decap_8 FILLER_8_2637 ();
 sg13g2_decap_8 FILLER_8_2644 ();
 sg13g2_decap_8 FILLER_8_2651 ();
 sg13g2_decap_8 FILLER_8_2658 ();
 sg13g2_decap_4 FILLER_8_2665 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_13 ();
 sg13g2_fill_2 FILLER_9_17 ();
 sg13g2_fill_1 FILLER_9_24 ();
 sg13g2_decap_8 FILLER_9_45 ();
 sg13g2_fill_2 FILLER_9_52 ();
 sg13g2_fill_1 FILLER_9_54 ();
 sg13g2_decap_4 FILLER_9_59 ();
 sg13g2_fill_1 FILLER_9_63 ();
 sg13g2_decap_4 FILLER_9_73 ();
 sg13g2_fill_2 FILLER_9_77 ();
 sg13g2_decap_4 FILLER_9_83 ();
 sg13g2_fill_1 FILLER_9_87 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_decap_8 FILLER_9_99 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_120 ();
 sg13g2_decap_4 FILLER_9_127 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_fill_1 FILLER_9_180 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_4 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_4 FILLER_9_259 ();
 sg13g2_fill_2 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_4 FILLER_9_275 ();
 sg13g2_fill_1 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_4 FILLER_9_291 ();
 sg13g2_fill_2 FILLER_9_295 ();
 sg13g2_fill_1 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_fill_2 FILLER_9_321 ();
 sg13g2_decap_4 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_fill_2 FILLER_9_366 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_fill_2 FILLER_9_383 ();
 sg13g2_fill_1 FILLER_9_385 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_422 ();
 sg13g2_decap_8 FILLER_9_429 ();
 sg13g2_fill_2 FILLER_9_436 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_fill_1 FILLER_9_475 ();
 sg13g2_fill_1 FILLER_9_480 ();
 sg13g2_fill_1 FILLER_9_495 ();
 sg13g2_fill_2 FILLER_9_505 ();
 sg13g2_fill_1 FILLER_9_507 ();
 sg13g2_decap_4 FILLER_9_512 ();
 sg13g2_fill_1 FILLER_9_516 ();
 sg13g2_fill_2 FILLER_9_582 ();
 sg13g2_fill_1 FILLER_9_584 ();
 sg13g2_fill_1 FILLER_9_591 ();
 sg13g2_fill_2 FILLER_9_598 ();
 sg13g2_decap_4 FILLER_9_613 ();
 sg13g2_fill_2 FILLER_9_617 ();
 sg13g2_decap_4 FILLER_9_623 ();
 sg13g2_decap_4 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_667 ();
 sg13g2_fill_1 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_722 ();
 sg13g2_decap_8 FILLER_9_729 ();
 sg13g2_fill_1 FILLER_9_736 ();
 sg13g2_decap_4 FILLER_9_751 ();
 sg13g2_fill_2 FILLER_9_755 ();
 sg13g2_fill_2 FILLER_9_788 ();
 sg13g2_fill_1 FILLER_9_790 ();
 sg13g2_fill_1 FILLER_9_838 ();
 sg13g2_decap_4 FILLER_9_843 ();
 sg13g2_fill_2 FILLER_9_881 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_8 FILLER_9_900 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_fill_1 FILLER_9_914 ();
 sg13g2_fill_2 FILLER_9_955 ();
 sg13g2_fill_1 FILLER_9_957 ();
 sg13g2_decap_4 FILLER_9_1015 ();
 sg13g2_decap_4 FILLER_9_1029 ();
 sg13g2_fill_2 FILLER_9_1033 ();
 sg13g2_fill_2 FILLER_9_1050 ();
 sg13g2_fill_1 FILLER_9_1052 ();
 sg13g2_decap_4 FILLER_9_1079 ();
 sg13g2_fill_1 FILLER_9_1083 ();
 sg13g2_decap_8 FILLER_9_1088 ();
 sg13g2_decap_8 FILLER_9_1095 ();
 sg13g2_fill_2 FILLER_9_1102 ();
 sg13g2_fill_2 FILLER_9_1148 ();
 sg13g2_fill_2 FILLER_9_1154 ();
 sg13g2_fill_1 FILLER_9_1156 ();
 sg13g2_decap_8 FILLER_9_1173 ();
 sg13g2_fill_2 FILLER_9_1180 ();
 sg13g2_fill_1 FILLER_9_1182 ();
 sg13g2_decap_4 FILLER_9_1191 ();
 sg13g2_fill_2 FILLER_9_1199 ();
 sg13g2_fill_1 FILLER_9_1201 ();
 sg13g2_fill_1 FILLER_9_1232 ();
 sg13g2_fill_1 FILLER_9_1245 ();
 sg13g2_decap_8 FILLER_9_1250 ();
 sg13g2_decap_4 FILLER_9_1257 ();
 sg13g2_fill_1 FILLER_9_1287 ();
 sg13g2_fill_1 FILLER_9_1314 ();
 sg13g2_fill_1 FILLER_9_1346 ();
 sg13g2_fill_2 FILLER_9_1351 ();
 sg13g2_fill_1 FILLER_9_1353 ();
 sg13g2_fill_1 FILLER_9_1411 ();
 sg13g2_decap_4 FILLER_9_1451 ();
 sg13g2_decap_8 FILLER_9_1469 ();
 sg13g2_decap_4 FILLER_9_1486 ();
 sg13g2_fill_1 FILLER_9_1490 ();
 sg13g2_decap_8 FILLER_9_1517 ();
 sg13g2_decap_4 FILLER_9_1524 ();
 sg13g2_fill_2 FILLER_9_1528 ();
 sg13g2_fill_2 FILLER_9_1534 ();
 sg13g2_fill_1 FILLER_9_1536 ();
 sg13g2_decap_4 FILLER_9_1546 ();
 sg13g2_fill_1 FILLER_9_1550 ();
 sg13g2_fill_2 FILLER_9_1568 ();
 sg13g2_fill_2 FILLER_9_1574 ();
 sg13g2_fill_1 FILLER_9_1604 ();
 sg13g2_fill_1 FILLER_9_1628 ();
 sg13g2_decap_8 FILLER_9_1638 ();
 sg13g2_fill_2 FILLER_9_1645 ();
 sg13g2_fill_1 FILLER_9_1647 ();
 sg13g2_fill_1 FILLER_9_1654 ();
 sg13g2_fill_1 FILLER_9_1662 ();
 sg13g2_fill_1 FILLER_9_1668 ();
 sg13g2_fill_2 FILLER_9_1704 ();
 sg13g2_fill_2 FILLER_9_1711 ();
 sg13g2_decap_4 FILLER_9_1722 ();
 sg13g2_fill_2 FILLER_9_1726 ();
 sg13g2_decap_8 FILLER_9_1736 ();
 sg13g2_fill_1 FILLER_9_1743 ();
 sg13g2_decap_8 FILLER_9_1748 ();
 sg13g2_decap_8 FILLER_9_1755 ();
 sg13g2_decap_8 FILLER_9_1762 ();
 sg13g2_decap_8 FILLER_9_1769 ();
 sg13g2_decap_8 FILLER_9_1776 ();
 sg13g2_decap_4 FILLER_9_1783 ();
 sg13g2_decap_8 FILLER_9_1805 ();
 sg13g2_decap_8 FILLER_9_1812 ();
 sg13g2_decap_8 FILLER_9_1819 ();
 sg13g2_decap_8 FILLER_9_1826 ();
 sg13g2_decap_4 FILLER_9_1833 ();
 sg13g2_decap_8 FILLER_9_1917 ();
 sg13g2_fill_1 FILLER_9_1924 ();
 sg13g2_fill_1 FILLER_9_1937 ();
 sg13g2_fill_2 FILLER_9_1954 ();
 sg13g2_fill_2 FILLER_9_1977 ();
 sg13g2_fill_1 FILLER_9_2030 ();
 sg13g2_fill_1 FILLER_9_2069 ();
 sg13g2_fill_2 FILLER_9_2074 ();
 sg13g2_fill_1 FILLER_9_2086 ();
 sg13g2_decap_8 FILLER_9_2108 ();
 sg13g2_decap_8 FILLER_9_2115 ();
 sg13g2_decap_8 FILLER_9_2122 ();
 sg13g2_decap_8 FILLER_9_2129 ();
 sg13g2_decap_4 FILLER_9_2136 ();
 sg13g2_fill_2 FILLER_9_2140 ();
 sg13g2_decap_8 FILLER_9_2166 ();
 sg13g2_fill_2 FILLER_9_2173 ();
 sg13g2_fill_1 FILLER_9_2175 ();
 sg13g2_fill_1 FILLER_9_2186 ();
 sg13g2_fill_1 FILLER_9_2197 ();
 sg13g2_fill_1 FILLER_9_2208 ();
 sg13g2_fill_2 FILLER_9_2219 ();
 sg13g2_fill_1 FILLER_9_2221 ();
 sg13g2_fill_2 FILLER_9_2278 ();
 sg13g2_decap_8 FILLER_9_2333 ();
 sg13g2_decap_8 FILLER_9_2340 ();
 sg13g2_decap_8 FILLER_9_2347 ();
 sg13g2_fill_2 FILLER_9_2354 ();
 sg13g2_fill_1 FILLER_9_2356 ();
 sg13g2_decap_8 FILLER_9_2377 ();
 sg13g2_fill_1 FILLER_9_2405 ();
 sg13g2_decap_8 FILLER_9_2445 ();
 sg13g2_decap_8 FILLER_9_2452 ();
 sg13g2_decap_8 FILLER_9_2459 ();
 sg13g2_decap_8 FILLER_9_2466 ();
 sg13g2_decap_8 FILLER_9_2473 ();
 sg13g2_decap_8 FILLER_9_2480 ();
 sg13g2_decap_8 FILLER_9_2487 ();
 sg13g2_decap_8 FILLER_9_2494 ();
 sg13g2_decap_8 FILLER_9_2501 ();
 sg13g2_decap_8 FILLER_9_2508 ();
 sg13g2_decap_8 FILLER_9_2515 ();
 sg13g2_decap_8 FILLER_9_2522 ();
 sg13g2_decap_8 FILLER_9_2529 ();
 sg13g2_decap_8 FILLER_9_2536 ();
 sg13g2_decap_8 FILLER_9_2543 ();
 sg13g2_decap_8 FILLER_9_2550 ();
 sg13g2_decap_8 FILLER_9_2557 ();
 sg13g2_decap_8 FILLER_9_2564 ();
 sg13g2_decap_8 FILLER_9_2571 ();
 sg13g2_decap_8 FILLER_9_2578 ();
 sg13g2_decap_8 FILLER_9_2585 ();
 sg13g2_decap_8 FILLER_9_2592 ();
 sg13g2_decap_8 FILLER_9_2599 ();
 sg13g2_decap_8 FILLER_9_2606 ();
 sg13g2_decap_8 FILLER_9_2613 ();
 sg13g2_decap_8 FILLER_9_2620 ();
 sg13g2_decap_8 FILLER_9_2627 ();
 sg13g2_decap_8 FILLER_9_2634 ();
 sg13g2_decap_8 FILLER_9_2641 ();
 sg13g2_decap_8 FILLER_9_2648 ();
 sg13g2_decap_8 FILLER_9_2655 ();
 sg13g2_decap_8 FILLER_9_2662 ();
 sg13g2_fill_1 FILLER_9_2669 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_67 ();
 sg13g2_fill_1 FILLER_10_82 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_2 FILLER_10_116 ();
 sg13g2_decap_4 FILLER_10_149 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_4 FILLER_10_354 ();
 sg13g2_fill_2 FILLER_10_392 ();
 sg13g2_fill_1 FILLER_10_394 ();
 sg13g2_decap_4 FILLER_10_415 ();
 sg13g2_fill_2 FILLER_10_423 ();
 sg13g2_fill_1 FILLER_10_425 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_fill_1 FILLER_10_438 ();
 sg13g2_decap_4 FILLER_10_455 ();
 sg13g2_fill_2 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_495 ();
 sg13g2_decap_8 FILLER_10_502 ();
 sg13g2_fill_2 FILLER_10_509 ();
 sg13g2_decap_4 FILLER_10_519 ();
 sg13g2_fill_1 FILLER_10_523 ();
 sg13g2_decap_8 FILLER_10_552 ();
 sg13g2_decap_8 FILLER_10_559 ();
 sg13g2_fill_2 FILLER_10_566 ();
 sg13g2_fill_1 FILLER_10_568 ();
 sg13g2_fill_2 FILLER_10_577 ();
 sg13g2_fill_2 FILLER_10_584 ();
 sg13g2_fill_1 FILLER_10_586 ();
 sg13g2_fill_2 FILLER_10_591 ();
 sg13g2_fill_1 FILLER_10_593 ();
 sg13g2_decap_8 FILLER_10_600 ();
 sg13g2_decap_8 FILLER_10_607 ();
 sg13g2_decap_8 FILLER_10_614 ();
 sg13g2_decap_8 FILLER_10_621 ();
 sg13g2_decap_4 FILLER_10_628 ();
 sg13g2_fill_1 FILLER_10_632 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_fill_2 FILLER_10_679 ();
 sg13g2_fill_1 FILLER_10_681 ();
 sg13g2_decap_4 FILLER_10_686 ();
 sg13g2_fill_2 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_702 ();
 sg13g2_decap_4 FILLER_10_709 ();
 sg13g2_decap_4 FILLER_10_717 ();
 sg13g2_fill_2 FILLER_10_721 ();
 sg13g2_fill_2 FILLER_10_733 ();
 sg13g2_fill_1 FILLER_10_735 ();
 sg13g2_decap_4 FILLER_10_788 ();
 sg13g2_decap_4 FILLER_10_828 ();
 sg13g2_fill_1 FILLER_10_832 ();
 sg13g2_decap_8 FILLER_10_863 ();
 sg13g2_fill_2 FILLER_10_870 ();
 sg13g2_fill_1 FILLER_10_872 ();
 sg13g2_decap_4 FILLER_10_883 ();
 sg13g2_fill_2 FILLER_10_887 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_fill_1 FILLER_10_936 ();
 sg13g2_fill_2 FILLER_10_945 ();
 sg13g2_fill_1 FILLER_10_947 ();
 sg13g2_decap_4 FILLER_10_958 ();
 sg13g2_fill_1 FILLER_10_962 ();
 sg13g2_decap_8 FILLER_10_985 ();
 sg13g2_decap_8 FILLER_10_992 ();
 sg13g2_decap_8 FILLER_10_999 ();
 sg13g2_decap_8 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1013 ();
 sg13g2_fill_2 FILLER_10_1020 ();
 sg13g2_fill_1 FILLER_10_1022 ();
 sg13g2_decap_8 FILLER_10_1033 ();
 sg13g2_decap_8 FILLER_10_1040 ();
 sg13g2_fill_2 FILLER_10_1103 ();
 sg13g2_fill_2 FILLER_10_1131 ();
 sg13g2_fill_1 FILLER_10_1133 ();
 sg13g2_fill_2 FILLER_10_1165 ();
 sg13g2_fill_1 FILLER_10_1172 ();
 sg13g2_fill_2 FILLER_10_1177 ();
 sg13g2_fill_1 FILLER_10_1179 ();
 sg13g2_fill_2 FILLER_10_1184 ();
 sg13g2_fill_1 FILLER_10_1186 ();
 sg13g2_decap_8 FILLER_10_1191 ();
 sg13g2_decap_8 FILLER_10_1198 ();
 sg13g2_decap_8 FILLER_10_1205 ();
 sg13g2_fill_2 FILLER_10_1252 ();
 sg13g2_fill_2 FILLER_10_1258 ();
 sg13g2_fill_2 FILLER_10_1273 ();
 sg13g2_decap_4 FILLER_10_1313 ();
 sg13g2_fill_1 FILLER_10_1317 ();
 sg13g2_fill_1 FILLER_10_1322 ();
 sg13g2_fill_1 FILLER_10_1328 ();
 sg13g2_fill_1 FILLER_10_1369 ();
 sg13g2_decap_8 FILLER_10_1374 ();
 sg13g2_decap_8 FILLER_10_1407 ();
 sg13g2_fill_2 FILLER_10_1414 ();
 sg13g2_decap_4 FILLER_10_1449 ();
 sg13g2_fill_2 FILLER_10_1458 ();
 sg13g2_fill_1 FILLER_10_1460 ();
 sg13g2_decap_8 FILLER_10_1473 ();
 sg13g2_decap_8 FILLER_10_1491 ();
 sg13g2_fill_1 FILLER_10_1502 ();
 sg13g2_decap_8 FILLER_10_1518 ();
 sg13g2_decap_8 FILLER_10_1525 ();
 sg13g2_fill_2 FILLER_10_1532 ();
 sg13g2_fill_1 FILLER_10_1534 ();
 sg13g2_decap_8 FILLER_10_1539 ();
 sg13g2_fill_2 FILLER_10_1546 ();
 sg13g2_fill_2 FILLER_10_1552 ();
 sg13g2_fill_1 FILLER_10_1554 ();
 sg13g2_decap_4 FILLER_10_1563 ();
 sg13g2_fill_2 FILLER_10_1578 ();
 sg13g2_fill_1 FILLER_10_1580 ();
 sg13g2_decap_4 FILLER_10_1607 ();
 sg13g2_fill_2 FILLER_10_1611 ();
 sg13g2_decap_4 FILLER_10_1617 ();
 sg13g2_fill_1 FILLER_10_1631 ();
 sg13g2_fill_2 FILLER_10_1636 ();
 sg13g2_decap_8 FILLER_10_1647 ();
 sg13g2_decap_4 FILLER_10_1654 ();
 sg13g2_fill_2 FILLER_10_1658 ();
 sg13g2_decap_8 FILLER_10_1664 ();
 sg13g2_decap_4 FILLER_10_1671 ();
 sg13g2_decap_8 FILLER_10_1679 ();
 sg13g2_decap_4 FILLER_10_1690 ();
 sg13g2_decap_4 FILLER_10_1700 ();
 sg13g2_fill_2 FILLER_10_1708 ();
 sg13g2_fill_1 FILLER_10_1710 ();
 sg13g2_fill_2 FILLER_10_1715 ();
 sg13g2_fill_1 FILLER_10_1717 ();
 sg13g2_fill_2 FILLER_10_1723 ();
 sg13g2_decap_8 FILLER_10_1729 ();
 sg13g2_decap_8 FILLER_10_1736 ();
 sg13g2_fill_2 FILLER_10_1743 ();
 sg13g2_fill_1 FILLER_10_1745 ();
 sg13g2_decap_8 FILLER_10_1756 ();
 sg13g2_fill_1 FILLER_10_1763 ();
 sg13g2_decap_8 FILLER_10_1768 ();
 sg13g2_decap_8 FILLER_10_1811 ();
 sg13g2_decap_8 FILLER_10_1818 ();
 sg13g2_decap_4 FILLER_10_1825 ();
 sg13g2_fill_2 FILLER_10_1859 ();
 sg13g2_fill_2 FILLER_10_1887 ();
 sg13g2_fill_1 FILLER_10_1889 ();
 sg13g2_fill_2 FILLER_10_1916 ();
 sg13g2_fill_1 FILLER_10_1943 ();
 sg13g2_fill_2 FILLER_10_1948 ();
 sg13g2_fill_1 FILLER_10_1950 ();
 sg13g2_fill_2 FILLER_10_1961 ();
 sg13g2_fill_1 FILLER_10_1963 ();
 sg13g2_decap_4 FILLER_10_2002 ();
 sg13g2_fill_1 FILLER_10_2006 ();
 sg13g2_fill_1 FILLER_10_2044 ();
 sg13g2_fill_1 FILLER_10_2073 ();
 sg13g2_decap_8 FILLER_10_2095 ();
 sg13g2_fill_2 FILLER_10_2102 ();
 sg13g2_fill_1 FILLER_10_2104 ();
 sg13g2_fill_2 FILLER_10_2109 ();
 sg13g2_fill_1 FILLER_10_2111 ();
 sg13g2_fill_1 FILLER_10_2120 ();
 sg13g2_fill_2 FILLER_10_2131 ();
 sg13g2_fill_1 FILLER_10_2133 ();
 sg13g2_decap_8 FILLER_10_2138 ();
 sg13g2_decap_8 FILLER_10_2145 ();
 sg13g2_fill_2 FILLER_10_2152 ();
 sg13g2_fill_1 FILLER_10_2154 ();
 sg13g2_fill_2 FILLER_10_2165 ();
 sg13g2_decap_8 FILLER_10_2197 ();
 sg13g2_decap_8 FILLER_10_2204 ();
 sg13g2_decap_4 FILLER_10_2211 ();
 sg13g2_decap_4 FILLER_10_2241 ();
 sg13g2_decap_8 FILLER_10_2258 ();
 sg13g2_decap_4 FILLER_10_2312 ();
 sg13g2_fill_1 FILLER_10_2316 ();
 sg13g2_fill_1 FILLER_10_2320 ();
 sg13g2_decap_8 FILLER_10_2361 ();
 sg13g2_decap_8 FILLER_10_2368 ();
 sg13g2_decap_8 FILLER_10_2375 ();
 sg13g2_decap_8 FILLER_10_2382 ();
 sg13g2_fill_1 FILLER_10_2389 ();
 sg13g2_decap_8 FILLER_10_2400 ();
 sg13g2_decap_8 FILLER_10_2407 ();
 sg13g2_decap_8 FILLER_10_2414 ();
 sg13g2_decap_8 FILLER_10_2421 ();
 sg13g2_decap_8 FILLER_10_2428 ();
 sg13g2_decap_8 FILLER_10_2435 ();
 sg13g2_decap_8 FILLER_10_2442 ();
 sg13g2_decap_8 FILLER_10_2449 ();
 sg13g2_decap_8 FILLER_10_2456 ();
 sg13g2_decap_8 FILLER_10_2463 ();
 sg13g2_decap_8 FILLER_10_2470 ();
 sg13g2_decap_8 FILLER_10_2477 ();
 sg13g2_decap_8 FILLER_10_2484 ();
 sg13g2_decap_8 FILLER_10_2491 ();
 sg13g2_decap_8 FILLER_10_2498 ();
 sg13g2_decap_8 FILLER_10_2505 ();
 sg13g2_decap_8 FILLER_10_2512 ();
 sg13g2_decap_8 FILLER_10_2519 ();
 sg13g2_decap_8 FILLER_10_2526 ();
 sg13g2_decap_8 FILLER_10_2533 ();
 sg13g2_decap_8 FILLER_10_2540 ();
 sg13g2_decap_8 FILLER_10_2547 ();
 sg13g2_decap_8 FILLER_10_2554 ();
 sg13g2_decap_8 FILLER_10_2561 ();
 sg13g2_decap_8 FILLER_10_2568 ();
 sg13g2_decap_8 FILLER_10_2575 ();
 sg13g2_decap_8 FILLER_10_2582 ();
 sg13g2_decap_8 FILLER_10_2589 ();
 sg13g2_decap_8 FILLER_10_2596 ();
 sg13g2_decap_8 FILLER_10_2603 ();
 sg13g2_decap_8 FILLER_10_2610 ();
 sg13g2_decap_8 FILLER_10_2617 ();
 sg13g2_decap_8 FILLER_10_2624 ();
 sg13g2_decap_8 FILLER_10_2631 ();
 sg13g2_decap_8 FILLER_10_2638 ();
 sg13g2_decap_8 FILLER_10_2645 ();
 sg13g2_decap_8 FILLER_10_2652 ();
 sg13g2_decap_8 FILLER_10_2659 ();
 sg13g2_decap_4 FILLER_10_2666 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_fill_2 FILLER_11_184 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_fill_1 FILLER_11_298 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_4 FILLER_11_383 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_4 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_472 ();
 sg13g2_decap_4 FILLER_11_479 ();
 sg13g2_fill_1 FILLER_11_483 ();
 sg13g2_decap_4 FILLER_11_488 ();
 sg13g2_fill_1 FILLER_11_492 ();
 sg13g2_fill_2 FILLER_11_521 ();
 sg13g2_fill_2 FILLER_11_531 ();
 sg13g2_fill_1 FILLER_11_533 ();
 sg13g2_decap_8 FILLER_11_540 ();
 sg13g2_decap_8 FILLER_11_547 ();
 sg13g2_decap_4 FILLER_11_565 ();
 sg13g2_fill_1 FILLER_11_569 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_4 FILLER_11_620 ();
 sg13g2_fill_2 FILLER_11_624 ();
 sg13g2_fill_1 FILLER_11_682 ();
 sg13g2_decap_8 FILLER_11_687 ();
 sg13g2_decap_8 FILLER_11_694 ();
 sg13g2_decap_4 FILLER_11_701 ();
 sg13g2_fill_2 FILLER_11_705 ();
 sg13g2_fill_2 FILLER_11_743 ();
 sg13g2_fill_1 FILLER_11_745 ();
 sg13g2_fill_2 FILLER_11_750 ();
 sg13g2_fill_1 FILLER_11_792 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_fill_2 FILLER_11_843 ();
 sg13g2_fill_1 FILLER_11_845 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_8 FILLER_11_857 ();
 sg13g2_decap_8 FILLER_11_864 ();
 sg13g2_decap_4 FILLER_11_871 ();
 sg13g2_fill_1 FILLER_11_875 ();
 sg13g2_fill_2 FILLER_11_912 ();
 sg13g2_fill_1 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_941 ();
 sg13g2_decap_8 FILLER_11_948 ();
 sg13g2_decap_4 FILLER_11_955 ();
 sg13g2_fill_1 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_975 ();
 sg13g2_decap_8 FILLER_11_982 ();
 sg13g2_fill_1 FILLER_11_989 ();
 sg13g2_decap_4 FILLER_11_995 ();
 sg13g2_fill_2 FILLER_11_999 ();
 sg13g2_decap_4 FILLER_11_1037 ();
 sg13g2_fill_1 FILLER_11_1051 ();
 sg13g2_fill_1 FILLER_11_1078 ();
 sg13g2_fill_2 FILLER_11_1201 ();
 sg13g2_fill_1 FILLER_11_1207 ();
 sg13g2_fill_1 FILLER_11_1217 ();
 sg13g2_fill_1 FILLER_11_1226 ();
 sg13g2_decap_8 FILLER_11_1257 ();
 sg13g2_fill_2 FILLER_11_1264 ();
 sg13g2_decap_4 FILLER_11_1279 ();
 sg13g2_fill_2 FILLER_11_1287 ();
 sg13g2_fill_1 FILLER_11_1289 ();
 sg13g2_fill_2 FILLER_11_1294 ();
 sg13g2_fill_1 FILLER_11_1296 ();
 sg13g2_decap_8 FILLER_11_1301 ();
 sg13g2_fill_2 FILLER_11_1308 ();
 sg13g2_decap_4 FILLER_11_1357 ();
 sg13g2_fill_2 FILLER_11_1361 ();
 sg13g2_decap_8 FILLER_11_1367 ();
 sg13g2_decap_4 FILLER_11_1374 ();
 sg13g2_fill_1 FILLER_11_1378 ();
 sg13g2_decap_8 FILLER_11_1384 ();
 sg13g2_decap_8 FILLER_11_1405 ();
 sg13g2_decap_4 FILLER_11_1426 ();
 sg13g2_fill_2 FILLER_11_1430 ();
 sg13g2_fill_1 FILLER_11_1444 ();
 sg13g2_fill_1 FILLER_11_1454 ();
 sg13g2_fill_1 FILLER_11_1459 ();
 sg13g2_fill_1 FILLER_11_1470 ();
 sg13g2_fill_1 FILLER_11_1483 ();
 sg13g2_fill_2 FILLER_11_1525 ();
 sg13g2_fill_1 FILLER_11_1527 ();
 sg13g2_decap_4 FILLER_11_1541 ();
 sg13g2_fill_1 FILLER_11_1571 ();
 sg13g2_fill_1 FILLER_11_1582 ();
 sg13g2_fill_1 FILLER_11_1588 ();
 sg13g2_decap_8 FILLER_11_1642 ();
 sg13g2_fill_1 FILLER_11_1649 ();
 sg13g2_fill_2 FILLER_11_1654 ();
 sg13g2_fill_1 FILLER_11_1656 ();
 sg13g2_decap_4 FILLER_11_1662 ();
 sg13g2_fill_1 FILLER_11_1666 ();
 sg13g2_decap_4 FILLER_11_1672 ();
 sg13g2_fill_1 FILLER_11_1676 ();
 sg13g2_fill_1 FILLER_11_1687 ();
 sg13g2_fill_1 FILLER_11_1709 ();
 sg13g2_fill_2 FILLER_11_1757 ();
 sg13g2_fill_1 FILLER_11_1759 ();
 sg13g2_fill_1 FILLER_11_1816 ();
 sg13g2_decap_4 FILLER_11_1863 ();
 sg13g2_fill_1 FILLER_11_1871 ();
 sg13g2_decap_4 FILLER_11_1931 ();
 sg13g2_fill_1 FILLER_11_1935 ();
 sg13g2_fill_2 FILLER_11_1940 ();
 sg13g2_fill_1 FILLER_11_1942 ();
 sg13g2_decap_4 FILLER_11_1946 ();
 sg13g2_fill_2 FILLER_11_1950 ();
 sg13g2_fill_2 FILLER_11_1956 ();
 sg13g2_fill_1 FILLER_11_1958 ();
 sg13g2_fill_2 FILLER_11_1985 ();
 sg13g2_decap_4 FILLER_11_1997 ();
 sg13g2_decap_8 FILLER_11_2011 ();
 sg13g2_fill_2 FILLER_11_2086 ();
 sg13g2_fill_1 FILLER_11_2124 ();
 sg13g2_decap_4 FILLER_11_2129 ();
 sg13g2_decap_8 FILLER_11_2190 ();
 sg13g2_decap_4 FILLER_11_2197 ();
 sg13g2_decap_8 FILLER_11_2211 ();
 sg13g2_decap_8 FILLER_11_2218 ();
 sg13g2_decap_8 FILLER_11_2225 ();
 sg13g2_decap_8 FILLER_11_2232 ();
 sg13g2_fill_1 FILLER_11_2239 ();
 sg13g2_fill_1 FILLER_11_2276 ();
 sg13g2_decap_8 FILLER_11_2297 ();
 sg13g2_fill_2 FILLER_11_2304 ();
 sg13g2_decap_8 FILLER_11_2363 ();
 sg13g2_decap_4 FILLER_11_2370 ();
 sg13g2_decap_8 FILLER_11_2384 ();
 sg13g2_decap_4 FILLER_11_2391 ();
 sg13g2_fill_2 FILLER_11_2395 ();
 sg13g2_decap_8 FILLER_11_2423 ();
 sg13g2_decap_8 FILLER_11_2430 ();
 sg13g2_decap_8 FILLER_11_2437 ();
 sg13g2_decap_8 FILLER_11_2444 ();
 sg13g2_decap_8 FILLER_11_2451 ();
 sg13g2_decap_8 FILLER_11_2458 ();
 sg13g2_decap_8 FILLER_11_2465 ();
 sg13g2_decap_8 FILLER_11_2472 ();
 sg13g2_decap_8 FILLER_11_2479 ();
 sg13g2_decap_8 FILLER_11_2486 ();
 sg13g2_decap_8 FILLER_11_2493 ();
 sg13g2_decap_8 FILLER_11_2500 ();
 sg13g2_decap_8 FILLER_11_2507 ();
 sg13g2_decap_8 FILLER_11_2514 ();
 sg13g2_decap_8 FILLER_11_2521 ();
 sg13g2_decap_8 FILLER_11_2528 ();
 sg13g2_decap_8 FILLER_11_2535 ();
 sg13g2_decap_8 FILLER_11_2542 ();
 sg13g2_decap_8 FILLER_11_2549 ();
 sg13g2_decap_8 FILLER_11_2556 ();
 sg13g2_decap_8 FILLER_11_2563 ();
 sg13g2_decap_8 FILLER_11_2570 ();
 sg13g2_decap_8 FILLER_11_2577 ();
 sg13g2_decap_8 FILLER_11_2584 ();
 sg13g2_decap_8 FILLER_11_2591 ();
 sg13g2_decap_8 FILLER_11_2598 ();
 sg13g2_decap_8 FILLER_11_2605 ();
 sg13g2_decap_8 FILLER_11_2612 ();
 sg13g2_decap_8 FILLER_11_2619 ();
 sg13g2_decap_8 FILLER_11_2626 ();
 sg13g2_decap_8 FILLER_11_2633 ();
 sg13g2_decap_8 FILLER_11_2640 ();
 sg13g2_decap_8 FILLER_11_2647 ();
 sg13g2_decap_8 FILLER_11_2654 ();
 sg13g2_decap_8 FILLER_11_2661 ();
 sg13g2_fill_2 FILLER_11_2668 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_12 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_decap_4 FILLER_12_64 ();
 sg13g2_fill_1 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_86 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_200 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_decap_4 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_252 ();
 sg13g2_fill_1 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_268 ();
 sg13g2_fill_2 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_decap_4 FILLER_12_311 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_fill_2 FILLER_12_351 ();
 sg13g2_decap_4 FILLER_12_361 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_decap_4 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_fill_2 FILLER_12_396 ();
 sg13g2_fill_2 FILLER_12_416 ();
 sg13g2_fill_1 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_fill_1 FILLER_12_515 ();
 sg13g2_fill_2 FILLER_12_538 ();
 sg13g2_decap_8 FILLER_12_544 ();
 sg13g2_decap_4 FILLER_12_551 ();
 sg13g2_fill_2 FILLER_12_555 ();
 sg13g2_decap_4 FILLER_12_603 ();
 sg13g2_fill_1 FILLER_12_607 ();
 sg13g2_decap_4 FILLER_12_621 ();
 sg13g2_fill_1 FILLER_12_625 ();
 sg13g2_fill_2 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_decap_4 FILLER_12_691 ();
 sg13g2_fill_2 FILLER_12_695 ();
 sg13g2_fill_2 FILLER_12_727 ();
 sg13g2_decap_4 FILLER_12_768 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_797 ();
 sg13g2_decap_4 FILLER_12_814 ();
 sg13g2_fill_2 FILLER_12_886 ();
 sg13g2_fill_1 FILLER_12_924 ();
 sg13g2_fill_1 FILLER_12_951 ();
 sg13g2_fill_1 FILLER_12_978 ();
 sg13g2_fill_1 FILLER_12_1048 ();
 sg13g2_fill_2 FILLER_12_1063 ();
 sg13g2_fill_1 FILLER_12_1065 ();
 sg13g2_fill_2 FILLER_12_1070 ();
 sg13g2_fill_2 FILLER_12_1082 ();
 sg13g2_fill_1 FILLER_12_1105 ();
 sg13g2_fill_1 FILLER_12_1118 ();
 sg13g2_fill_2 FILLER_12_1149 ();
 sg13g2_fill_1 FILLER_12_1151 ();
 sg13g2_fill_1 FILLER_12_1157 ();
 sg13g2_decap_4 FILLER_12_1257 ();
 sg13g2_fill_2 FILLER_12_1261 ();
 sg13g2_fill_2 FILLER_12_1276 ();
 sg13g2_decap_8 FILLER_12_1282 ();
 sg13g2_decap_8 FILLER_12_1289 ();
 sg13g2_fill_1 FILLER_12_1296 ();
 sg13g2_decap_4 FILLER_12_1301 ();
 sg13g2_fill_2 FILLER_12_1305 ();
 sg13g2_decap_8 FILLER_12_1337 ();
 sg13g2_fill_2 FILLER_12_1344 ();
 sg13g2_decap_8 FILLER_12_1367 ();
 sg13g2_fill_2 FILLER_12_1374 ();
 sg13g2_fill_1 FILLER_12_1376 ();
 sg13g2_decap_8 FILLER_12_1413 ();
 sg13g2_decap_8 FILLER_12_1420 ();
 sg13g2_decap_8 FILLER_12_1427 ();
 sg13g2_fill_1 FILLER_12_1434 ();
 sg13g2_decap_4 FILLER_12_1510 ();
 sg13g2_fill_2 FILLER_12_1519 ();
 sg13g2_decap_8 FILLER_12_1526 ();
 sg13g2_decap_4 FILLER_12_1533 ();
 sg13g2_fill_2 FILLER_12_1537 ();
 sg13g2_fill_1 FILLER_12_1543 ();
 sg13g2_fill_1 FILLER_12_1570 ();
 sg13g2_fill_1 FILLER_12_1581 ();
 sg13g2_decap_4 FILLER_12_1592 ();
 sg13g2_fill_1 FILLER_12_1596 ();
 sg13g2_fill_2 FILLER_12_1601 ();
 sg13g2_fill_1 FILLER_12_1603 ();
 sg13g2_fill_1 FILLER_12_1624 ();
 sg13g2_fill_1 FILLER_12_1633 ();
 sg13g2_fill_1 FILLER_12_1645 ();
 sg13g2_fill_1 FILLER_12_1651 ();
 sg13g2_fill_1 FILLER_12_1704 ();
 sg13g2_decap_4 FILLER_12_1757 ();
 sg13g2_fill_1 FILLER_12_1796 ();
 sg13g2_fill_2 FILLER_12_1831 ();
 sg13g2_fill_1 FILLER_12_1833 ();
 sg13g2_fill_2 FILLER_12_1860 ();
 sg13g2_decap_4 FILLER_12_1877 ();
 sg13g2_fill_1 FILLER_12_1881 ();
 sg13g2_decap_8 FILLER_12_1886 ();
 sg13g2_fill_2 FILLER_12_1901 ();
 sg13g2_fill_1 FILLER_12_1939 ();
 sg13g2_fill_1 FILLER_12_2008 ();
 sg13g2_fill_2 FILLER_12_2059 ();
 sg13g2_fill_1 FILLER_12_2094 ();
 sg13g2_fill_2 FILLER_12_2100 ();
 sg13g2_fill_1 FILLER_12_2102 ();
 sg13g2_fill_2 FILLER_12_2113 ();
 sg13g2_fill_1 FILLER_12_2115 ();
 sg13g2_fill_2 FILLER_12_2168 ();
 sg13g2_fill_1 FILLER_12_2170 ();
 sg13g2_decap_8 FILLER_12_2179 ();
 sg13g2_decap_4 FILLER_12_2186 ();
 sg13g2_fill_1 FILLER_12_2190 ();
 sg13g2_decap_4 FILLER_12_2201 ();
 sg13g2_decap_4 FILLER_12_2261 ();
 sg13g2_fill_1 FILLER_12_2265 ();
 sg13g2_fill_2 FILLER_12_2270 ();
 sg13g2_fill_1 FILLER_12_2282 ();
 sg13g2_fill_1 FILLER_12_2309 ();
 sg13g2_fill_2 FILLER_12_2314 ();
 sg13g2_fill_1 FILLER_12_2326 ();
 sg13g2_fill_2 FILLER_12_2353 ();
 sg13g2_decap_8 FILLER_12_2433 ();
 sg13g2_decap_8 FILLER_12_2440 ();
 sg13g2_decap_8 FILLER_12_2447 ();
 sg13g2_decap_8 FILLER_12_2454 ();
 sg13g2_decap_8 FILLER_12_2461 ();
 sg13g2_decap_8 FILLER_12_2468 ();
 sg13g2_decap_8 FILLER_12_2475 ();
 sg13g2_decap_8 FILLER_12_2482 ();
 sg13g2_decap_8 FILLER_12_2489 ();
 sg13g2_fill_2 FILLER_12_2496 ();
 sg13g2_decap_8 FILLER_12_2501 ();
 sg13g2_decap_4 FILLER_12_2508 ();
 sg13g2_fill_1 FILLER_12_2512 ();
 sg13g2_decap_8 FILLER_12_2517 ();
 sg13g2_decap_8 FILLER_12_2524 ();
 sg13g2_decap_8 FILLER_12_2531 ();
 sg13g2_decap_8 FILLER_12_2538 ();
 sg13g2_decap_8 FILLER_12_2545 ();
 sg13g2_decap_8 FILLER_12_2552 ();
 sg13g2_decap_8 FILLER_12_2572 ();
 sg13g2_decap_8 FILLER_12_2579 ();
 sg13g2_decap_8 FILLER_12_2586 ();
 sg13g2_decap_8 FILLER_12_2593 ();
 sg13g2_fill_2 FILLER_12_2600 ();
 sg13g2_fill_1 FILLER_12_2602 ();
 sg13g2_decap_8 FILLER_12_2607 ();
 sg13g2_decap_8 FILLER_12_2614 ();
 sg13g2_decap_8 FILLER_12_2621 ();
 sg13g2_decap_8 FILLER_12_2628 ();
 sg13g2_decap_8 FILLER_12_2635 ();
 sg13g2_decap_8 FILLER_12_2642 ();
 sg13g2_decap_8 FILLER_12_2649 ();
 sg13g2_decap_8 FILLER_12_2656 ();
 sg13g2_decap_8 FILLER_12_2663 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_15 ();
 sg13g2_decap_4 FILLER_13_22 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_decap_8 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_decap_4 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_237 ();
 sg13g2_decap_4 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_decap_4 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_decap_4 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_329 ();
 sg13g2_fill_1 FILLER_13_357 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_404 ();
 sg13g2_fill_2 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_4 FILLER_13_481 ();
 sg13g2_decap_4 FILLER_13_573 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_fill_2 FILLER_13_605 ();
 sg13g2_fill_1 FILLER_13_607 ();
 sg13g2_fill_1 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_decap_8 FILLER_13_681 ();
 sg13g2_fill_2 FILLER_13_688 ();
 sg13g2_fill_1 FILLER_13_690 ();
 sg13g2_fill_2 FILLER_13_695 ();
 sg13g2_decap_8 FILLER_13_744 ();
 sg13g2_fill_1 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_4 FILLER_13_784 ();
 sg13g2_fill_1 FILLER_13_788 ();
 sg13g2_fill_2 FILLER_13_815 ();
 sg13g2_fill_1 FILLER_13_817 ();
 sg13g2_fill_2 FILLER_13_823 ();
 sg13g2_fill_2 FILLER_13_864 ();
 sg13g2_decap_8 FILLER_13_937 ();
 sg13g2_decap_8 FILLER_13_944 ();
 sg13g2_decap_4 FILLER_13_951 ();
 sg13g2_fill_1 FILLER_13_955 ();
 sg13g2_decap_4 FILLER_13_1077 ();
 sg13g2_fill_2 FILLER_13_1081 ();
 sg13g2_fill_1 FILLER_13_1087 ();
 sg13g2_fill_1 FILLER_13_1121 ();
 sg13g2_fill_2 FILLER_13_1127 ();
 sg13g2_fill_2 FILLER_13_1154 ();
 sg13g2_fill_1 FILLER_13_1187 ();
 sg13g2_decap_8 FILLER_13_1209 ();
 sg13g2_decap_8 FILLER_13_1216 ();
 sg13g2_decap_8 FILLER_13_1223 ();
 sg13g2_decap_8 FILLER_13_1230 ();
 sg13g2_decap_8 FILLER_13_1237 ();
 sg13g2_fill_2 FILLER_13_1244 ();
 sg13g2_fill_2 FILLER_13_1277 ();
 sg13g2_fill_1 FILLER_13_1279 ();
 sg13g2_decap_8 FILLER_13_1314 ();
 sg13g2_decap_4 FILLER_13_1321 ();
 sg13g2_decap_4 FILLER_13_1346 ();
 sg13g2_fill_1 FILLER_13_1350 ();
 sg13g2_decap_4 FILLER_13_1358 ();
 sg13g2_fill_1 FILLER_13_1392 ();
 sg13g2_decap_8 FILLER_13_1419 ();
 sg13g2_decap_4 FILLER_13_1426 ();
 sg13g2_fill_2 FILLER_13_1430 ();
 sg13g2_fill_1 FILLER_13_1493 ();
 sg13g2_decap_4 FILLER_13_1504 ();
 sg13g2_fill_1 FILLER_13_1508 ();
 sg13g2_decap_4 FILLER_13_1514 ();
 sg13g2_decap_8 FILLER_13_1522 ();
 sg13g2_decap_4 FILLER_13_1529 ();
 sg13g2_fill_1 FILLER_13_1533 ();
 sg13g2_decap_4 FILLER_13_1538 ();
 sg13g2_fill_2 FILLER_13_1542 ();
 sg13g2_fill_2 FILLER_13_1555 ();
 sg13g2_fill_1 FILLER_13_1557 ();
 sg13g2_decap_4 FILLER_13_1562 ();
 sg13g2_fill_2 FILLER_13_1566 ();
 sg13g2_fill_2 FILLER_13_1572 ();
 sg13g2_decap_8 FILLER_13_1595 ();
 sg13g2_decap_4 FILLER_13_1606 ();
 sg13g2_fill_2 FILLER_13_1610 ();
 sg13g2_decap_8 FILLER_13_1622 ();
 sg13g2_decap_8 FILLER_13_1665 ();
 sg13g2_fill_1 FILLER_13_1672 ();
 sg13g2_fill_1 FILLER_13_1710 ();
 sg13g2_fill_1 FILLER_13_1722 ();
 sg13g2_fill_2 FILLER_13_1729 ();
 sg13g2_decap_8 FILLER_13_1752 ();
 sg13g2_decap_4 FILLER_13_1759 ();
 sg13g2_fill_2 FILLER_13_1763 ();
 sg13g2_fill_2 FILLER_13_1769 ();
 sg13g2_fill_1 FILLER_13_1771 ();
 sg13g2_fill_1 FILLER_13_1789 ();
 sg13g2_decap_8 FILLER_13_1824 ();
 sg13g2_decap_8 FILLER_13_1831 ();
 sg13g2_fill_2 FILLER_13_1842 ();
 sg13g2_decap_4 FILLER_13_1848 ();
 sg13g2_decap_4 FILLER_13_1862 ();
 sg13g2_decap_8 FILLER_13_1893 ();
 sg13g2_decap_8 FILLER_13_1900 ();
 sg13g2_decap_4 FILLER_13_1907 ();
 sg13g2_fill_2 FILLER_13_1911 ();
 sg13g2_fill_2 FILLER_13_1977 ();
 sg13g2_fill_1 FILLER_13_1979 ();
 sg13g2_fill_1 FILLER_13_2010 ();
 sg13g2_fill_1 FILLER_13_2047 ();
 sg13g2_fill_2 FILLER_13_2059 ();
 sg13g2_fill_2 FILLER_13_2071 ();
 sg13g2_fill_1 FILLER_13_2083 ();
 sg13g2_fill_1 FILLER_13_2110 ();
 sg13g2_fill_1 FILLER_13_2137 ();
 sg13g2_fill_1 FILLER_13_2142 ();
 sg13g2_fill_1 FILLER_13_2174 ();
 sg13g2_fill_1 FILLER_13_2201 ();
 sg13g2_fill_1 FILLER_13_2238 ();
 sg13g2_fill_2 FILLER_13_2243 ();
 sg13g2_fill_1 FILLER_13_2245 ();
 sg13g2_fill_1 FILLER_13_2250 ();
 sg13g2_decap_4 FILLER_13_2287 ();
 sg13g2_fill_2 FILLER_13_2291 ();
 sg13g2_fill_2 FILLER_13_2314 ();
 sg13g2_decap_8 FILLER_13_2372 ();
 sg13g2_fill_1 FILLER_13_2379 ();
 sg13g2_fill_2 FILLER_13_2405 ();
 sg13g2_fill_2 FILLER_13_2433 ();
 sg13g2_decap_8 FILLER_13_2439 ();
 sg13g2_decap_8 FILLER_13_2446 ();
 sg13g2_decap_4 FILLER_13_2453 ();
 sg13g2_fill_2 FILLER_13_2457 ();
 sg13g2_fill_2 FILLER_13_2504 ();
 sg13g2_decap_8 FILLER_13_2532 ();
 sg13g2_decap_8 FILLER_13_2539 ();
 sg13g2_decap_8 FILLER_13_2552 ();
 sg13g2_fill_2 FILLER_13_2559 ();
 sg13g2_decap_8 FILLER_13_2587 ();
 sg13g2_fill_2 FILLER_13_2594 ();
 sg13g2_decap_8 FILLER_13_2622 ();
 sg13g2_decap_8 FILLER_13_2629 ();
 sg13g2_decap_8 FILLER_13_2636 ();
 sg13g2_decap_8 FILLER_13_2643 ();
 sg13g2_decap_8 FILLER_13_2650 ();
 sg13g2_decap_8 FILLER_13_2657 ();
 sg13g2_decap_4 FILLER_13_2664 ();
 sg13g2_fill_2 FILLER_13_2668 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_44 ();
 sg13g2_decap_8 FILLER_14_50 ();
 sg13g2_fill_1 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_62 ();
 sg13g2_fill_2 FILLER_14_67 ();
 sg13g2_fill_2 FILLER_14_73 ();
 sg13g2_decap_8 FILLER_14_79 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_decap_4 FILLER_14_131 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_decap_4 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_177 ();
 sg13g2_fill_2 FILLER_14_204 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_1 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_decap_4 FILLER_14_305 ();
 sg13g2_fill_2 FILLER_14_309 ();
 sg13g2_fill_2 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_fill_2 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_2 FILLER_14_385 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_439 ();
 sg13g2_decap_4 FILLER_14_446 ();
 sg13g2_fill_1 FILLER_14_450 ();
 sg13g2_fill_2 FILLER_14_460 ();
 sg13g2_fill_1 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_fill_2 FILLER_14_483 ();
 sg13g2_fill_1 FILLER_14_485 ();
 sg13g2_fill_2 FILLER_14_536 ();
 sg13g2_fill_2 FILLER_14_662 ();
 sg13g2_fill_2 FILLER_14_678 ();
 sg13g2_fill_1 FILLER_14_680 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_fill_2 FILLER_14_706 ();
 sg13g2_fill_2 FILLER_14_712 ();
 sg13g2_fill_1 FILLER_14_714 ();
 sg13g2_fill_1 FILLER_14_725 ();
 sg13g2_fill_2 FILLER_14_736 ();
 sg13g2_fill_1 FILLER_14_738 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_782 ();
 sg13g2_fill_1 FILLER_14_789 ();
 sg13g2_fill_1 FILLER_14_826 ();
 sg13g2_fill_1 FILLER_14_867 ();
 sg13g2_fill_1 FILLER_14_872 ();
 sg13g2_decap_4 FILLER_14_907 ();
 sg13g2_decap_4 FILLER_14_919 ();
 sg13g2_fill_2 FILLER_14_923 ();
 sg13g2_decap_8 FILLER_14_929 ();
 sg13g2_fill_1 FILLER_14_936 ();
 sg13g2_fill_1 FILLER_14_940 ();
 sg13g2_fill_2 FILLER_14_945 ();
 sg13g2_decap_8 FILLER_14_951 ();
 sg13g2_fill_2 FILLER_14_958 ();
 sg13g2_fill_1 FILLER_14_960 ();
 sg13g2_decap_8 FILLER_14_991 ();
 sg13g2_decap_4 FILLER_14_998 ();
 sg13g2_fill_2 FILLER_14_1002 ();
 sg13g2_decap_8 FILLER_14_1034 ();
 sg13g2_decap_8 FILLER_14_1041 ();
 sg13g2_decap_4 FILLER_14_1048 ();
 sg13g2_fill_1 FILLER_14_1052 ();
 sg13g2_fill_2 FILLER_14_1111 ();
 sg13g2_fill_1 FILLER_14_1113 ();
 sg13g2_fill_2 FILLER_14_1153 ();
 sg13g2_fill_1 FILLER_14_1155 ();
 sg13g2_fill_2 FILLER_14_1166 ();
 sg13g2_fill_1 FILLER_14_1172 ();
 sg13g2_fill_1 FILLER_14_1177 ();
 sg13g2_fill_1 FILLER_14_1187 ();
 sg13g2_decap_4 FILLER_14_1196 ();
 sg13g2_decap_8 FILLER_14_1204 ();
 sg13g2_decap_4 FILLER_14_1211 ();
 sg13g2_fill_2 FILLER_14_1219 ();
 sg13g2_fill_2 FILLER_14_1225 ();
 sg13g2_fill_1 FILLER_14_1227 ();
 sg13g2_decap_8 FILLER_14_1241 ();
 sg13g2_decap_8 FILLER_14_1248 ();
 sg13g2_decap_8 FILLER_14_1255 ();
 sg13g2_decap_4 FILLER_14_1267 ();
 sg13g2_decap_8 FILLER_14_1357 ();
 sg13g2_fill_2 FILLER_14_1364 ();
 sg13g2_fill_1 FILLER_14_1366 ();
 sg13g2_decap_4 FILLER_14_1379 ();
 sg13g2_fill_2 FILLER_14_1383 ();
 sg13g2_decap_8 FILLER_14_1410 ();
 sg13g2_decap_4 FILLER_14_1417 ();
 sg13g2_fill_2 FILLER_14_1457 ();
 sg13g2_fill_1 FILLER_14_1472 ();
 sg13g2_fill_1 FILLER_14_1480 ();
 sg13g2_fill_1 FILLER_14_1507 ();
 sg13g2_decap_4 FILLER_14_1529 ();
 sg13g2_fill_1 FILLER_14_1533 ();
 sg13g2_decap_4 FILLER_14_1538 ();
 sg13g2_fill_1 FILLER_14_1556 ();
 sg13g2_fill_2 FILLER_14_1567 ();
 sg13g2_fill_2 FILLER_14_1575 ();
 sg13g2_fill_1 FILLER_14_1577 ();
 sg13g2_decap_4 FILLER_14_1583 ();
 sg13g2_fill_1 FILLER_14_1697 ();
 sg13g2_fill_1 FILLER_14_1703 ();
 sg13g2_fill_1 FILLER_14_1708 ();
 sg13g2_fill_2 FILLER_14_1714 ();
 sg13g2_fill_1 FILLER_14_1720 ();
 sg13g2_decap_8 FILLER_14_1725 ();
 sg13g2_decap_4 FILLER_14_1732 ();
 sg13g2_fill_2 FILLER_14_1736 ();
 sg13g2_decap_8 FILLER_14_1742 ();
 sg13g2_decap_8 FILLER_14_1749 ();
 sg13g2_fill_2 FILLER_14_1790 ();
 sg13g2_fill_2 FILLER_14_1796 ();
 sg13g2_fill_2 FILLER_14_1802 ();
 sg13g2_fill_2 FILLER_14_1814 ();
 sg13g2_fill_1 FILLER_14_1816 ();
 sg13g2_decap_4 FILLER_14_1843 ();
 sg13g2_fill_2 FILLER_14_1847 ();
 sg13g2_decap_8 FILLER_14_1885 ();
 sg13g2_decap_8 FILLER_14_1892 ();
 sg13g2_fill_1 FILLER_14_1899 ();
 sg13g2_decap_4 FILLER_14_1910 ();
 sg13g2_fill_1 FILLER_14_1914 ();
 sg13g2_fill_1 FILLER_14_1925 ();
 sg13g2_fill_2 FILLER_14_1947 ();
 sg13g2_fill_1 FILLER_14_1949 ();
 sg13g2_fill_1 FILLER_14_2082 ();
 sg13g2_decap_8 FILLER_14_2152 ();
 sg13g2_decap_4 FILLER_14_2159 ();
 sg13g2_decap_8 FILLER_14_2173 ();
 sg13g2_fill_2 FILLER_14_2180 ();
 sg13g2_decap_4 FILLER_14_2186 ();
 sg13g2_fill_1 FILLER_14_2190 ();
 sg13g2_fill_2 FILLER_14_2201 ();
 sg13g2_fill_2 FILLER_14_2207 ();
 sg13g2_fill_2 FILLER_14_2235 ();
 sg13g2_fill_1 FILLER_14_2331 ();
 sg13g2_decap_8 FILLER_14_2368 ();
 sg13g2_decap_8 FILLER_14_2375 ();
 sg13g2_decap_8 FILLER_14_2382 ();
 sg13g2_decap_8 FILLER_14_2455 ();
 sg13g2_fill_2 FILLER_14_2462 ();
 sg13g2_fill_1 FILLER_14_2464 ();
 sg13g2_fill_1 FILLER_14_2550 ();
 sg13g2_fill_2 FILLER_14_2607 ();
 sg13g2_decap_8 FILLER_14_2635 ();
 sg13g2_decap_8 FILLER_14_2642 ();
 sg13g2_decap_8 FILLER_14_2649 ();
 sg13g2_decap_8 FILLER_14_2656 ();
 sg13g2_decap_8 FILLER_14_2663 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_decap_4 FILLER_15_120 ();
 sg13g2_fill_2 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_fill_1 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_15_415 ();
 sg13g2_decap_4 FILLER_15_429 ();
 sg13g2_fill_1 FILLER_15_433 ();
 sg13g2_decap_4 FILLER_15_444 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_4 FILLER_15_480 ();
 sg13g2_fill_1 FILLER_15_484 ();
 sg13g2_fill_2 FILLER_15_497 ();
 sg13g2_fill_1 FILLER_15_499 ();
 sg13g2_fill_2 FILLER_15_539 ();
 sg13g2_fill_1 FILLER_15_545 ();
 sg13g2_decap_8 FILLER_15_554 ();
 sg13g2_decap_8 FILLER_15_561 ();
 sg13g2_decap_4 FILLER_15_568 ();
 sg13g2_decap_8 FILLER_15_576 ();
 sg13g2_decap_8 FILLER_15_583 ();
 sg13g2_decap_8 FILLER_15_590 ();
 sg13g2_decap_8 FILLER_15_601 ();
 sg13g2_fill_1 FILLER_15_608 ();
 sg13g2_fill_1 FILLER_15_617 ();
 sg13g2_fill_1 FILLER_15_628 ();
 sg13g2_fill_1 FILLER_15_634 ();
 sg13g2_fill_1 FILLER_15_642 ();
 sg13g2_fill_2 FILLER_15_653 ();
 sg13g2_fill_1 FILLER_15_660 ();
 sg13g2_fill_2 FILLER_15_667 ();
 sg13g2_fill_1 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_678 ();
 sg13g2_decap_8 FILLER_15_685 ();
 sg13g2_fill_2 FILLER_15_692 ();
 sg13g2_fill_1 FILLER_15_694 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_fill_1 FILLER_15_749 ();
 sg13g2_fill_1 FILLER_15_780 ();
 sg13g2_fill_1 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_862 ();
 sg13g2_fill_2 FILLER_15_869 ();
 sg13g2_fill_2 FILLER_15_881 ();
 sg13g2_decap_4 FILLER_15_887 ();
 sg13g2_fill_1 FILLER_15_925 ();
 sg13g2_fill_1 FILLER_15_976 ();
 sg13g2_decap_8 FILLER_15_1038 ();
 sg13g2_decap_8 FILLER_15_1045 ();
 sg13g2_decap_4 FILLER_15_1052 ();
 sg13g2_fill_2 FILLER_15_1056 ();
 sg13g2_decap_8 FILLER_15_1067 ();
 sg13g2_fill_2 FILLER_15_1078 ();
 sg13g2_fill_2 FILLER_15_1106 ();
 sg13g2_fill_2 FILLER_15_1146 ();
 sg13g2_fill_1 FILLER_15_1148 ();
 sg13g2_fill_2 FILLER_15_1170 ();
 sg13g2_fill_1 FILLER_15_1172 ();
 sg13g2_decap_4 FILLER_15_1254 ();
 sg13g2_fill_1 FILLER_15_1309 ();
 sg13g2_fill_1 FILLER_15_1318 ();
 sg13g2_fill_1 FILLER_15_1333 ();
 sg13g2_fill_1 FILLER_15_1338 ();
 sg13g2_decap_4 FILLER_15_1360 ();
 sg13g2_fill_1 FILLER_15_1364 ();
 sg13g2_fill_2 FILLER_15_1375 ();
 sg13g2_decap_8 FILLER_15_1412 ();
 sg13g2_decap_8 FILLER_15_1419 ();
 sg13g2_fill_2 FILLER_15_1444 ();
 sg13g2_fill_1 FILLER_15_1446 ();
 sg13g2_fill_1 FILLER_15_1452 ();
 sg13g2_fill_1 FILLER_15_1462 ();
 sg13g2_fill_2 FILLER_15_1468 ();
 sg13g2_fill_1 FILLER_15_1543 ();
 sg13g2_fill_1 FILLER_15_1557 ();
 sg13g2_fill_1 FILLER_15_1573 ();
 sg13g2_fill_2 FILLER_15_1588 ();
 sg13g2_fill_1 FILLER_15_1590 ();
 sg13g2_fill_2 FILLER_15_1596 ();
 sg13g2_fill_1 FILLER_15_1652 ();
 sg13g2_decap_8 FILLER_15_1665 ();
 sg13g2_decap_4 FILLER_15_1672 ();
 sg13g2_fill_1 FILLER_15_1676 ();
 sg13g2_decap_4 FILLER_15_1681 ();
 sg13g2_decap_8 FILLER_15_1690 ();
 sg13g2_decap_4 FILLER_15_1697 ();
 sg13g2_fill_1 FILLER_15_1701 ();
 sg13g2_decap_4 FILLER_15_1752 ();
 sg13g2_fill_1 FILLER_15_1756 ();
 sg13g2_fill_1 FILLER_15_1792 ();
 sg13g2_fill_1 FILLER_15_1797 ();
 sg13g2_fill_2 FILLER_15_1802 ();
 sg13g2_fill_1 FILLER_15_1804 ();
 sg13g2_decap_8 FILLER_15_1835 ();
 sg13g2_fill_2 FILLER_15_1893 ();
 sg13g2_fill_1 FILLER_15_1895 ();
 sg13g2_decap_8 FILLER_15_1922 ();
 sg13g2_fill_1 FILLER_15_1929 ();
 sg13g2_decap_8 FILLER_15_1940 ();
 sg13g2_decap_8 FILLER_15_1951 ();
 sg13g2_fill_1 FILLER_15_1958 ();
 sg13g2_decap_8 FILLER_15_1963 ();
 sg13g2_fill_2 FILLER_15_1970 ();
 sg13g2_fill_2 FILLER_15_1988 ();
 sg13g2_fill_2 FILLER_15_1993 ();
 sg13g2_fill_1 FILLER_15_2015 ();
 sg13g2_fill_2 FILLER_15_2041 ();
 sg13g2_fill_1 FILLER_15_2047 ();
 sg13g2_fill_1 FILLER_15_2111 ();
 sg13g2_decap_8 FILLER_15_2122 ();
 sg13g2_decap_4 FILLER_15_2133 ();
 sg13g2_fill_1 FILLER_15_2137 ();
 sg13g2_decap_8 FILLER_15_2146 ();
 sg13g2_fill_1 FILLER_15_2153 ();
 sg13g2_fill_2 FILLER_15_2175 ();
 sg13g2_fill_1 FILLER_15_2177 ();
 sg13g2_decap_8 FILLER_15_2182 ();
 sg13g2_decap_8 FILLER_15_2189 ();
 sg13g2_fill_2 FILLER_15_2196 ();
 sg13g2_decap_8 FILLER_15_2235 ();
 sg13g2_decap_4 FILLER_15_2242 ();
 sg13g2_fill_1 FILLER_15_2286 ();
 sg13g2_fill_2 FILLER_15_2291 ();
 sg13g2_fill_1 FILLER_15_2293 ();
 sg13g2_fill_2 FILLER_15_2304 ();
 sg13g2_fill_1 FILLER_15_2306 ();
 sg13g2_fill_2 FILLER_15_2310 ();
 sg13g2_fill_1 FILLER_15_2312 ();
 sg13g2_decap_8 FILLER_15_2317 ();
 sg13g2_fill_2 FILLER_15_2328 ();
 sg13g2_fill_1 FILLER_15_2330 ();
 sg13g2_fill_2 FILLER_15_2362 ();
 sg13g2_fill_1 FILLER_15_2364 ();
 sg13g2_decap_8 FILLER_15_2369 ();
 sg13g2_decap_8 FILLER_15_2376 ();
 sg13g2_decap_8 FILLER_15_2383 ();
 sg13g2_decap_4 FILLER_15_2390 ();
 sg13g2_fill_1 FILLER_15_2394 ();
 sg13g2_decap_8 FILLER_15_2405 ();
 sg13g2_decap_4 FILLER_15_2412 ();
 sg13g2_fill_2 FILLER_15_2416 ();
 sg13g2_fill_1 FILLER_15_2474 ();
 sg13g2_fill_1 FILLER_15_2538 ();
 sg13g2_fill_2 FILLER_15_2549 ();
 sg13g2_fill_1 FILLER_15_2581 ();
 sg13g2_fill_1 FILLER_15_2587 ();
 sg13g2_fill_2 FILLER_15_2592 ();
 sg13g2_decap_8 FILLER_15_2629 ();
 sg13g2_decap_8 FILLER_15_2636 ();
 sg13g2_fill_2 FILLER_15_2643 ();
 sg13g2_fill_1 FILLER_15_2645 ();
 sg13g2_decap_8 FILLER_15_2650 ();
 sg13g2_decap_8 FILLER_15_2657 ();
 sg13g2_decap_4 FILLER_15_2664 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_18 ();
 sg13g2_fill_2 FILLER_16_24 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_103 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_301 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_4 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_4 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_436 ();
 sg13g2_fill_2 FILLER_16_463 ();
 sg13g2_fill_1 FILLER_16_491 ();
 sg13g2_fill_1 FILLER_16_496 ();
 sg13g2_fill_2 FILLER_16_505 ();
 sg13g2_fill_2 FILLER_16_512 ();
 sg13g2_fill_1 FILLER_16_514 ();
 sg13g2_fill_2 FILLER_16_523 ();
 sg13g2_decap_8 FILLER_16_556 ();
 sg13g2_fill_2 FILLER_16_589 ();
 sg13g2_fill_1 FILLER_16_591 ();
 sg13g2_decap_8 FILLER_16_596 ();
 sg13g2_fill_2 FILLER_16_603 ();
 sg13g2_fill_1 FILLER_16_605 ();
 sg13g2_decap_4 FILLER_16_621 ();
 sg13g2_fill_2 FILLER_16_625 ();
 sg13g2_fill_2 FILLER_16_631 ();
 sg13g2_fill_1 FILLER_16_638 ();
 sg13g2_fill_2 FILLER_16_643 ();
 sg13g2_fill_1 FILLER_16_655 ();
 sg13g2_fill_2 FILLER_16_661 ();
 sg13g2_fill_1 FILLER_16_663 ();
 sg13g2_decap_4 FILLER_16_668 ();
 sg13g2_decap_4 FILLER_16_676 ();
 sg13g2_fill_2 FILLER_16_720 ();
 sg13g2_fill_1 FILLER_16_722 ();
 sg13g2_fill_1 FILLER_16_857 ();
 sg13g2_fill_2 FILLER_16_872 ();
 sg13g2_fill_1 FILLER_16_874 ();
 sg13g2_decap_8 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_4 FILLER_16_914 ();
 sg13g2_fill_1 FILLER_16_918 ();
 sg13g2_decap_8 FILLER_16_977 ();
 sg13g2_fill_2 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_990 ();
 sg13g2_decap_8 FILLER_16_997 ();
 sg13g2_decap_8 FILLER_16_1004 ();
 sg13g2_decap_8 FILLER_16_1011 ();
 sg13g2_decap_8 FILLER_16_1018 ();
 sg13g2_decap_8 FILLER_16_1025 ();
 sg13g2_decap_4 FILLER_16_1068 ();
 sg13g2_fill_2 FILLER_16_1072 ();
 sg13g2_fill_2 FILLER_16_1095 ();
 sg13g2_fill_1 FILLER_16_1097 ();
 sg13g2_decap_4 FILLER_16_1108 ();
 sg13g2_fill_2 FILLER_16_1112 ();
 sg13g2_fill_2 FILLER_16_1149 ();
 sg13g2_decap_4 FILLER_16_1155 ();
 sg13g2_fill_2 FILLER_16_1159 ();
 sg13g2_fill_1 FILLER_16_1192 ();
 sg13g2_fill_2 FILLER_16_1208 ();
 sg13g2_fill_1 FILLER_16_1210 ();
 sg13g2_fill_1 FILLER_16_1221 ();
 sg13g2_decap_8 FILLER_16_1256 ();
 sg13g2_fill_1 FILLER_16_1286 ();
 sg13g2_fill_2 FILLER_16_1292 ();
 sg13g2_fill_1 FILLER_16_1333 ();
 sg13g2_fill_1 FILLER_16_1365 ();
 sg13g2_fill_1 FILLER_16_1370 ();
 sg13g2_decap_8 FILLER_16_1421 ();
 sg13g2_fill_2 FILLER_16_1428 ();
 sg13g2_fill_1 FILLER_16_1430 ();
 sg13g2_decap_4 FILLER_16_1436 ();
 sg13g2_fill_1 FILLER_16_1440 ();
 sg13g2_fill_2 FILLER_16_1451 ();
 sg13g2_fill_1 FILLER_16_1457 ();
 sg13g2_fill_1 FILLER_16_1474 ();
 sg13g2_fill_2 FILLER_16_1480 ();
 sg13g2_fill_2 FILLER_16_1495 ();
 sg13g2_fill_1 FILLER_16_1497 ();
 sg13g2_decap_4 FILLER_16_1502 ();
 sg13g2_fill_2 FILLER_16_1506 ();
 sg13g2_fill_2 FILLER_16_1512 ();
 sg13g2_fill_1 FILLER_16_1537 ();
 sg13g2_fill_1 FILLER_16_1549 ();
 sg13g2_fill_1 FILLER_16_1567 ();
 sg13g2_fill_2 FILLER_16_1608 ();
 sg13g2_fill_1 FILLER_16_1618 ();
 sg13g2_decap_4 FILLER_16_1623 ();
 sg13g2_fill_1 FILLER_16_1627 ();
 sg13g2_fill_1 FILLER_16_1647 ();
 sg13g2_fill_1 FILLER_16_1652 ();
 sg13g2_fill_1 FILLER_16_1658 ();
 sg13g2_decap_8 FILLER_16_1663 ();
 sg13g2_fill_2 FILLER_16_1670 ();
 sg13g2_fill_1 FILLER_16_1672 ();
 sg13g2_decap_4 FILLER_16_1683 ();
 sg13g2_fill_2 FILLER_16_1687 ();
 sg13g2_decap_8 FILLER_16_1694 ();
 sg13g2_decap_4 FILLER_16_1701 ();
 sg13g2_decap_8 FILLER_16_1740 ();
 sg13g2_decap_8 FILLER_16_1747 ();
 sg13g2_decap_8 FILLER_16_1754 ();
 sg13g2_fill_2 FILLER_16_1761 ();
 sg13g2_decap_4 FILLER_16_1767 ();
 sg13g2_decap_4 FILLER_16_1785 ();
 sg13g2_decap_4 FILLER_16_1809 ();
 sg13g2_fill_2 FILLER_16_1817 ();
 sg13g2_fill_1 FILLER_16_1819 ();
 sg13g2_fill_2 FILLER_16_1924 ();
 sg13g2_fill_2 FILLER_16_1978 ();
 sg13g2_fill_2 FILLER_16_1999 ();
 sg13g2_fill_2 FILLER_16_2026 ();
 sg13g2_fill_2 FILLER_16_2063 ();
 sg13g2_fill_1 FILLER_16_2163 ();
 sg13g2_fill_2 FILLER_16_2168 ();
 sg13g2_fill_2 FILLER_16_2196 ();
 sg13g2_fill_2 FILLER_16_2202 ();
 sg13g2_fill_2 FILLER_16_2233 ();
 sg13g2_fill_1 FILLER_16_2284 ();
 sg13g2_fill_2 FILLER_16_2295 ();
 sg13g2_fill_1 FILLER_16_2297 ();
 sg13g2_fill_2 FILLER_16_2346 ();
 sg13g2_fill_1 FILLER_16_2348 ();
 sg13g2_decap_8 FILLER_16_2389 ();
 sg13g2_decap_8 FILLER_16_2396 ();
 sg13g2_decap_8 FILLER_16_2403 ();
 sg13g2_fill_2 FILLER_16_2410 ();
 sg13g2_fill_1 FILLER_16_2439 ();
 sg13g2_fill_1 FILLER_16_2479 ();
 sg13g2_fill_1 FILLER_16_2549 ();
 sg13g2_fill_1 FILLER_16_2555 ();
 sg13g2_decap_8 FILLER_16_2568 ();
 sg13g2_fill_1 FILLER_16_2575 ();
 sg13g2_decap_4 FILLER_16_2585 ();
 sg13g2_decap_4 FILLER_16_2612 ();
 sg13g2_fill_1 FILLER_16_2621 ();
 sg13g2_fill_1 FILLER_16_2626 ();
 sg13g2_fill_1 FILLER_16_2632 ();
 sg13g2_fill_2 FILLER_16_2637 ();
 sg13g2_decap_4 FILLER_16_2665 ();
 sg13g2_fill_1 FILLER_16_2669 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_32 ();
 sg13g2_fill_2 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_71 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_4 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_2 FILLER_17_101 ();
 sg13g2_decap_4 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_fill_2 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_298 ();
 sg13g2_fill_1 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_decap_4 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_416 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_decap_8 FILLER_17_429 ();
 sg13g2_fill_1 FILLER_17_436 ();
 sg13g2_fill_1 FILLER_17_474 ();
 sg13g2_fill_2 FILLER_17_479 ();
 sg13g2_fill_2 FILLER_17_486 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_decap_4 FILLER_17_495 ();
 sg13g2_fill_2 FILLER_17_507 ();
 sg13g2_fill_1 FILLER_17_509 ();
 sg13g2_decap_8 FILLER_17_524 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_542 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_fill_2 FILLER_17_560 ();
 sg13g2_fill_2 FILLER_17_566 ();
 sg13g2_fill_1 FILLER_17_568 ();
 sg13g2_fill_2 FILLER_17_573 ();
 sg13g2_fill_1 FILLER_17_575 ();
 sg13g2_decap_4 FILLER_17_602 ();
 sg13g2_fill_2 FILLER_17_606 ();
 sg13g2_decap_4 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_628 ();
 sg13g2_fill_2 FILLER_17_639 ();
 sg13g2_fill_1 FILLER_17_641 ();
 sg13g2_fill_2 FILLER_17_646 ();
 sg13g2_fill_1 FILLER_17_652 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_fill_1 FILLER_17_690 ();
 sg13g2_fill_2 FILLER_17_735 ();
 sg13g2_fill_1 FILLER_17_737 ();
 sg13g2_decap_8 FILLER_17_748 ();
 sg13g2_decap_4 FILLER_17_755 ();
 sg13g2_fill_2 FILLER_17_763 ();
 sg13g2_decap_4 FILLER_17_786 ();
 sg13g2_fill_2 FILLER_17_790 ();
 sg13g2_fill_1 FILLER_17_806 ();
 sg13g2_fill_1 FILLER_17_811 ();
 sg13g2_fill_2 FILLER_17_822 ();
 sg13g2_fill_2 FILLER_17_829 ();
 sg13g2_fill_2 FILLER_17_852 ();
 sg13g2_fill_1 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_898 ();
 sg13g2_fill_1 FILLER_17_905 ();
 sg13g2_fill_1 FILLER_17_944 ();
 sg13g2_decap_4 FILLER_17_981 ();
 sg13g2_fill_2 FILLER_17_1034 ();
 sg13g2_decap_8 FILLER_17_1066 ();
 sg13g2_decap_8 FILLER_17_1073 ();
 sg13g2_fill_2 FILLER_17_1080 ();
 sg13g2_fill_1 FILLER_17_1108 ();
 sg13g2_fill_2 FILLER_17_1122 ();
 sg13g2_fill_1 FILLER_17_1124 ();
 sg13g2_decap_4 FILLER_17_1133 ();
 sg13g2_fill_1 FILLER_17_1137 ();
 sg13g2_fill_2 FILLER_17_1143 ();
 sg13g2_fill_1 FILLER_17_1145 ();
 sg13g2_fill_2 FILLER_17_1175 ();
 sg13g2_fill_1 FILLER_17_1177 ();
 sg13g2_fill_1 FILLER_17_1204 ();
 sg13g2_fill_2 FILLER_17_1213 ();
 sg13g2_fill_1 FILLER_17_1228 ();
 sg13g2_fill_1 FILLER_17_1233 ();
 sg13g2_fill_1 FILLER_17_1302 ();
 sg13g2_fill_1 FILLER_17_1329 ();
 sg13g2_fill_2 FILLER_17_1366 ();
 sg13g2_fill_1 FILLER_17_1368 ();
 sg13g2_fill_2 FILLER_17_1395 ();
 sg13g2_fill_2 FILLER_17_1402 ();
 sg13g2_fill_1 FILLER_17_1404 ();
 sg13g2_fill_1 FILLER_17_1431 ();
 sg13g2_fill_1 FILLER_17_1442 ();
 sg13g2_fill_1 FILLER_17_1469 ();
 sg13g2_fill_2 FILLER_17_1475 ();
 sg13g2_decap_8 FILLER_17_1481 ();
 sg13g2_decap_4 FILLER_17_1488 ();
 sg13g2_fill_1 FILLER_17_1492 ();
 sg13g2_decap_4 FILLER_17_1503 ();
 sg13g2_fill_1 FILLER_17_1507 ();
 sg13g2_decap_8 FILLER_17_1513 ();
 sg13g2_fill_2 FILLER_17_1525 ();
 sg13g2_decap_4 FILLER_17_1546 ();
 sg13g2_fill_1 FILLER_17_1558 ();
 sg13g2_fill_1 FILLER_17_1587 ();
 sg13g2_fill_2 FILLER_17_1596 ();
 sg13g2_decap_4 FILLER_17_1606 ();
 sg13g2_fill_2 FILLER_17_1610 ();
 sg13g2_fill_1 FILLER_17_1616 ();
 sg13g2_fill_2 FILLER_17_1622 ();
 sg13g2_fill_2 FILLER_17_1630 ();
 sg13g2_fill_2 FILLER_17_1663 ();
 sg13g2_fill_2 FILLER_17_1699 ();
 sg13g2_fill_1 FILLER_17_1705 ();
 sg13g2_fill_2 FILLER_17_1727 ();
 sg13g2_decap_4 FILLER_17_1735 ();
 sg13g2_fill_1 FILLER_17_1739 ();
 sg13g2_decap_8 FILLER_17_1744 ();
 sg13g2_decap_4 FILLER_17_1751 ();
 sg13g2_fill_1 FILLER_17_1755 ();
 sg13g2_fill_2 FILLER_17_1761 ();
 sg13g2_decap_8 FILLER_17_1768 ();
 sg13g2_decap_8 FILLER_17_1775 ();
 sg13g2_fill_1 FILLER_17_1782 ();
 sg13g2_decap_8 FILLER_17_1788 ();
 sg13g2_fill_2 FILLER_17_1795 ();
 sg13g2_decap_8 FILLER_17_1818 ();
 sg13g2_fill_1 FILLER_17_1825 ();
 sg13g2_decap_8 FILLER_17_1846 ();
 sg13g2_decap_8 FILLER_17_1853 ();
 sg13g2_fill_2 FILLER_17_1860 ();
 sg13g2_decap_8 FILLER_17_1888 ();
 sg13g2_fill_2 FILLER_17_1895 ();
 sg13g2_fill_1 FILLER_17_1897 ();
 sg13g2_fill_2 FILLER_17_1937 ();
 sg13g2_decap_8 FILLER_17_1943 ();
 sg13g2_decap_4 FILLER_17_1950 ();
 sg13g2_fill_2 FILLER_17_1997 ();
 sg13g2_fill_1 FILLER_17_2003 ();
 sg13g2_fill_1 FILLER_17_2043 ();
 sg13g2_decap_4 FILLER_17_2076 ();
 sg13g2_decap_8 FILLER_17_2084 ();
 sg13g2_fill_1 FILLER_17_2091 ();
 sg13g2_fill_1 FILLER_17_2102 ();
 sg13g2_decap_8 FILLER_17_2124 ();
 sg13g2_decap_8 FILLER_17_2131 ();
 sg13g2_decap_8 FILLER_17_2138 ();
 sg13g2_fill_1 FILLER_17_2149 ();
 sg13g2_decap_4 FILLER_17_2184 ();
 sg13g2_fill_2 FILLER_17_2227 ();
 sg13g2_fill_1 FILLER_17_2229 ();
 sg13g2_decap_8 FILLER_17_2256 ();
 sg13g2_fill_2 FILLER_17_2263 ();
 sg13g2_decap_8 FILLER_17_2308 ();
 sg13g2_decap_8 FILLER_17_2315 ();
 sg13g2_decap_8 FILLER_17_2322 ();
 sg13g2_fill_2 FILLER_17_2329 ();
 sg13g2_fill_1 FILLER_17_2331 ();
 sg13g2_decap_4 FILLER_17_2337 ();
 sg13g2_fill_2 FILLER_17_2341 ();
 sg13g2_decap_8 FILLER_17_2347 ();
 sg13g2_decap_8 FILLER_17_2354 ();
 sg13g2_decap_4 FILLER_17_2361 ();
 sg13g2_fill_1 FILLER_17_2365 ();
 sg13g2_fill_1 FILLER_17_2402 ();
 sg13g2_fill_2 FILLER_17_2453 ();
 sg13g2_fill_2 FILLER_17_2510 ();
 sg13g2_fill_2 FILLER_17_2523 ();
 sg13g2_fill_1 FILLER_17_2538 ();
 sg13g2_fill_1 FILLER_17_2550 ();
 sg13g2_fill_2 FILLER_17_2568 ();
 sg13g2_fill_1 FILLER_17_2570 ();
 sg13g2_decap_8 FILLER_17_2589 ();
 sg13g2_decap_4 FILLER_17_2596 ();
 sg13g2_fill_1 FILLER_17_2600 ();
 sg13g2_decap_8 FILLER_17_2627 ();
 sg13g2_fill_1 FILLER_17_2634 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_13 ();
 sg13g2_decap_8 FILLER_18_20 ();
 sg13g2_decap_8 FILLER_18_27 ();
 sg13g2_decap_4 FILLER_18_34 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_decap_8 FILLER_18_44 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_decap_4 FILLER_18_88 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_2 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_282 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_decap_4 FILLER_18_330 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_447 ();
 sg13g2_decap_4 FILLER_18_454 ();
 sg13g2_fill_1 FILLER_18_458 ();
 sg13g2_decap_8 FILLER_18_495 ();
 sg13g2_decap_8 FILLER_18_502 ();
 sg13g2_decap_8 FILLER_18_509 ();
 sg13g2_decap_8 FILLER_18_516 ();
 sg13g2_decap_8 FILLER_18_523 ();
 sg13g2_fill_2 FILLER_18_530 ();
 sg13g2_fill_2 FILLER_18_536 ();
 sg13g2_fill_1 FILLER_18_538 ();
 sg13g2_fill_2 FILLER_18_544 ();
 sg13g2_fill_1 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_591 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_fill_2 FILLER_18_605 ();
 sg13g2_fill_1 FILLER_18_607 ();
 sg13g2_decap_4 FILLER_18_634 ();
 sg13g2_fill_2 FILLER_18_646 ();
 sg13g2_fill_1 FILLER_18_648 ();
 sg13g2_fill_1 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_4 FILLER_18_710 ();
 sg13g2_fill_2 FILLER_18_764 ();
 sg13g2_decap_8 FILLER_18_774 ();
 sg13g2_fill_1 FILLER_18_781 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_4 FILLER_18_822 ();
 sg13g2_fill_2 FILLER_18_826 ();
 sg13g2_decap_4 FILLER_18_831 ();
 sg13g2_fill_2 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_848 ();
 sg13g2_fill_2 FILLER_18_855 ();
 sg13g2_fill_1 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_868 ();
 sg13g2_fill_2 FILLER_18_908 ();
 sg13g2_fill_1 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_968 ();
 sg13g2_fill_1 FILLER_18_975 ();
 sg13g2_fill_2 FILLER_18_988 ();
 sg13g2_fill_2 FILLER_18_1032 ();
 sg13g2_fill_1 FILLER_18_1034 ();
 sg13g2_decap_4 FILLER_18_1039 ();
 sg13g2_fill_1 FILLER_18_1043 ();
 sg13g2_fill_2 FILLER_18_1048 ();
 sg13g2_fill_1 FILLER_18_1050 ();
 sg13g2_decap_4 FILLER_18_1055 ();
 sg13g2_fill_2 FILLER_18_1059 ();
 sg13g2_fill_2 FILLER_18_1102 ();
 sg13g2_decap_4 FILLER_18_1108 ();
 sg13g2_decap_8 FILLER_18_1116 ();
 sg13g2_fill_1 FILLER_18_1123 ();
 sg13g2_decap_8 FILLER_18_1127 ();
 sg13g2_decap_8 FILLER_18_1134 ();
 sg13g2_fill_2 FILLER_18_1141 ();
 sg13g2_decap_4 FILLER_18_1151 ();
 sg13g2_fill_2 FILLER_18_1198 ();
 sg13g2_fill_2 FILLER_18_1221 ();
 sg13g2_fill_1 FILLER_18_1235 ();
 sg13g2_decap_4 FILLER_18_1240 ();
 sg13g2_decap_8 FILLER_18_1248 ();
 sg13g2_fill_1 FILLER_18_1255 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_8 FILLER_18_1267 ();
 sg13g2_decap_4 FILLER_18_1274 ();
 sg13g2_fill_2 FILLER_18_1278 ();
 sg13g2_fill_1 FILLER_18_1309 ();
 sg13g2_fill_2 FILLER_18_1322 ();
 sg13g2_fill_2 FILLER_18_1328 ();
 sg13g2_fill_2 FILLER_18_1390 ();
 sg13g2_fill_1 FILLER_18_1392 ();
 sg13g2_fill_1 FILLER_18_1397 ();
 sg13g2_decap_8 FILLER_18_1419 ();
 sg13g2_fill_1 FILLER_18_1426 ();
 sg13g2_fill_2 FILLER_18_1453 ();
 sg13g2_fill_1 FILLER_18_1455 ();
 sg13g2_fill_2 FILLER_18_1466 ();
 sg13g2_decap_4 FILLER_18_1498 ();
 sg13g2_decap_4 FILLER_18_1507 ();
 sg13g2_decap_4 FILLER_18_1516 ();
 sg13g2_fill_2 FILLER_18_1520 ();
 sg13g2_decap_4 FILLER_18_1525 ();
 sg13g2_decap_4 FILLER_18_1544 ();
 sg13g2_fill_1 FILLER_18_1567 ();
 sg13g2_fill_1 FILLER_18_1582 ();
 sg13g2_fill_2 FILLER_18_1626 ();
 sg13g2_decap_8 FILLER_18_1654 ();
 sg13g2_decap_4 FILLER_18_1661 ();
 sg13g2_fill_1 FILLER_18_1665 ();
 sg13g2_decap_8 FILLER_18_1753 ();
 sg13g2_decap_8 FILLER_18_1760 ();
 sg13g2_decap_4 FILLER_18_1767 ();
 sg13g2_fill_2 FILLER_18_1771 ();
 sg13g2_decap_8 FILLER_18_1787 ();
 sg13g2_decap_8 FILLER_18_1794 ();
 sg13g2_decap_8 FILLER_18_1801 ();
 sg13g2_decap_8 FILLER_18_1808 ();
 sg13g2_fill_2 FILLER_18_1815 ();
 sg13g2_fill_1 FILLER_18_1817 ();
 sg13g2_decap_8 FILLER_18_1840 ();
 sg13g2_decap_8 FILLER_18_1847 ();
 sg13g2_decap_8 FILLER_18_1854 ();
 sg13g2_decap_4 FILLER_18_1861 ();
 sg13g2_fill_1 FILLER_18_1865 ();
 sg13g2_decap_8 FILLER_18_1884 ();
 sg13g2_decap_8 FILLER_18_1891 ();
 sg13g2_fill_2 FILLER_18_1898 ();
 sg13g2_fill_1 FILLER_18_1900 ();
 sg13g2_decap_4 FILLER_18_1906 ();
 sg13g2_decap_4 FILLER_18_1914 ();
 sg13g2_fill_1 FILLER_18_1918 ();
 sg13g2_fill_2 FILLER_18_1923 ();
 sg13g2_fill_1 FILLER_18_1943 ();
 sg13g2_fill_2 FILLER_18_1970 ();
 sg13g2_decap_4 FILLER_18_2039 ();
 sg13g2_fill_1 FILLER_18_2043 ();
 sg13g2_fill_1 FILLER_18_2117 ();
 sg13g2_fill_1 FILLER_18_2148 ();
 sg13g2_fill_2 FILLER_18_2179 ();
 sg13g2_fill_1 FILLER_18_2181 ();
 sg13g2_fill_2 FILLER_18_2324 ();
 sg13g2_decap_8 FILLER_18_2362 ();
 sg13g2_decap_8 FILLER_18_2369 ();
 sg13g2_decap_4 FILLER_18_2376 ();
 sg13g2_fill_2 FILLER_18_2380 ();
 sg13g2_fill_2 FILLER_18_2390 ();
 sg13g2_fill_1 FILLER_18_2428 ();
 sg13g2_fill_2 FILLER_18_2469 ();
 sg13g2_fill_2 FILLER_18_2480 ();
 sg13g2_fill_1 FILLER_18_2487 ();
 sg13g2_fill_1 FILLER_18_2503 ();
 sg13g2_fill_1 FILLER_18_2521 ();
 sg13g2_fill_2 FILLER_18_2552 ();
 sg13g2_fill_1 FILLER_18_2580 ();
 sg13g2_decap_8 FILLER_18_2662 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_29 ();
 sg13g2_decap_8 FILLER_19_36 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_104 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_178 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_fill_2 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_fill_2 FILLER_19_448 ();
 sg13g2_fill_1 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_507 ();
 sg13g2_decap_8 FILLER_19_516 ();
 sg13g2_fill_2 FILLER_19_557 ();
 sg13g2_fill_2 FILLER_19_599 ();
 sg13g2_fill_1 FILLER_19_632 ();
 sg13g2_fill_1 FILLER_19_638 ();
 sg13g2_fill_2 FILLER_19_686 ();
 sg13g2_fill_1 FILLER_19_688 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_fill_1 FILLER_19_735 ();
 sg13g2_fill_2 FILLER_19_787 ();
 sg13g2_fill_1 FILLER_19_793 ();
 sg13g2_decap_8 FILLER_19_820 ();
 sg13g2_fill_1 FILLER_19_827 ();
 sg13g2_fill_2 FILLER_19_838 ();
 sg13g2_fill_1 FILLER_19_840 ();
 sg13g2_fill_2 FILLER_19_919 ();
 sg13g2_fill_1 FILLER_19_935 ();
 sg13g2_fill_2 FILLER_19_942 ();
 sg13g2_fill_2 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_19_1035 ();
 sg13g2_fill_2 FILLER_19_1042 ();
 sg13g2_decap_8 FILLER_19_1070 ();
 sg13g2_decap_4 FILLER_19_1151 ();
 sg13g2_fill_1 FILLER_19_1163 ();
 sg13g2_fill_2 FILLER_19_1191 ();
 sg13g2_fill_1 FILLER_19_1193 ();
 sg13g2_fill_1 FILLER_19_1223 ();
 sg13g2_decap_4 FILLER_19_1268 ();
 sg13g2_fill_1 FILLER_19_1321 ();
 sg13g2_decap_8 FILLER_19_1340 ();
 sg13g2_decap_8 FILLER_19_1347 ();
 sg13g2_decap_4 FILLER_19_1354 ();
 sg13g2_fill_2 FILLER_19_1358 ();
 sg13g2_fill_2 FILLER_19_1374 ();
 sg13g2_fill_1 FILLER_19_1376 ();
 sg13g2_fill_2 FILLER_19_1428 ();
 sg13g2_fill_1 FILLER_19_1430 ();
 sg13g2_fill_2 FILLER_19_1461 ();
 sg13g2_decap_8 FILLER_19_1467 ();
 sg13g2_decap_4 FILLER_19_1474 ();
 sg13g2_fill_1 FILLER_19_1478 ();
 sg13g2_decap_8 FILLER_19_1484 ();
 sg13g2_decap_8 FILLER_19_1491 ();
 sg13g2_fill_2 FILLER_19_1635 ();
 sg13g2_fill_2 FILLER_19_1641 ();
 sg13g2_decap_8 FILLER_19_1647 ();
 sg13g2_decap_4 FILLER_19_1654 ();
 sg13g2_fill_2 FILLER_19_1662 ();
 sg13g2_fill_1 FILLER_19_1679 ();
 sg13g2_fill_1 FILLER_19_1685 ();
 sg13g2_fill_1 FILLER_19_1690 ();
 sg13g2_fill_2 FILLER_19_1697 ();
 sg13g2_fill_1 FILLER_19_1720 ();
 sg13g2_decap_8 FILLER_19_1746 ();
 sg13g2_decap_4 FILLER_19_1753 ();
 sg13g2_fill_1 FILLER_19_1797 ();
 sg13g2_decap_8 FILLER_19_1824 ();
 sg13g2_decap_4 FILLER_19_1857 ();
 sg13g2_fill_1 FILLER_19_1861 ();
 sg13g2_decap_8 FILLER_19_1898 ();
 sg13g2_fill_2 FILLER_19_1905 ();
 sg13g2_fill_1 FILLER_19_1907 ();
 sg13g2_decap_4 FILLER_19_1940 ();
 sg13g2_fill_1 FILLER_19_1949 ();
 sg13g2_fill_2 FILLER_19_1954 ();
 sg13g2_fill_2 FILLER_19_1960 ();
 sg13g2_fill_1 FILLER_19_1962 ();
 sg13g2_fill_2 FILLER_19_1990 ();
 sg13g2_fill_1 FILLER_19_2049 ();
 sg13g2_decap_8 FILLER_19_2060 ();
 sg13g2_fill_1 FILLER_19_2067 ();
 sg13g2_fill_1 FILLER_19_2072 ();
 sg13g2_fill_1 FILLER_19_2109 ();
 sg13g2_fill_1 FILLER_19_2114 ();
 sg13g2_decap_4 FILLER_19_2141 ();
 sg13g2_fill_1 FILLER_19_2168 ();
 sg13g2_fill_1 FILLER_19_2208 ();
 sg13g2_fill_1 FILLER_19_2368 ();
 sg13g2_fill_2 FILLER_19_2373 ();
 sg13g2_fill_1 FILLER_19_2375 ();
 sg13g2_decap_4 FILLER_19_2435 ();
 sg13g2_fill_2 FILLER_19_2453 ();
 sg13g2_fill_1 FILLER_19_2455 ();
 sg13g2_fill_1 FILLER_19_2584 ();
 sg13g2_fill_1 FILLER_19_2590 ();
 sg13g2_fill_2 FILLER_19_2621 ();
 sg13g2_fill_2 FILLER_19_2649 ();
 sg13g2_decap_8 FILLER_19_2655 ();
 sg13g2_decap_8 FILLER_19_2662 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_18 ();
 sg13g2_fill_1 FILLER_20_45 ();
 sg13g2_decap_8 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_90 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_4 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_325 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_decap_4 FILLER_20_344 ();
 sg13g2_decap_4 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_372 ();
 sg13g2_decap_4 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_fill_2 FILLER_20_443 ();
 sg13g2_fill_1 FILLER_20_453 ();
 sg13g2_fill_1 FILLER_20_480 ();
 sg13g2_fill_1 FILLER_20_490 ();
 sg13g2_fill_1 FILLER_20_496 ();
 sg13g2_fill_2 FILLER_20_523 ();
 sg13g2_fill_1 FILLER_20_525 ();
 sg13g2_fill_2 FILLER_20_561 ();
 sg13g2_fill_1 FILLER_20_574 ();
 sg13g2_fill_2 FILLER_20_597 ();
 sg13g2_decap_8 FILLER_20_607 ();
 sg13g2_fill_1 FILLER_20_614 ();
 sg13g2_fill_2 FILLER_20_623 ();
 sg13g2_fill_1 FILLER_20_633 ();
 sg13g2_fill_2 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_8 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_fill_2 FILLER_20_740 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_fill_2 FILLER_20_785 ();
 sg13g2_fill_1 FILLER_20_787 ();
 sg13g2_decap_4 FILLER_20_834 ();
 sg13g2_fill_2 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_fill_2 FILLER_20_876 ();
 sg13g2_decap_8 FILLER_20_904 ();
 sg13g2_fill_2 FILLER_20_911 ();
 sg13g2_fill_1 FILLER_20_913 ();
 sg13g2_fill_2 FILLER_20_963 ();
 sg13g2_fill_2 FILLER_20_979 ();
 sg13g2_decap_4 FILLER_20_1034 ();
 sg13g2_fill_1 FILLER_20_1068 ();
 sg13g2_decap_8 FILLER_20_1108 ();
 sg13g2_decap_8 FILLER_20_1115 ();
 sg13g2_fill_2 FILLER_20_1122 ();
 sg13g2_fill_1 FILLER_20_1127 ();
 sg13g2_decap_8 FILLER_20_1172 ();
 sg13g2_decap_4 FILLER_20_1193 ();
 sg13g2_fill_2 FILLER_20_1257 ();
 sg13g2_fill_2 FILLER_20_1264 ();
 sg13g2_fill_1 FILLER_20_1266 ();
 sg13g2_fill_2 FILLER_20_1293 ();
 sg13g2_fill_2 FILLER_20_1321 ();
 sg13g2_fill_1 FILLER_20_1323 ();
 sg13g2_decap_8 FILLER_20_1360 ();
 sg13g2_decap_8 FILLER_20_1367 ();
 sg13g2_decap_8 FILLER_20_1374 ();
 sg13g2_decap_8 FILLER_20_1381 ();
 sg13g2_fill_2 FILLER_20_1388 ();
 sg13g2_fill_1 FILLER_20_1390 ();
 sg13g2_fill_2 FILLER_20_1396 ();
 sg13g2_decap_4 FILLER_20_1419 ();
 sg13g2_fill_2 FILLER_20_1423 ();
 sg13g2_decap_8 FILLER_20_1435 ();
 sg13g2_decap_8 FILLER_20_1442 ();
 sg13g2_decap_8 FILLER_20_1449 ();
 sg13g2_decap_4 FILLER_20_1456 ();
 sg13g2_fill_1 FILLER_20_1460 ();
 sg13g2_decap_4 FILLER_20_1482 ();
 sg13g2_fill_1 FILLER_20_1486 ();
 sg13g2_decap_4 FILLER_20_1492 ();
 sg13g2_fill_1 FILLER_20_1496 ();
 sg13g2_fill_1 FILLER_20_1500 ();
 sg13g2_decap_8 FILLER_20_1521 ();
 sg13g2_fill_1 FILLER_20_1561 ();
 sg13g2_fill_1 FILLER_20_1587 ();
 sg13g2_fill_2 FILLER_20_1611 ();
 sg13g2_fill_1 FILLER_20_1639 ();
 sg13g2_fill_2 FILLER_20_1643 ();
 sg13g2_decap_8 FILLER_20_1651 ();
 sg13g2_decap_4 FILLER_20_1658 ();
 sg13g2_fill_2 FILLER_20_1662 ();
 sg13g2_fill_2 FILLER_20_1679 ();
 sg13g2_fill_1 FILLER_20_1681 ();
 sg13g2_decap_4 FILLER_20_1708 ();
 sg13g2_decap_8 FILLER_20_1725 ();
 sg13g2_decap_4 FILLER_20_1732 ();
 sg13g2_decap_4 FILLER_20_1744 ();
 sg13g2_fill_1 FILLER_20_1779 ();
 sg13g2_fill_1 FILLER_20_1806 ();
 sg13g2_fill_1 FILLER_20_1817 ();
 sg13g2_decap_4 FILLER_20_1870 ();
 sg13g2_decap_8 FILLER_20_1940 ();
 sg13g2_decap_8 FILLER_20_1947 ();
 sg13g2_decap_8 FILLER_20_1954 ();
 sg13g2_fill_1 FILLER_20_1961 ();
 sg13g2_decap_8 FILLER_20_1966 ();
 sg13g2_decap_8 FILLER_20_1973 ();
 sg13g2_fill_1 FILLER_20_1980 ();
 sg13g2_fill_2 FILLER_20_1994 ();
 sg13g2_fill_1 FILLER_20_2022 ();
 sg13g2_fill_1 FILLER_20_2033 ();
 sg13g2_fill_1 FILLER_20_2096 ();
 sg13g2_decap_8 FILLER_20_2127 ();
 sg13g2_fill_2 FILLER_20_2134 ();
 sg13g2_fill_1 FILLER_20_2136 ();
 sg13g2_fill_2 FILLER_20_2142 ();
 sg13g2_decap_4 FILLER_20_2154 ();
 sg13g2_fill_1 FILLER_20_2162 ();
 sg13g2_fill_2 FILLER_20_2180 ();
 sg13g2_fill_1 FILLER_20_2190 ();
 sg13g2_fill_2 FILLER_20_2251 ();
 sg13g2_fill_2 FILLER_20_2269 ();
 sg13g2_fill_1 FILLER_20_2307 ();
 sg13g2_decap_8 FILLER_20_2344 ();
 sg13g2_decap_8 FILLER_20_2377 ();
 sg13g2_fill_2 FILLER_20_2384 ();
 sg13g2_fill_1 FILLER_20_2463 ();
 sg13g2_decap_8 FILLER_20_2468 ();
 sg13g2_fill_1 FILLER_20_2475 ();
 sg13g2_fill_1 FILLER_20_2512 ();
 sg13g2_fill_1 FILLER_20_2519 ();
 sg13g2_fill_2 FILLER_20_2530 ();
 sg13g2_fill_2 FILLER_20_2537 ();
 sg13g2_fill_1 FILLER_20_2547 ();
 sg13g2_fill_1 FILLER_20_2564 ();
 sg13g2_fill_1 FILLER_20_2595 ();
 sg13g2_fill_2 FILLER_20_2600 ();
 sg13g2_fill_1 FILLER_20_2623 ();
 sg13g2_fill_2 FILLER_20_2633 ();
 sg13g2_decap_8 FILLER_20_2639 ();
 sg13g2_fill_2 FILLER_20_2646 ();
 sg13g2_decap_8 FILLER_20_2652 ();
 sg13g2_decap_8 FILLER_20_2659 ();
 sg13g2_decap_4 FILLER_20_2666 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_fill_2 FILLER_21_65 ();
 sg13g2_fill_1 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_80 ();
 sg13g2_decap_8 FILLER_21_86 ();
 sg13g2_decap_4 FILLER_21_93 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_fill_2 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_299 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_363 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_383 ();
 sg13g2_fill_1 FILLER_21_389 ();
 sg13g2_fill_1 FILLER_21_395 ();
 sg13g2_fill_2 FILLER_21_413 ();
 sg13g2_fill_1 FILLER_21_449 ();
 sg13g2_fill_2 FILLER_21_454 ();
 sg13g2_decap_4 FILLER_21_460 ();
 sg13g2_fill_2 FILLER_21_468 ();
 sg13g2_fill_1 FILLER_21_470 ();
 sg13g2_decap_4 FILLER_21_548 ();
 sg13g2_fill_1 FILLER_21_552 ();
 sg13g2_fill_2 FILLER_21_579 ();
 sg13g2_fill_1 FILLER_21_584 ();
 sg13g2_fill_1 FILLER_21_599 ();
 sg13g2_fill_2 FILLER_21_643 ();
 sg13g2_fill_1 FILLER_21_686 ();
 sg13g2_fill_1 FILLER_21_713 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_fill_2 FILLER_21_732 ();
 sg13g2_fill_2 FILLER_21_744 ();
 sg13g2_fill_1 FILLER_21_750 ();
 sg13g2_fill_2 FILLER_21_777 ();
 sg13g2_fill_2 FILLER_21_820 ();
 sg13g2_fill_1 FILLER_21_825 ();
 sg13g2_fill_2 FILLER_21_840 ();
 sg13g2_decap_4 FILLER_21_868 ();
 sg13g2_fill_2 FILLER_21_882 ();
 sg13g2_fill_1 FILLER_21_884 ();
 sg13g2_fill_2 FILLER_21_889 ();
 sg13g2_fill_1 FILLER_21_938 ();
 sg13g2_fill_1 FILLER_21_955 ();
 sg13g2_fill_2 FILLER_21_1008 ();
 sg13g2_fill_1 FILLER_21_1082 ();
 sg13g2_fill_1 FILLER_21_1107 ();
 sg13g2_fill_2 FILLER_21_1134 ();
 sg13g2_fill_1 FILLER_21_1136 ();
 sg13g2_fill_2 FILLER_21_1166 ();
 sg13g2_decap_8 FILLER_21_1215 ();
 sg13g2_decap_4 FILLER_21_1222 ();
 sg13g2_fill_2 FILLER_21_1278 ();
 sg13g2_fill_1 FILLER_21_1280 ();
 sg13g2_decap_8 FILLER_21_1364 ();
 sg13g2_decap_4 FILLER_21_1371 ();
 sg13g2_fill_1 FILLER_21_1375 ();
 sg13g2_decap_8 FILLER_21_1416 ();
 sg13g2_fill_2 FILLER_21_1431 ();
 sg13g2_decap_4 FILLER_21_1484 ();
 sg13g2_fill_2 FILLER_21_1488 ();
 sg13g2_fill_2 FILLER_21_1528 ();
 sg13g2_fill_2 FILLER_21_1543 ();
 sg13g2_fill_1 FILLER_21_1545 ();
 sg13g2_fill_1 FILLER_21_1555 ();
 sg13g2_fill_1 FILLER_21_1594 ();
 sg13g2_fill_2 FILLER_21_1605 ();
 sg13g2_fill_2 FILLER_21_1613 ();
 sg13g2_fill_1 FILLER_21_1615 ();
 sg13g2_fill_1 FILLER_21_1658 ();
 sg13g2_fill_2 FILLER_21_1675 ();
 sg13g2_decap_4 FILLER_21_1700 ();
 sg13g2_fill_1 FILLER_21_1724 ();
 sg13g2_decap_8 FILLER_21_1730 ();
 sg13g2_decap_8 FILLER_21_1737 ();
 sg13g2_fill_2 FILLER_21_1744 ();
 sg13g2_fill_2 FILLER_21_1755 ();
 sg13g2_fill_1 FILLER_21_1757 ();
 sg13g2_fill_1 FILLER_21_1763 ();
 sg13g2_fill_1 FILLER_21_1778 ();
 sg13g2_fill_1 FILLER_21_1815 ();
 sg13g2_decap_8 FILLER_21_1871 ();
 sg13g2_fill_2 FILLER_21_1878 ();
 sg13g2_decap_4 FILLER_21_1897 ();
 sg13g2_fill_1 FILLER_21_1905 ();
 sg13g2_fill_1 FILLER_21_1916 ();
 sg13g2_decap_8 FILLER_21_1943 ();
 sg13g2_decap_4 FILLER_21_1950 ();
 sg13g2_decap_8 FILLER_21_1958 ();
 sg13g2_decap_8 FILLER_21_2005 ();
 sg13g2_fill_2 FILLER_21_2012 ();
 sg13g2_fill_1 FILLER_21_2082 ();
 sg13g2_decap_8 FILLER_21_2099 ();
 sg13g2_decap_8 FILLER_21_2106 ();
 sg13g2_decap_8 FILLER_21_2113 ();
 sg13g2_decap_8 FILLER_21_2120 ();
 sg13g2_decap_8 FILLER_21_2127 ();
 sg13g2_decap_4 FILLER_21_2134 ();
 sg13g2_fill_2 FILLER_21_2138 ();
 sg13g2_fill_1 FILLER_21_2150 ();
 sg13g2_fill_2 FILLER_21_2161 ();
 sg13g2_fill_1 FILLER_21_2163 ();
 sg13g2_decap_8 FILLER_21_2168 ();
 sg13g2_fill_2 FILLER_21_2175 ();
 sg13g2_decap_8 FILLER_21_2180 ();
 sg13g2_fill_2 FILLER_21_2187 ();
 sg13g2_fill_1 FILLER_21_2202 ();
 sg13g2_decap_8 FILLER_21_2206 ();
 sg13g2_decap_8 FILLER_21_2213 ();
 sg13g2_fill_2 FILLER_21_2286 ();
 sg13g2_fill_2 FILLER_21_2298 ();
 sg13g2_fill_1 FILLER_21_2300 ();
 sg13g2_decap_8 FILLER_21_2311 ();
 sg13g2_decap_8 FILLER_21_2318 ();
 sg13g2_decap_8 FILLER_21_2329 ();
 sg13g2_decap_8 FILLER_21_2336 ();
 sg13g2_fill_1 FILLER_21_2343 ();
 sg13g2_decap_8 FILLER_21_2380 ();
 sg13g2_fill_2 FILLER_21_2387 ();
 sg13g2_fill_1 FILLER_21_2389 ();
 sg13g2_decap_8 FILLER_21_2400 ();
 sg13g2_decap_4 FILLER_21_2417 ();
 sg13g2_fill_2 FILLER_21_2421 ();
 sg13g2_decap_4 FILLER_21_2453 ();
 sg13g2_fill_1 FILLER_21_2457 ();
 sg13g2_decap_4 FILLER_21_2463 ();
 sg13g2_decap_8 FILLER_21_2604 ();
 sg13g2_decap_8 FILLER_21_2611 ();
 sg13g2_decap_8 FILLER_21_2618 ();
 sg13g2_decap_8 FILLER_21_2625 ();
 sg13g2_fill_1 FILLER_21_2632 ();
 sg13g2_fill_2 FILLER_21_2668 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_fill_1 FILLER_22_16 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_45 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_60 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_76 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_decap_4 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_decap_4 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_449 ();
 sg13g2_decap_8 FILLER_22_467 ();
 sg13g2_decap_4 FILLER_22_474 ();
 sg13g2_fill_2 FILLER_22_478 ();
 sg13g2_fill_2 FILLER_22_497 ();
 sg13g2_fill_1 FILLER_22_508 ();
 sg13g2_fill_1 FILLER_22_514 ();
 sg13g2_fill_1 FILLER_22_520 ();
 sg13g2_fill_1 FILLER_22_529 ();
 sg13g2_fill_1 FILLER_22_534 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_4 FILLER_22_550 ();
 sg13g2_fill_2 FILLER_22_589 ();
 sg13g2_fill_2 FILLER_22_596 ();
 sg13g2_fill_1 FILLER_22_598 ();
 sg13g2_decap_4 FILLER_22_607 ();
 sg13g2_fill_2 FILLER_22_670 ();
 sg13g2_fill_2 FILLER_22_680 ();
 sg13g2_fill_1 FILLER_22_689 ();
 sg13g2_fill_1 FILLER_22_694 ();
 sg13g2_fill_1 FILLER_22_700 ();
 sg13g2_fill_2 FILLER_22_705 ();
 sg13g2_decap_4 FILLER_22_733 ();
 sg13g2_fill_1 FILLER_22_737 ();
 sg13g2_fill_1 FILLER_22_768 ();
 sg13g2_fill_2 FILLER_22_779 ();
 sg13g2_fill_2 FILLER_22_785 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_fill_2 FILLER_22_798 ();
 sg13g2_fill_1 FILLER_22_800 ();
 sg13g2_fill_2 FILLER_22_811 ();
 sg13g2_fill_1 FILLER_22_813 ();
 sg13g2_fill_1 FILLER_22_821 ();
 sg13g2_fill_2 FILLER_22_829 ();
 sg13g2_fill_1 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_fill_2 FILLER_22_886 ();
 sg13g2_fill_2 FILLER_22_896 ();
 sg13g2_fill_2 FILLER_22_940 ();
 sg13g2_fill_2 FILLER_22_984 ();
 sg13g2_fill_2 FILLER_22_1058 ();
 sg13g2_fill_2 FILLER_22_1101 ();
 sg13g2_fill_1 FILLER_22_1128 ();
 sg13g2_fill_1 FILLER_22_1155 ();
 sg13g2_fill_2 FILLER_22_1193 ();
 sg13g2_decap_4 FILLER_22_1199 ();
 sg13g2_fill_2 FILLER_22_1203 ();
 sg13g2_decap_8 FILLER_22_1209 ();
 sg13g2_decap_4 FILLER_22_1216 ();
 sg13g2_fill_2 FILLER_22_1220 ();
 sg13g2_decap_4 FILLER_22_1227 ();
 sg13g2_fill_1 FILLER_22_1231 ();
 sg13g2_fill_2 FILLER_22_1240 ();
 sg13g2_fill_1 FILLER_22_1246 ();
 sg13g2_decap_4 FILLER_22_1259 ();
 sg13g2_decap_8 FILLER_22_1267 ();
 sg13g2_decap_8 FILLER_22_1278 ();
 sg13g2_decap_8 FILLER_22_1285 ();
 sg13g2_fill_1 FILLER_22_1292 ();
 sg13g2_fill_2 FILLER_22_1302 ();
 sg13g2_fill_1 FILLER_22_1317 ();
 sg13g2_fill_2 FILLER_22_1322 ();
 sg13g2_fill_1 FILLER_22_1324 ();
 sg13g2_fill_2 FILLER_22_1346 ();
 sg13g2_fill_2 FILLER_22_1374 ();
 sg13g2_fill_1 FILLER_22_1376 ();
 sg13g2_fill_2 FILLER_22_1403 ();
 sg13g2_fill_1 FILLER_22_1405 ();
 sg13g2_fill_2 FILLER_22_1432 ();
 sg13g2_fill_1 FILLER_22_1500 ();
 sg13g2_fill_1 FILLER_22_1631 ();
 sg13g2_fill_1 FILLER_22_1663 ();
 sg13g2_fill_1 FILLER_22_1676 ();
 sg13g2_decap_8 FILLER_22_1737 ();
 sg13g2_fill_2 FILLER_22_1744 ();
 sg13g2_fill_1 FILLER_22_1746 ();
 sg13g2_fill_1 FILLER_22_1751 ();
 sg13g2_fill_1 FILLER_22_1769 ();
 sg13g2_fill_1 FILLER_22_1783 ();
 sg13g2_fill_1 FILLER_22_1810 ();
 sg13g2_fill_2 FILLER_22_1821 ();
 sg13g2_fill_2 FILLER_22_1833 ();
 sg13g2_fill_2 FILLER_22_1839 ();
 sg13g2_fill_2 FILLER_22_1860 ();
 sg13g2_fill_1 FILLER_22_1892 ();
 sg13g2_fill_1 FILLER_22_1903 ();
 sg13g2_decap_4 FILLER_22_1908 ();
 sg13g2_fill_1 FILLER_22_1912 ();
 sg13g2_decap_8 FILLER_22_1949 ();
 sg13g2_decap_4 FILLER_22_1960 ();
 sg13g2_decap_4 FILLER_22_1974 ();
 sg13g2_decap_4 FILLER_22_1982 ();
 sg13g2_fill_2 FILLER_22_1990 ();
 sg13g2_decap_4 FILLER_22_1996 ();
 sg13g2_fill_2 FILLER_22_2004 ();
 sg13g2_fill_1 FILLER_22_2006 ();
 sg13g2_decap_4 FILLER_22_2021 ();
 sg13g2_decap_8 FILLER_22_2033 ();
 sg13g2_fill_2 FILLER_22_2046 ();
 sg13g2_decap_4 FILLER_22_2055 ();
 sg13g2_fill_1 FILLER_22_2092 ();
 sg13g2_decap_8 FILLER_22_2119 ();
 sg13g2_decap_4 FILLER_22_2126 ();
 sg13g2_fill_2 FILLER_22_2130 ();
 sg13g2_fill_2 FILLER_22_2184 ();
 sg13g2_fill_2 FILLER_22_2216 ();
 sg13g2_fill_1 FILLER_22_2218 ();
 sg13g2_fill_1 FILLER_22_2236 ();
 sg13g2_decap_8 FILLER_22_2313 ();
 sg13g2_fill_2 FILLER_22_2320 ();
 sg13g2_decap_4 FILLER_22_2332 ();
 sg13g2_fill_2 FILLER_22_2336 ();
 sg13g2_decap_8 FILLER_22_2342 ();
 sg13g2_decap_8 FILLER_22_2349 ();
 sg13g2_decap_4 FILLER_22_2356 ();
 sg13g2_fill_1 FILLER_22_2360 ();
 sg13g2_decap_8 FILLER_22_2397 ();
 sg13g2_fill_2 FILLER_22_2404 ();
 sg13g2_decap_4 FILLER_22_2429 ();
 sg13g2_fill_1 FILLER_22_2433 ();
 sg13g2_decap_4 FILLER_22_2454 ();
 sg13g2_fill_2 FILLER_22_2458 ();
 sg13g2_fill_2 FILLER_22_2469 ();
 sg13g2_fill_1 FILLER_22_2471 ();
 sg13g2_fill_1 FILLER_22_2481 ();
 sg13g2_fill_2 FILLER_22_2487 ();
 sg13g2_decap_8 FILLER_22_2499 ();
 sg13g2_decap_4 FILLER_22_2506 ();
 sg13g2_fill_1 FILLER_22_2510 ();
 sg13g2_fill_1 FILLER_22_2527 ();
 sg13g2_fill_2 FILLER_22_2533 ();
 sg13g2_fill_1 FILLER_22_2535 ();
 sg13g2_fill_1 FILLER_22_2553 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_64 ();
 sg13g2_fill_1 FILLER_23_66 ();
 sg13g2_fill_1 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_decap_4 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_162 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_2 FILLER_23_192 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_decap_4 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_fill_1 FILLER_23_424 ();
 sg13g2_fill_2 FILLER_23_435 ();
 sg13g2_fill_1 FILLER_23_437 ();
 sg13g2_fill_1 FILLER_23_474 ();
 sg13g2_fill_2 FILLER_23_479 ();
 sg13g2_fill_2 FILLER_23_485 ();
 sg13g2_fill_1 FILLER_23_487 ();
 sg13g2_fill_2 FILLER_23_514 ();
 sg13g2_fill_1 FILLER_23_516 ();
 sg13g2_decap_8 FILLER_23_521 ();
 sg13g2_decap_8 FILLER_23_528 ();
 sg13g2_fill_1 FILLER_23_535 ();
 sg13g2_fill_2 FILLER_23_631 ();
 sg13g2_fill_2 FILLER_23_649 ();
 sg13g2_fill_1 FILLER_23_679 ();
 sg13g2_fill_1 FILLER_23_685 ();
 sg13g2_decap_4 FILLER_23_700 ();
 sg13g2_fill_1 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_fill_1 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_797 ();
 sg13g2_fill_1 FILLER_23_804 ();
 sg13g2_fill_2 FILLER_23_815 ();
 sg13g2_fill_2 FILLER_23_820 ();
 sg13g2_fill_1 FILLER_23_859 ();
 sg13g2_fill_2 FILLER_23_880 ();
 sg13g2_fill_1 FILLER_23_882 ();
 sg13g2_fill_2 FILLER_23_904 ();
 sg13g2_fill_2 FILLER_23_912 ();
 sg13g2_fill_2 FILLER_23_937 ();
 sg13g2_fill_2 FILLER_23_951 ();
 sg13g2_fill_1 FILLER_23_998 ();
 sg13g2_decap_4 FILLER_23_1030 ();
 sg13g2_fill_1 FILLER_23_1034 ();
 sg13g2_fill_2 FILLER_23_1042 ();
 sg13g2_fill_1 FILLER_23_1091 ();
 sg13g2_decap_8 FILLER_23_1095 ();
 sg13g2_decap_8 FILLER_23_1102 ();
 sg13g2_decap_4 FILLER_23_1109 ();
 sg13g2_fill_1 FILLER_23_1113 ();
 sg13g2_fill_2 FILLER_23_1136 ();
 sg13g2_fill_1 FILLER_23_1138 ();
 sg13g2_fill_2 FILLER_23_1160 ();
 sg13g2_fill_1 FILLER_23_1162 ();
 sg13g2_fill_2 FILLER_23_1171 ();
 sg13g2_fill_1 FILLER_23_1173 ();
 sg13g2_fill_2 FILLER_23_1192 ();
 sg13g2_decap_4 FILLER_23_1198 ();
 sg13g2_fill_1 FILLER_23_1207 ();
 sg13g2_fill_1 FILLER_23_1213 ();
 sg13g2_decap_8 FILLER_23_1253 ();
 sg13g2_decap_8 FILLER_23_1265 ();
 sg13g2_decap_8 FILLER_23_1276 ();
 sg13g2_fill_2 FILLER_23_1283 ();
 sg13g2_fill_1 FILLER_23_1285 ();
 sg13g2_fill_2 FILLER_23_1290 ();
 sg13g2_decap_4 FILLER_23_1295 ();
 sg13g2_fill_1 FILLER_23_1299 ();
 sg13g2_decap_8 FILLER_23_1314 ();
 sg13g2_fill_1 FILLER_23_1321 ();
 sg13g2_fill_1 FILLER_23_1340 ();
 sg13g2_fill_2 FILLER_23_1349 ();
 sg13g2_fill_1 FILLER_23_1351 ();
 sg13g2_decap_8 FILLER_23_1356 ();
 sg13g2_decap_8 FILLER_23_1363 ();
 sg13g2_fill_1 FILLER_23_1370 ();
 sg13g2_decap_4 FILLER_23_1379 ();
 sg13g2_decap_4 FILLER_23_1470 ();
 sg13g2_fill_1 FILLER_23_1481 ();
 sg13g2_fill_1 FILLER_23_1496 ();
 sg13g2_fill_1 FILLER_23_1504 ();
 sg13g2_fill_1 FILLER_23_1513 ();
 sg13g2_fill_1 FILLER_23_1548 ();
 sg13g2_fill_1 FILLER_23_1554 ();
 sg13g2_fill_2 FILLER_23_1583 ();
 sg13g2_fill_1 FILLER_23_1625 ();
 sg13g2_fill_2 FILLER_23_1642 ();
 sg13g2_fill_1 FILLER_23_1644 ();
 sg13g2_fill_1 FILLER_23_1652 ();
 sg13g2_fill_2 FILLER_23_1674 ();
 sg13g2_fill_1 FILLER_23_1723 ();
 sg13g2_fill_1 FILLER_23_1729 ();
 sg13g2_fill_1 FILLER_23_1736 ();
 sg13g2_fill_2 FILLER_23_1770 ();
 sg13g2_fill_1 FILLER_23_1772 ();
 sg13g2_fill_2 FILLER_23_1787 ();
 sg13g2_decap_4 FILLER_23_1793 ();
 sg13g2_decap_8 FILLER_23_1807 ();
 sg13g2_decap_4 FILLER_23_1814 ();
 sg13g2_fill_2 FILLER_23_1818 ();
 sg13g2_decap_4 FILLER_23_1824 ();
 sg13g2_fill_1 FILLER_23_1828 ();
 sg13g2_fill_1 FILLER_23_1839 ();
 sg13g2_fill_2 FILLER_23_1846 ();
 sg13g2_fill_2 FILLER_23_1869 ();
 sg13g2_fill_1 FILLER_23_1875 ();
 sg13g2_fill_2 FILLER_23_1931 ();
 sg13g2_fill_1 FILLER_23_1933 ();
 sg13g2_decap_8 FILLER_23_2000 ();
 sg13g2_decap_8 FILLER_23_2043 ();
 sg13g2_decap_4 FILLER_23_2050 ();
 sg13g2_fill_1 FILLER_23_2054 ();
 sg13g2_fill_1 FILLER_23_2063 ();
 sg13g2_decap_8 FILLER_23_2072 ();
 sg13g2_decap_8 FILLER_23_2083 ();
 sg13g2_decap_4 FILLER_23_2090 ();
 sg13g2_fill_1 FILLER_23_2094 ();
 sg13g2_decap_8 FILLER_23_2098 ();
 sg13g2_decap_8 FILLER_23_2105 ();
 sg13g2_fill_1 FILLER_23_2112 ();
 sg13g2_decap_4 FILLER_23_2175 ();
 sg13g2_fill_1 FILLER_23_2179 ();
 sg13g2_fill_1 FILLER_23_2206 ();
 sg13g2_fill_1 FILLER_23_2238 ();
 sg13g2_fill_2 FILLER_23_2302 ();
 sg13g2_fill_1 FILLER_23_2325 ();
 sg13g2_fill_2 FILLER_23_2357 ();
 sg13g2_fill_1 FILLER_23_2359 ();
 sg13g2_decap_8 FILLER_23_2364 ();
 sg13g2_decap_8 FILLER_23_2371 ();
 sg13g2_fill_2 FILLER_23_2382 ();
 sg13g2_fill_1 FILLER_23_2420 ();
 sg13g2_fill_1 FILLER_23_2482 ();
 sg13g2_decap_4 FILLER_23_2489 ();
 sg13g2_fill_2 FILLER_23_2493 ();
 sg13g2_fill_2 FILLER_23_2507 ();
 sg13g2_fill_1 FILLER_23_2516 ();
 sg13g2_fill_1 FILLER_23_2557 ();
 sg13g2_decap_8 FILLER_23_2661 ();
 sg13g2_fill_2 FILLER_23_2668 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_33 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_78 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_decap_4 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_168 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_fill_1 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_decap_4 FILLER_24_381 ();
 sg13g2_fill_1 FILLER_24_385 ();
 sg13g2_fill_2 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_419 ();
 sg13g2_fill_1 FILLER_24_460 ();
 sg13g2_fill_1 FILLER_24_497 ();
 sg13g2_fill_1 FILLER_24_550 ();
 sg13g2_fill_2 FILLER_24_621 ();
 sg13g2_fill_1 FILLER_24_630 ();
 sg13g2_fill_2 FILLER_24_636 ();
 sg13g2_fill_1 FILLER_24_648 ();
 sg13g2_decap_4 FILLER_24_678 ();
 sg13g2_fill_1 FILLER_24_696 ();
 sg13g2_decap_8 FILLER_24_702 ();
 sg13g2_decap_8 FILLER_24_709 ();
 sg13g2_fill_1 FILLER_24_720 ();
 sg13g2_fill_1 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_fill_2 FILLER_24_774 ();
 sg13g2_fill_2 FILLER_24_780 ();
 sg13g2_fill_1 FILLER_24_782 ();
 sg13g2_fill_2 FILLER_24_793 ();
 sg13g2_fill_1 FILLER_24_795 ();
 sg13g2_fill_1 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_24_856 ();
 sg13g2_fill_1 FILLER_24_904 ();
 sg13g2_fill_1 FILLER_24_956 ();
 sg13g2_fill_2 FILLER_24_1032 ();
 sg13g2_fill_1 FILLER_24_1039 ();
 sg13g2_decap_4 FILLER_24_1123 ();
 sg13g2_fill_2 FILLER_24_1136 ();
 sg13g2_fill_2 FILLER_24_1142 ();
 sg13g2_fill_1 FILLER_24_1144 ();
 sg13g2_fill_1 FILLER_24_1174 ();
 sg13g2_fill_1 FILLER_24_1222 ();
 sg13g2_fill_2 FILLER_24_1302 ();
 sg13g2_fill_1 FILLER_24_1307 ();
 sg13g2_fill_1 FILLER_24_1329 ();
 sg13g2_fill_1 FILLER_24_1335 ();
 sg13g2_decap_8 FILLER_24_1362 ();
 sg13g2_decap_8 FILLER_24_1369 ();
 sg13g2_fill_2 FILLER_24_1376 ();
 sg13g2_fill_2 FILLER_24_1387 ();
 sg13g2_fill_1 FILLER_24_1389 ();
 sg13g2_fill_2 FILLER_24_1400 ();
 sg13g2_fill_1 FILLER_24_1402 ();
 sg13g2_decap_8 FILLER_24_1429 ();
 sg13g2_fill_2 FILLER_24_1436 ();
 sg13g2_fill_1 FILLER_24_1476 ();
 sg13g2_fill_2 FILLER_24_1485 ();
 sg13g2_fill_2 FILLER_24_1495 ();
 sg13g2_fill_2 FILLER_24_1504 ();
 sg13g2_fill_2 FILLER_24_1526 ();
 sg13g2_decap_4 FILLER_24_1563 ();
 sg13g2_fill_1 FILLER_24_1567 ();
 sg13g2_fill_2 FILLER_24_1575 ();
 sg13g2_fill_2 FILLER_24_1595 ();
 sg13g2_fill_1 FILLER_24_1602 ();
 sg13g2_fill_2 FILLER_24_1611 ();
 sg13g2_fill_1 FILLER_24_1613 ();
 sg13g2_fill_1 FILLER_24_1645 ();
 sg13g2_decap_4 FILLER_24_1660 ();
 sg13g2_fill_1 FILLER_24_1736 ();
 sg13g2_fill_1 FILLER_24_1742 ();
 sg13g2_fill_1 FILLER_24_1769 ();
 sg13g2_fill_1 FILLER_24_1780 ();
 sg13g2_fill_1 FILLER_24_1785 ();
 sg13g2_fill_1 FILLER_24_1811 ();
 sg13g2_decap_4 FILLER_24_1822 ();
 sg13g2_fill_2 FILLER_24_1826 ();
 sg13g2_decap_4 FILLER_24_1832 ();
 sg13g2_fill_1 FILLER_24_1836 ();
 sg13g2_fill_2 FILLER_24_1879 ();
 sg13g2_fill_1 FILLER_24_1881 ();
 sg13g2_decap_8 FILLER_24_1918 ();
 sg13g2_decap_4 FILLER_24_1925 ();
 sg13g2_decap_8 FILLER_24_1933 ();
 sg13g2_decap_4 FILLER_24_1940 ();
 sg13g2_fill_2 FILLER_24_1944 ();
 sg13g2_fill_2 FILLER_24_1960 ();
 sg13g2_fill_1 FILLER_24_1983 ();
 sg13g2_decap_8 FILLER_24_2010 ();
 sg13g2_fill_1 FILLER_24_2017 ();
 sg13g2_fill_2 FILLER_24_2038 ();
 sg13g2_fill_1 FILLER_24_2040 ();
 sg13g2_fill_1 FILLER_24_2051 ();
 sg13g2_fill_1 FILLER_24_2104 ();
 sg13g2_decap_8 FILLER_24_2113 ();
 sg13g2_decap_4 FILLER_24_2120 ();
 sg13g2_fill_1 FILLER_24_2124 ();
 sg13g2_decap_4 FILLER_24_2134 ();
 sg13g2_fill_1 FILLER_24_2138 ();
 sg13g2_fill_1 FILLER_24_2143 ();
 sg13g2_fill_1 FILLER_24_2165 ();
 sg13g2_fill_2 FILLER_24_2223 ();
 sg13g2_fill_1 FILLER_24_2225 ();
 sg13g2_fill_1 FILLER_24_2248 ();
 sg13g2_fill_2 FILLER_24_2274 ();
 sg13g2_fill_1 FILLER_24_2276 ();
 sg13g2_fill_2 FILLER_24_2303 ();
 sg13g2_fill_1 FILLER_24_2326 ();
 sg13g2_fill_1 FILLER_24_2384 ();
 sg13g2_decap_8 FILLER_24_2427 ();
 sg13g2_decap_8 FILLER_24_2434 ();
 sg13g2_decap_8 FILLER_24_2453 ();
 sg13g2_decap_4 FILLER_24_2464 ();
 sg13g2_fill_2 FILLER_24_2473 ();
 sg13g2_fill_2 FILLER_24_2481 ();
 sg13g2_fill_1 FILLER_24_2483 ();
 sg13g2_fill_2 FILLER_24_2488 ();
 sg13g2_fill_1 FILLER_24_2537 ();
 sg13g2_fill_1 FILLER_24_2546 ();
 sg13g2_fill_2 FILLER_24_2578 ();
 sg13g2_fill_1 FILLER_24_2593 ();
 sg13g2_fill_2 FILLER_24_2603 ();
 sg13g2_fill_1 FILLER_24_2622 ();
 sg13g2_fill_1 FILLER_24_2629 ();
 sg13g2_fill_1 FILLER_24_2637 ();
 sg13g2_decap_8 FILLER_24_2645 ();
 sg13g2_decap_8 FILLER_24_2652 ();
 sg13g2_decap_8 FILLER_24_2659 ();
 sg13g2_decap_4 FILLER_24_2666 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_33 ();
 sg13g2_fill_2 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_fill_1 FILLER_25_96 ();
 sg13g2_decap_4 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_312 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_fill_1 FILLER_25_430 ();
 sg13g2_decap_8 FILLER_25_435 ();
 sg13g2_decap_8 FILLER_25_442 ();
 sg13g2_decap_8 FILLER_25_449 ();
 sg13g2_fill_1 FILLER_25_461 ();
 sg13g2_fill_1 FILLER_25_479 ();
 sg13g2_decap_8 FILLER_25_484 ();
 sg13g2_fill_2 FILLER_25_491 ();
 sg13g2_fill_1 FILLER_25_497 ();
 sg13g2_fill_1 FILLER_25_502 ();
 sg13g2_fill_1 FILLER_25_507 ();
 sg13g2_fill_1 FILLER_25_512 ();
 sg13g2_fill_2 FILLER_25_518 ();
 sg13g2_fill_2 FILLER_25_565 ();
 sg13g2_fill_2 FILLER_25_575 ();
 sg13g2_fill_2 FILLER_25_594 ();
 sg13g2_fill_1 FILLER_25_631 ();
 sg13g2_fill_2 FILLER_25_635 ();
 sg13g2_fill_1 FILLER_25_647 ();
 sg13g2_fill_1 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_678 ();
 sg13g2_fill_1 FILLER_25_685 ();
 sg13g2_fill_2 FILLER_25_693 ();
 sg13g2_fill_1 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_4 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_796 ();
 sg13g2_fill_1 FILLER_25_856 ();
 sg13g2_fill_1 FILLER_25_909 ();
 sg13g2_fill_1 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_1005 ();
 sg13g2_decap_4 FILLER_25_1012 ();
 sg13g2_fill_2 FILLER_25_1026 ();
 sg13g2_fill_1 FILLER_25_1033 ();
 sg13g2_fill_1 FILLER_25_1039 ();
 sg13g2_decap_4 FILLER_25_1047 ();
 sg13g2_fill_1 FILLER_25_1051 ();
 sg13g2_fill_2 FILLER_25_1075 ();
 sg13g2_fill_1 FILLER_25_1103 ();
 sg13g2_fill_2 FILLER_25_1114 ();
 sg13g2_fill_2 FILLER_25_1175 ();
 sg13g2_fill_2 FILLER_25_1203 ();
 sg13g2_fill_2 FILLER_25_1209 ();
 sg13g2_fill_2 FILLER_25_1215 ();
 sg13g2_fill_1 FILLER_25_1217 ();
 sg13g2_fill_2 FILLER_25_1290 ();
 sg13g2_fill_1 FILLER_25_1326 ();
 sg13g2_fill_1 FILLER_25_1337 ();
 sg13g2_fill_1 FILLER_25_1342 ();
 sg13g2_fill_2 FILLER_25_1369 ();
 sg13g2_fill_2 FILLER_25_1385 ();
 sg13g2_fill_2 FILLER_25_1418 ();
 sg13g2_fill_1 FILLER_25_1420 ();
 sg13g2_fill_1 FILLER_25_1488 ();
 sg13g2_fill_1 FILLER_25_1497 ();
 sg13g2_fill_1 FILLER_25_1531 ();
 sg13g2_decap_8 FILLER_25_1552 ();
 sg13g2_decap_8 FILLER_25_1559 ();
 sg13g2_decap_8 FILLER_25_1566 ();
 sg13g2_fill_1 FILLER_25_1590 ();
 sg13g2_fill_1 FILLER_25_1596 ();
 sg13g2_fill_2 FILLER_25_1605 ();
 sg13g2_decap_4 FILLER_25_1645 ();
 sg13g2_decap_4 FILLER_25_1686 ();
 sg13g2_fill_1 FILLER_25_1720 ();
 sg13g2_fill_2 FILLER_25_1725 ();
 sg13g2_fill_1 FILLER_25_1746 ();
 sg13g2_fill_1 FILLER_25_1756 ();
 sg13g2_fill_1 FILLER_25_1762 ();
 sg13g2_decap_4 FILLER_25_1776 ();
 sg13g2_fill_1 FILLER_25_1780 ();
 sg13g2_fill_1 FILLER_25_1807 ();
 sg13g2_fill_1 FILLER_25_1818 ();
 sg13g2_fill_2 FILLER_25_1845 ();
 sg13g2_fill_2 FILLER_25_1894 ();
 sg13g2_fill_1 FILLER_25_1931 ();
 sg13g2_decap_8 FILLER_25_1957 ();
 sg13g2_decap_4 FILLER_25_1964 ();
 sg13g2_fill_1 FILLER_25_1968 ();
 sg13g2_fill_1 FILLER_25_2007 ();
 sg13g2_fill_1 FILLER_25_2017 ();
 sg13g2_fill_1 FILLER_25_2028 ();
 sg13g2_fill_1 FILLER_25_2065 ();
 sg13g2_fill_2 FILLER_25_2128 ();
 sg13g2_decap_8 FILLER_25_2134 ();
 sg13g2_decap_4 FILLER_25_2141 ();
 sg13g2_fill_1 FILLER_25_2145 ();
 sg13g2_fill_2 FILLER_25_2160 ();
 sg13g2_fill_2 FILLER_25_2300 ();
 sg13g2_fill_1 FILLER_25_2333 ();
 sg13g2_decap_8 FILLER_25_2374 ();
 sg13g2_decap_8 FILLER_25_2381 ();
 sg13g2_decap_8 FILLER_25_2388 ();
 sg13g2_decap_8 FILLER_25_2395 ();
 sg13g2_fill_1 FILLER_25_2402 ();
 sg13g2_decap_4 FILLER_25_2413 ();
 sg13g2_fill_1 FILLER_25_2417 ();
 sg13g2_decap_8 FILLER_25_2448 ();
 sg13g2_fill_1 FILLER_25_2455 ();
 sg13g2_fill_2 FILLER_25_2461 ();
 sg13g2_fill_2 FILLER_25_2468 ();
 sg13g2_decap_4 FILLER_25_2507 ();
 sg13g2_fill_1 FILLER_25_2511 ();
 sg13g2_fill_2 FILLER_25_2518 ();
 sg13g2_fill_1 FILLER_25_2520 ();
 sg13g2_fill_1 FILLER_25_2565 ();
 sg13g2_fill_2 FILLER_25_2605 ();
 sg13g2_fill_2 FILLER_25_2642 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_114 ();
 sg13g2_decap_4 FILLER_26_121 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_decap_8 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_decap_4 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_396 ();
 sg13g2_fill_1 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_428 ();
 sg13g2_fill_1 FILLER_26_440 ();
 sg13g2_decap_8 FILLER_26_450 ();
 sg13g2_decap_8 FILLER_26_457 ();
 sg13g2_fill_1 FILLER_26_464 ();
 sg13g2_decap_4 FILLER_26_473 ();
 sg13g2_fill_2 FILLER_26_477 ();
 sg13g2_decap_8 FILLER_26_514 ();
 sg13g2_fill_2 FILLER_26_552 ();
 sg13g2_fill_2 FILLER_26_558 ();
 sg13g2_fill_2 FILLER_26_569 ();
 sg13g2_fill_2 FILLER_26_658 ();
 sg13g2_decap_4 FILLER_26_677 ();
 sg13g2_fill_2 FILLER_26_681 ();
 sg13g2_fill_2 FILLER_26_695 ();
 sg13g2_fill_1 FILLER_26_697 ();
 sg13g2_fill_2 FILLER_26_729 ();
 sg13g2_fill_2 FILLER_26_761 ();
 sg13g2_fill_2 FILLER_26_814 ();
 sg13g2_fill_1 FILLER_26_816 ();
 sg13g2_fill_2 FILLER_26_827 ();
 sg13g2_fill_2 FILLER_26_842 ();
 sg13g2_fill_1 FILLER_26_870 ();
 sg13g2_fill_2 FILLER_26_901 ();
 sg13g2_fill_2 FILLER_26_932 ();
 sg13g2_fill_1 FILLER_26_964 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_fill_2 FILLER_26_1029 ();
 sg13g2_fill_2 FILLER_26_1042 ();
 sg13g2_fill_2 FILLER_26_1047 ();
 sg13g2_decap_8 FILLER_26_1062 ();
 sg13g2_fill_2 FILLER_26_1069 ();
 sg13g2_decap_8 FILLER_26_1075 ();
 sg13g2_fill_1 FILLER_26_1082 ();
 sg13g2_decap_8 FILLER_26_1198 ();
 sg13g2_decap_8 FILLER_26_1205 ();
 sg13g2_fill_2 FILLER_26_1242 ();
 sg13g2_fill_1 FILLER_26_1244 ();
 sg13g2_decap_4 FILLER_26_1249 ();
 sg13g2_fill_1 FILLER_26_1284 ();
 sg13g2_decap_4 FILLER_26_1345 ();
 sg13g2_fill_2 FILLER_26_1349 ();
 sg13g2_decap_8 FILLER_26_1355 ();
 sg13g2_fill_2 FILLER_26_1392 ();
 sg13g2_decap_8 FILLER_26_1398 ();
 sg13g2_fill_1 FILLER_26_1405 ();
 sg13g2_fill_2 FILLER_26_1439 ();
 sg13g2_fill_2 FILLER_26_1446 ();
 sg13g2_fill_2 FILLER_26_1481 ();
 sg13g2_decap_4 FILLER_26_1560 ();
 sg13g2_fill_1 FILLER_26_1564 ();
 sg13g2_fill_1 FILLER_26_1584 ();
 sg13g2_fill_1 FILLER_26_1608 ();
 sg13g2_fill_1 FILLER_26_1639 ();
 sg13g2_decap_8 FILLER_26_1644 ();
 sg13g2_decap_4 FILLER_26_1651 ();
 sg13g2_fill_1 FILLER_26_1655 ();
 sg13g2_decap_8 FILLER_26_1661 ();
 sg13g2_decap_4 FILLER_26_1668 ();
 sg13g2_fill_2 FILLER_26_1672 ();
 sg13g2_decap_8 FILLER_26_1679 ();
 sg13g2_decap_8 FILLER_26_1686 ();
 sg13g2_decap_4 FILLER_26_1693 ();
 sg13g2_fill_1 FILLER_26_1697 ();
 sg13g2_fill_2 FILLER_26_1719 ();
 sg13g2_fill_1 FILLER_26_1721 ();
 sg13g2_fill_1 FILLER_26_1734 ();
 sg13g2_fill_1 FILLER_26_1751 ();
 sg13g2_decap_4 FILLER_26_1760 ();
 sg13g2_fill_2 FILLER_26_1774 ();
 sg13g2_decap_8 FILLER_26_1794 ();
 sg13g2_fill_1 FILLER_26_1801 ();
 sg13g2_fill_1 FILLER_26_1852 ();
 sg13g2_fill_1 FILLER_26_1857 ();
 sg13g2_decap_8 FILLER_26_1884 ();
 sg13g2_fill_2 FILLER_26_1891 ();
 sg13g2_fill_1 FILLER_26_1893 ();
 sg13g2_fill_2 FILLER_26_1904 ();
 sg13g2_decap_8 FILLER_26_1937 ();
 sg13g2_fill_2 FILLER_26_1944 ();
 sg13g2_fill_1 FILLER_26_1946 ();
 sg13g2_fill_1 FILLER_26_1951 ();
 sg13g2_fill_1 FILLER_26_1961 ();
 sg13g2_fill_2 FILLER_26_1970 ();
 sg13g2_fill_2 FILLER_26_2054 ();
 sg13g2_fill_1 FILLER_26_2056 ();
 sg13g2_fill_2 FILLER_26_2093 ();
 sg13g2_decap_4 FILLER_26_2129 ();
 sg13g2_decap_4 FILLER_26_2138 ();
 sg13g2_fill_2 FILLER_26_2150 ();
 sg13g2_fill_1 FILLER_26_2152 ();
 sg13g2_decap_4 FILLER_26_2163 ();
 sg13g2_fill_2 FILLER_26_2167 ();
 sg13g2_fill_2 FILLER_26_2180 ();
 sg13g2_fill_2 FILLER_26_2190 ();
 sg13g2_fill_2 FILLER_26_2207 ();
 sg13g2_fill_1 FILLER_26_2249 ();
 sg13g2_decap_8 FILLER_26_2273 ();
 sg13g2_decap_4 FILLER_26_2280 ();
 sg13g2_fill_2 FILLER_26_2287 ();
 sg13g2_fill_1 FILLER_26_2289 ();
 sg13g2_fill_2 FILLER_26_2294 ();
 sg13g2_decap_8 FILLER_26_2304 ();
 sg13g2_fill_2 FILLER_26_2311 ();
 sg13g2_decap_8 FILLER_26_2317 ();
 sg13g2_decap_8 FILLER_26_2324 ();
 sg13g2_decap_8 FILLER_26_2331 ();
 sg13g2_decap_8 FILLER_26_2338 ();
 sg13g2_decap_4 FILLER_26_2345 ();
 sg13g2_fill_1 FILLER_26_2349 ();
 sg13g2_decap_8 FILLER_26_2355 ();
 sg13g2_decap_8 FILLER_26_2362 ();
 sg13g2_decap_8 FILLER_26_2369 ();
 sg13g2_decap_8 FILLER_26_2376 ();
 sg13g2_decap_4 FILLER_26_2383 ();
 sg13g2_fill_2 FILLER_26_2387 ();
 sg13g2_fill_2 FILLER_26_2397 ();
 sg13g2_fill_2 FILLER_26_2404 ();
 sg13g2_fill_1 FILLER_26_2406 ();
 sg13g2_fill_2 FILLER_26_2433 ();
 sg13g2_fill_1 FILLER_26_2435 ();
 sg13g2_decap_8 FILLER_26_2449 ();
 sg13g2_decap_4 FILLER_26_2456 ();
 sg13g2_decap_4 FILLER_26_2465 ();
 sg13g2_fill_2 FILLER_26_2473 ();
 sg13g2_fill_1 FILLER_26_2506 ();
 sg13g2_fill_1 FILLER_26_2520 ();
 sg13g2_fill_1 FILLER_26_2529 ();
 sg13g2_fill_1 FILLER_26_2553 ();
 sg13g2_fill_2 FILLER_26_2575 ();
 sg13g2_fill_1 FILLER_26_2632 ();
 sg13g2_fill_2 FILLER_26_2667 ();
 sg13g2_fill_1 FILLER_26_2669 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_68 ();
 sg13g2_decap_4 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_decap_4 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_4 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_27_442 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_fill_1 FILLER_27_462 ();
 sg13g2_fill_2 FILLER_27_520 ();
 sg13g2_fill_1 FILLER_27_522 ();
 sg13g2_fill_1 FILLER_27_532 ();
 sg13g2_fill_1 FILLER_27_537 ();
 sg13g2_fill_1 FILLER_27_549 ();
 sg13g2_fill_2 FILLER_27_595 ();
 sg13g2_fill_1 FILLER_27_597 ();
 sg13g2_fill_2 FILLER_27_606 ();
 sg13g2_fill_2 FILLER_27_621 ();
 sg13g2_fill_2 FILLER_27_627 ();
 sg13g2_fill_2 FILLER_27_635 ();
 sg13g2_decap_4 FILLER_27_663 ();
 sg13g2_fill_2 FILLER_27_667 ();
 sg13g2_decap_4 FILLER_27_679 ();
 sg13g2_fill_2 FILLER_27_683 ();
 sg13g2_decap_8 FILLER_27_690 ();
 sg13g2_fill_2 FILLER_27_697 ();
 sg13g2_fill_1 FILLER_27_699 ();
 sg13g2_fill_2 FILLER_27_726 ();
 sg13g2_fill_1 FILLER_27_728 ();
 sg13g2_fill_2 FILLER_27_736 ();
 sg13g2_fill_1 FILLER_27_742 ();
 sg13g2_fill_1 FILLER_27_797 ();
 sg13g2_fill_2 FILLER_27_808 ();
 sg13g2_fill_1 FILLER_27_853 ();
 sg13g2_fill_1 FILLER_27_884 ();
 sg13g2_fill_1 FILLER_27_889 ();
 sg13g2_fill_1 FILLER_27_900 ();
 sg13g2_fill_1 FILLER_27_933 ();
 sg13g2_fill_2 FILLER_27_1024 ();
 sg13g2_fill_2 FILLER_27_1029 ();
 sg13g2_fill_1 FILLER_27_1031 ();
 sg13g2_fill_2 FILLER_27_1099 ();
 sg13g2_fill_1 FILLER_27_1122 ();
 sg13g2_fill_1 FILLER_27_1127 ();
 sg13g2_fill_1 FILLER_27_1154 ();
 sg13g2_fill_2 FILLER_27_1163 ();
 sg13g2_fill_2 FILLER_27_1191 ();
 sg13g2_fill_2 FILLER_27_1198 ();
 sg13g2_decap_4 FILLER_27_1204 ();
 sg13g2_fill_2 FILLER_27_1212 ();
 sg13g2_fill_2 FILLER_27_1219 ();
 sg13g2_decap_4 FILLER_27_1225 ();
 sg13g2_fill_1 FILLER_27_1233 ();
 sg13g2_decap_4 FILLER_27_1238 ();
 sg13g2_fill_1 FILLER_27_1246 ();
 sg13g2_fill_1 FILLER_27_1298 ();
 sg13g2_decap_8 FILLER_27_1304 ();
 sg13g2_fill_1 FILLER_27_1311 ();
 sg13g2_decap_8 FILLER_27_1342 ();
 sg13g2_decap_8 FILLER_27_1349 ();
 sg13g2_decap_4 FILLER_27_1356 ();
 sg13g2_fill_1 FILLER_27_1360 ();
 sg13g2_fill_1 FILLER_27_1384 ();
 sg13g2_fill_2 FILLER_27_1411 ();
 sg13g2_fill_1 FILLER_27_1423 ();
 sg13g2_fill_2 FILLER_27_1439 ();
 sg13g2_fill_1 FILLER_27_1496 ();
 sg13g2_fill_1 FILLER_27_1505 ();
 sg13g2_fill_1 FILLER_27_1521 ();
 sg13g2_fill_2 FILLER_27_1548 ();
 sg13g2_fill_2 FILLER_27_1555 ();
 sg13g2_fill_1 FILLER_27_1557 ();
 sg13g2_fill_2 FILLER_27_1563 ();
 sg13g2_fill_1 FILLER_27_1565 ();
 sg13g2_decap_8 FILLER_27_1571 ();
 sg13g2_fill_2 FILLER_27_1578 ();
 sg13g2_fill_1 FILLER_27_1580 ();
 sg13g2_fill_1 FILLER_27_1585 ();
 sg13g2_decap_8 FILLER_27_1590 ();
 sg13g2_fill_2 FILLER_27_1600 ();
 sg13g2_fill_1 FILLER_27_1602 ();
 sg13g2_fill_2 FILLER_27_1633 ();
 sg13g2_fill_1 FILLER_27_1635 ();
 sg13g2_fill_2 FILLER_27_1649 ();
 sg13g2_fill_1 FILLER_27_1651 ();
 sg13g2_decap_8 FILLER_27_1660 ();
 sg13g2_decap_8 FILLER_27_1667 ();
 sg13g2_decap_4 FILLER_27_1678 ();
 sg13g2_fill_1 FILLER_27_1682 ();
 sg13g2_decap_8 FILLER_27_1709 ();
 sg13g2_decap_8 FILLER_27_1716 ();
 sg13g2_decap_8 FILLER_27_1723 ();
 sg13g2_fill_2 FILLER_27_1730 ();
 sg13g2_fill_2 FILLER_27_1739 ();
 sg13g2_fill_1 FILLER_27_1741 ();
 sg13g2_decap_8 FILLER_27_1784 ();
 sg13g2_decap_8 FILLER_27_1791 ();
 sg13g2_decap_8 FILLER_27_1798 ();
 sg13g2_decap_4 FILLER_27_1809 ();
 sg13g2_fill_2 FILLER_27_1818 ();
 sg13g2_decap_8 FILLER_27_1875 ();
 sg13g2_fill_2 FILLER_27_1882 ();
 sg13g2_fill_2 FILLER_27_1914 ();
 sg13g2_fill_2 FILLER_27_1920 ();
 sg13g2_decap_8 FILLER_27_1957 ();
 sg13g2_decap_8 FILLER_27_1964 ();
 sg13g2_fill_1 FILLER_27_1971 ();
 sg13g2_decap_8 FILLER_27_2040 ();
 sg13g2_fill_2 FILLER_27_2047 ();
 sg13g2_fill_1 FILLER_27_2049 ();
 sg13g2_fill_2 FILLER_27_2075 ();
 sg13g2_fill_2 FILLER_27_2092 ();
 sg13g2_fill_1 FILLER_27_2104 ();
 sg13g2_fill_2 FILLER_27_2131 ();
 sg13g2_fill_1 FILLER_27_2138 ();
 sg13g2_fill_2 FILLER_27_2165 ();
 sg13g2_fill_1 FILLER_27_2203 ();
 sg13g2_fill_2 FILLER_27_2264 ();
 sg13g2_fill_1 FILLER_27_2266 ();
 sg13g2_fill_2 FILLER_27_2274 ();
 sg13g2_fill_1 FILLER_27_2276 ();
 sg13g2_fill_2 FILLER_27_2291 ();
 sg13g2_fill_1 FILLER_27_2293 ();
 sg13g2_decap_8 FILLER_27_2340 ();
 sg13g2_decap_8 FILLER_27_2347 ();
 sg13g2_fill_2 FILLER_27_2354 ();
 sg13g2_fill_1 FILLER_27_2364 ();
 sg13g2_fill_2 FILLER_27_2369 ();
 sg13g2_fill_2 FILLER_27_2375 ();
 sg13g2_fill_2 FILLER_27_2382 ();
 sg13g2_fill_1 FILLER_27_2388 ();
 sg13g2_fill_2 FILLER_27_2423 ();
 sg13g2_fill_1 FILLER_27_2425 ();
 sg13g2_fill_1 FILLER_27_2491 ();
 sg13g2_fill_1 FILLER_27_2557 ();
 sg13g2_fill_1 FILLER_27_2602 ();
 sg13g2_fill_1 FILLER_27_2626 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_5 ();
 sg13g2_fill_2 FILLER_28_17 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_decap_4 FILLER_28_285 ();
 sg13g2_fill_2 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_2 FILLER_28_424 ();
 sg13g2_fill_1 FILLER_28_426 ();
 sg13g2_fill_2 FILLER_28_457 ();
 sg13g2_fill_1 FILLER_28_489 ();
 sg13g2_fill_1 FILLER_28_495 ();
 sg13g2_decap_4 FILLER_28_508 ();
 sg13g2_fill_2 FILLER_28_521 ();
 sg13g2_decap_4 FILLER_28_527 ();
 sg13g2_fill_1 FILLER_28_531 ();
 sg13g2_fill_1 FILLER_28_536 ();
 sg13g2_decap_4 FILLER_28_585 ();
 sg13g2_fill_1 FILLER_28_589 ();
 sg13g2_decap_4 FILLER_28_595 ();
 sg13g2_fill_2 FILLER_28_599 ();
 sg13g2_fill_1 FILLER_28_605 ();
 sg13g2_fill_2 FILLER_28_623 ();
 sg13g2_fill_1 FILLER_28_637 ();
 sg13g2_fill_1 FILLER_28_644 ();
 sg13g2_decap_4 FILLER_28_660 ();
 sg13g2_fill_2 FILLER_28_701 ();
 sg13g2_fill_1 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_712 ();
 sg13g2_decap_4 FILLER_28_719 ();
 sg13g2_decap_4 FILLER_28_736 ();
 sg13g2_fill_2 FILLER_28_740 ();
 sg13g2_decap_4 FILLER_28_747 ();
 sg13g2_fill_1 FILLER_28_751 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_4 FILLER_28_763 ();
 sg13g2_fill_1 FILLER_28_767 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_4 FILLER_28_809 ();
 sg13g2_fill_1 FILLER_28_813 ();
 sg13g2_fill_1 FILLER_28_889 ();
 sg13g2_fill_1 FILLER_28_926 ();
 sg13g2_fill_1 FILLER_28_976 ();
 sg13g2_fill_2 FILLER_28_1003 ();
 sg13g2_fill_1 FILLER_28_1031 ();
 sg13g2_decap_4 FILLER_28_1120 ();
 sg13g2_fill_1 FILLER_28_1148 ();
 sg13g2_fill_2 FILLER_28_1182 ();
 sg13g2_fill_1 FILLER_28_1184 ();
 sg13g2_fill_1 FILLER_28_1190 ();
 sg13g2_fill_1 FILLER_28_1217 ();
 sg13g2_fill_2 FILLER_28_1222 ();
 sg13g2_fill_2 FILLER_28_1234 ();
 sg13g2_fill_1 FILLER_28_1262 ();
 sg13g2_decap_4 FILLER_28_1327 ();
 sg13g2_decap_8 FILLER_28_1334 ();
 sg13g2_fill_1 FILLER_28_1341 ();
 sg13g2_fill_2 FILLER_28_1346 ();
 sg13g2_fill_1 FILLER_28_1374 ();
 sg13g2_decap_4 FILLER_28_1413 ();
 sg13g2_fill_1 FILLER_28_1417 ();
 sg13g2_fill_2 FILLER_28_1434 ();
 sg13g2_fill_2 FILLER_28_1440 ();
 sg13g2_fill_1 FILLER_28_1445 ();
 sg13g2_fill_2 FILLER_28_1462 ();
 sg13g2_fill_1 FILLER_28_1476 ();
 sg13g2_fill_1 FILLER_28_1523 ();
 sg13g2_fill_2 FILLER_28_1537 ();
 sg13g2_decap_4 FILLER_28_1588 ();
 sg13g2_fill_2 FILLER_28_1592 ();
 sg13g2_decap_4 FILLER_28_1607 ();
 sg13g2_decap_4 FILLER_28_1620 ();
 sg13g2_fill_2 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_fill_2 FILLER_28_1638 ();
 sg13g2_decap_8 FILLER_28_1644 ();
 sg13g2_decap_8 FILLER_28_1651 ();
 sg13g2_decap_4 FILLER_28_1658 ();
 sg13g2_fill_1 FILLER_28_1662 ();
 sg13g2_decap_4 FILLER_28_1668 ();
 sg13g2_fill_1 FILLER_28_1672 ();
 sg13g2_decap_8 FILLER_28_1703 ();
 sg13g2_decap_8 FILLER_28_1710 ();
 sg13g2_decap_8 FILLER_28_1717 ();
 sg13g2_decap_8 FILLER_28_1724 ();
 sg13g2_decap_4 FILLER_28_1731 ();
 sg13g2_decap_8 FILLER_28_1743 ();
 sg13g2_decap_8 FILLER_28_1750 ();
 sg13g2_decap_4 FILLER_28_1761 ();
 sg13g2_fill_1 FILLER_28_1765 ();
 sg13g2_fill_2 FILLER_28_1792 ();
 sg13g2_fill_2 FILLER_28_1799 ();
 sg13g2_fill_1 FILLER_28_1801 ();
 sg13g2_decap_8 FILLER_28_1806 ();
 sg13g2_decap_4 FILLER_28_1813 ();
 sg13g2_fill_1 FILLER_28_1817 ();
 sg13g2_fill_2 FILLER_28_1823 ();
 sg13g2_fill_1 FILLER_28_1825 ();
 sg13g2_fill_2 FILLER_28_1833 ();
 sg13g2_fill_2 FILLER_28_1883 ();
 sg13g2_decap_8 FILLER_28_1905 ();
 sg13g2_fill_2 FILLER_28_1912 ();
 sg13g2_fill_1 FILLER_28_1928 ();
 sg13g2_fill_1 FILLER_28_1933 ();
 sg13g2_fill_2 FILLER_28_1960 ();
 sg13g2_fill_1 FILLER_28_1962 ();
 sg13g2_decap_8 FILLER_28_2021 ();
 sg13g2_decap_4 FILLER_28_2028 ();
 sg13g2_fill_2 FILLER_28_2032 ();
 sg13g2_decap_4 FILLER_28_2042 ();
 sg13g2_fill_2 FILLER_28_2103 ();
 sg13g2_fill_2 FILLER_28_2170 ();
 sg13g2_fill_2 FILLER_28_2182 ();
 sg13g2_fill_1 FILLER_28_2203 ();
 sg13g2_decap_8 FILLER_28_2261 ();
 sg13g2_decap_4 FILLER_28_2268 ();
 sg13g2_fill_2 FILLER_28_2272 ();
 sg13g2_fill_2 FILLER_28_2297 ();
 sg13g2_fill_1 FILLER_28_2299 ();
 sg13g2_fill_2 FILLER_28_2329 ();
 sg13g2_fill_1 FILLER_28_2331 ();
 sg13g2_decap_8 FILLER_28_2342 ();
 sg13g2_fill_1 FILLER_28_2349 ();
 sg13g2_fill_2 FILLER_28_2435 ();
 sg13g2_fill_2 FILLER_28_2443 ();
 sg13g2_fill_2 FILLER_28_2449 ();
 sg13g2_fill_1 FILLER_28_2456 ();
 sg13g2_decap_4 FILLER_28_2460 ();
 sg13g2_fill_2 FILLER_28_2464 ();
 sg13g2_fill_1 FILLER_28_2494 ();
 sg13g2_fill_2 FILLER_28_2500 ();
 sg13g2_fill_1 FILLER_28_2502 ();
 sg13g2_fill_2 FILLER_28_2511 ();
 sg13g2_fill_1 FILLER_28_2547 ();
 sg13g2_fill_1 FILLER_28_2587 ();
 sg13g2_fill_1 FILLER_28_2592 ();
 sg13g2_fill_2 FILLER_28_2616 ();
 sg13g2_decap_4 FILLER_28_2664 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_decap_4 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_1 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_422 ();
 sg13g2_fill_2 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_29_470 ();
 sg13g2_fill_1 FILLER_29_487 ();
 sg13g2_decap_4 FILLER_29_492 ();
 sg13g2_decap_8 FILLER_29_500 ();
 sg13g2_decap_8 FILLER_29_507 ();
 sg13g2_fill_2 FILLER_29_514 ();
 sg13g2_fill_1 FILLER_29_516 ();
 sg13g2_decap_8 FILLER_29_531 ();
 sg13g2_decap_8 FILLER_29_538 ();
 sg13g2_decap_8 FILLER_29_545 ();
 sg13g2_fill_2 FILLER_29_552 ();
 sg13g2_fill_1 FILLER_29_554 ();
 sg13g2_fill_1 FILLER_29_568 ();
 sg13g2_fill_1 FILLER_29_605 ();
 sg13g2_fill_1 FILLER_29_617 ();
 sg13g2_fill_1 FILLER_29_628 ();
 sg13g2_fill_2 FILLER_29_639 ();
 sg13g2_fill_2 FILLER_29_658 ();
 sg13g2_fill_1 FILLER_29_660 ();
 sg13g2_fill_2 FILLER_29_666 ();
 sg13g2_fill_2 FILLER_29_698 ();
 sg13g2_fill_2 FILLER_29_738 ();
 sg13g2_fill_1 FILLER_29_740 ();
 sg13g2_decap_8 FILLER_29_771 ();
 sg13g2_decap_4 FILLER_29_778 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_4 FILLER_29_807 ();
 sg13g2_fill_1 FILLER_29_815 ();
 sg13g2_fill_1 FILLER_29_886 ();
 sg13g2_fill_1 FILLER_29_900 ();
 sg13g2_fill_2 FILLER_29_927 ();
 sg13g2_fill_1 FILLER_29_934 ();
 sg13g2_fill_1 FILLER_29_974 ();
 sg13g2_fill_1 FILLER_29_979 ();
 sg13g2_fill_1 FILLER_29_987 ();
 sg13g2_fill_1 FILLER_29_998 ();
 sg13g2_fill_1 FILLER_29_1016 ();
 sg13g2_fill_2 FILLER_29_1051 ();
 sg13g2_fill_2 FILLER_29_1082 ();
 sg13g2_fill_2 FILLER_29_1091 ();
 sg13g2_fill_2 FILLER_29_1097 ();
 sg13g2_fill_1 FILLER_29_1135 ();
 sg13g2_fill_2 FILLER_29_1185 ();
 sg13g2_fill_2 FILLER_29_1269 ();
 sg13g2_decap_8 FILLER_29_1297 ();
 sg13g2_decap_8 FILLER_29_1304 ();
 sg13g2_fill_2 FILLER_29_1311 ();
 sg13g2_decap_8 FILLER_29_1316 ();
 sg13g2_fill_1 FILLER_29_1323 ();
 sg13g2_fill_1 FILLER_29_1344 ();
 sg13g2_decap_4 FILLER_29_1359 ();
 sg13g2_fill_2 FILLER_29_1379 ();
 sg13g2_fill_2 FILLER_29_1405 ();
 sg13g2_fill_2 FILLER_29_1445 ();
 sg13g2_fill_2 FILLER_29_1495 ();
 sg13g2_fill_1 FILLER_29_1509 ();
 sg13g2_fill_2 FILLER_29_1534 ();
 sg13g2_fill_2 FILLER_29_1541 ();
 sg13g2_fill_1 FILLER_29_1576 ();
 sg13g2_fill_2 FILLER_29_1595 ();
 sg13g2_decap_8 FILLER_29_1612 ();
 sg13g2_decap_8 FILLER_29_1619 ();
 sg13g2_decap_8 FILLER_29_1626 ();
 sg13g2_decap_8 FILLER_29_1633 ();
 sg13g2_decap_8 FILLER_29_1640 ();
 sg13g2_decap_8 FILLER_29_1647 ();
 sg13g2_decap_4 FILLER_29_1654 ();
 sg13g2_decap_4 FILLER_29_1663 ();
 sg13g2_fill_2 FILLER_29_1667 ();
 sg13g2_decap_8 FILLER_29_1695 ();
 sg13g2_decap_8 FILLER_29_1702 ();
 sg13g2_fill_2 FILLER_29_1709 ();
 sg13g2_fill_1 FILLER_29_1711 ();
 sg13g2_decap_4 FILLER_29_1717 ();
 sg13g2_fill_1 FILLER_29_1721 ();
 sg13g2_decap_8 FILLER_29_1726 ();
 sg13g2_decap_8 FILLER_29_1733 ();
 sg13g2_decap_8 FILLER_29_1740 ();
 sg13g2_decap_8 FILLER_29_1747 ();
 sg13g2_decap_4 FILLER_29_1758 ();
 sg13g2_decap_8 FILLER_29_1823 ();
 sg13g2_fill_2 FILLER_29_1859 ();
 sg13g2_decap_4 FILLER_29_1955 ();
 sg13g2_fill_2 FILLER_29_1959 ();
 sg13g2_fill_2 FILLER_29_1971 ();
 sg13g2_fill_2 FILLER_29_1994 ();
 sg13g2_decap_8 FILLER_29_2000 ();
 sg13g2_fill_1 FILLER_29_2007 ();
 sg13g2_decap_4 FILLER_29_2016 ();
 sg13g2_decap_4 FILLER_29_2024 ();
 sg13g2_decap_4 FILLER_29_2036 ();
 sg13g2_fill_1 FILLER_29_2040 ();
 sg13g2_fill_1 FILLER_29_2045 ();
 sg13g2_decap_4 FILLER_29_2156 ();
 sg13g2_fill_2 FILLER_29_2160 ();
 sg13g2_decap_8 FILLER_29_2260 ();
 sg13g2_fill_2 FILLER_29_2267 ();
 sg13g2_fill_1 FILLER_29_2269 ();
 sg13g2_fill_2 FILLER_29_2358 ();
 sg13g2_fill_1 FILLER_29_2417 ();
 sg13g2_fill_1 FILLER_29_2442 ();
 sg13g2_decap_4 FILLER_29_2453 ();
 sg13g2_decap_4 FILLER_29_2466 ();
 sg13g2_decap_4 FILLER_29_2474 ();
 sg13g2_fill_2 FILLER_29_2495 ();
 sg13g2_fill_1 FILLER_29_2497 ();
 sg13g2_fill_1 FILLER_29_2511 ();
 sg13g2_fill_1 FILLER_29_2520 ();
 sg13g2_fill_1 FILLER_29_2530 ();
 sg13g2_fill_1 FILLER_29_2544 ();
 sg13g2_fill_2 FILLER_29_2591 ();
 sg13g2_fill_1 FILLER_29_2635 ();
 sg13g2_fill_2 FILLER_29_2640 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_61 ();
 sg13g2_fill_2 FILLER_30_66 ();
 sg13g2_fill_1 FILLER_30_68 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_decap_4 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_159 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_384 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_431 ();
 sg13g2_fill_2 FILLER_30_498 ();
 sg13g2_decap_8 FILLER_30_530 ();
 sg13g2_decap_8 FILLER_30_537 ();
 sg13g2_decap_8 FILLER_30_544 ();
 sg13g2_decap_4 FILLER_30_551 ();
 sg13g2_fill_1 FILLER_30_555 ();
 sg13g2_fill_1 FILLER_30_569 ();
 sg13g2_fill_1 FILLER_30_580 ();
 sg13g2_fill_1 FILLER_30_586 ();
 sg13g2_fill_2 FILLER_30_613 ();
 sg13g2_fill_1 FILLER_30_632 ();
 sg13g2_fill_1 FILLER_30_659 ();
 sg13g2_fill_1 FILLER_30_692 ();
 sg13g2_decap_4 FILLER_30_753 ();
 sg13g2_fill_1 FILLER_30_766 ();
 sg13g2_decap_4 FILLER_30_772 ();
 sg13g2_fill_1 FILLER_30_776 ();
 sg13g2_decap_8 FILLER_30_783 ();
 sg13g2_fill_1 FILLER_30_790 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_fill_2 FILLER_30_835 ();
 sg13g2_fill_1 FILLER_30_867 ();
 sg13g2_fill_2 FILLER_30_894 ();
 sg13g2_fill_1 FILLER_30_938 ();
 sg13g2_fill_1 FILLER_30_987 ();
 sg13g2_fill_1 FILLER_30_1010 ();
 sg13g2_fill_1 FILLER_30_1021 ();
 sg13g2_fill_1 FILLER_30_1055 ();
 sg13g2_fill_2 FILLER_30_1083 ();
 sg13g2_fill_2 FILLER_30_1120 ();
 sg13g2_fill_1 FILLER_30_1125 ();
 sg13g2_fill_2 FILLER_30_1189 ();
 sg13g2_fill_1 FILLER_30_1191 ();
 sg13g2_fill_2 FILLER_30_1260 ();
 sg13g2_fill_1 FILLER_30_1305 ();
 sg13g2_decap_4 FILLER_30_1326 ();
 sg13g2_fill_1 FILLER_30_1330 ();
 sg13g2_decap_4 FILLER_30_1334 ();
 sg13g2_fill_1 FILLER_30_1470 ();
 sg13g2_fill_1 FILLER_30_1486 ();
 sg13g2_fill_1 FILLER_30_1496 ();
 sg13g2_fill_1 FILLER_30_1516 ();
 sg13g2_fill_1 FILLER_30_1521 ();
 sg13g2_decap_4 FILLER_30_1566 ();
 sg13g2_fill_1 FILLER_30_1570 ();
 sg13g2_fill_2 FILLER_30_1579 ();
 sg13g2_fill_1 FILLER_30_1581 ();
 sg13g2_decap_4 FILLER_30_1599 ();
 sg13g2_fill_1 FILLER_30_1603 ();
 sg13g2_decap_8 FILLER_30_1608 ();
 sg13g2_decap_8 FILLER_30_1615 ();
 sg13g2_decap_8 FILLER_30_1622 ();
 sg13g2_decap_4 FILLER_30_1629 ();
 sg13g2_fill_1 FILLER_30_1633 ();
 sg13g2_decap_4 FILLER_30_1654 ();
 sg13g2_fill_1 FILLER_30_1658 ();
 sg13g2_decap_4 FILLER_30_1672 ();
 sg13g2_fill_2 FILLER_30_1676 ();
 sg13g2_decap_4 FILLER_30_1682 ();
 sg13g2_decap_8 FILLER_30_1720 ();
 sg13g2_decap_8 FILLER_30_1727 ();
 sg13g2_fill_2 FILLER_30_1734 ();
 sg13g2_fill_2 FILLER_30_1745 ();
 sg13g2_fill_1 FILLER_30_1747 ();
 sg13g2_fill_1 FILLER_30_1870 ();
 sg13g2_fill_2 FILLER_30_1897 ();
 sg13g2_fill_1 FILLER_30_1946 ();
 sg13g2_fill_2 FILLER_30_1951 ();
 sg13g2_fill_2 FILLER_30_1963 ();
 sg13g2_decap_8 FILLER_30_1985 ();
 sg13g2_decap_4 FILLER_30_1992 ();
 sg13g2_fill_2 FILLER_30_2040 ();
 sg13g2_fill_1 FILLER_30_2042 ();
 sg13g2_decap_4 FILLER_30_2069 ();
 sg13g2_fill_2 FILLER_30_2073 ();
 sg13g2_fill_2 FILLER_30_2101 ();
 sg13g2_fill_1 FILLER_30_2108 ();
 sg13g2_fill_2 FILLER_30_2124 ();
 sg13g2_fill_1 FILLER_30_2126 ();
 sg13g2_fill_2 FILLER_30_2188 ();
 sg13g2_decap_4 FILLER_30_2278 ();
 sg13g2_fill_2 FILLER_30_2312 ();
 sg13g2_fill_1 FILLER_30_2314 ();
 sg13g2_decap_4 FILLER_30_2319 ();
 sg13g2_fill_2 FILLER_30_2323 ();
 sg13g2_fill_2 FILLER_30_2359 ();
 sg13g2_fill_2 FILLER_30_2375 ();
 sg13g2_fill_1 FILLER_30_2421 ();
 sg13g2_decap_4 FILLER_30_2452 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_87 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_174 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_258 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_2 FILLER_31_288 ();
 sg13g2_fill_1 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_decap_4 FILLER_31_350 ();
 sg13g2_fill_2 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_decap_4 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_31_416 ();
 sg13g2_fill_2 FILLER_31_422 ();
 sg13g2_decap_8 FILLER_31_491 ();
 sg13g2_decap_8 FILLER_31_498 ();
 sg13g2_fill_1 FILLER_31_505 ();
 sg13g2_fill_2 FILLER_31_532 ();
 sg13g2_fill_1 FILLER_31_578 ();
 sg13g2_fill_1 FILLER_31_601 ();
 sg13g2_fill_2 FILLER_31_630 ();
 sg13g2_fill_1 FILLER_31_685 ();
 sg13g2_fill_1 FILLER_31_695 ();
 sg13g2_fill_2 FILLER_31_714 ();
 sg13g2_fill_1 FILLER_31_720 ();
 sg13g2_fill_2 FILLER_31_727 ();
 sg13g2_fill_2 FILLER_31_734 ();
 sg13g2_fill_1 FILLER_31_736 ();
 sg13g2_fill_2 FILLER_31_741 ();
 sg13g2_fill_1 FILLER_31_743 ();
 sg13g2_fill_2 FILLER_31_788 ();
 sg13g2_fill_1 FILLER_31_795 ();
 sg13g2_fill_2 FILLER_31_822 ();
 sg13g2_fill_1 FILLER_31_834 ();
 sg13g2_fill_2 FILLER_31_925 ();
 sg13g2_fill_1 FILLER_31_950 ();
 sg13g2_fill_2 FILLER_31_977 ();
 sg13g2_fill_2 FILLER_31_983 ();
 sg13g2_fill_2 FILLER_31_989 ();
 sg13g2_fill_1 FILLER_31_1043 ();
 sg13g2_fill_1 FILLER_31_1091 ();
 sg13g2_fill_2 FILLER_31_1109 ();
 sg13g2_fill_1 FILLER_31_1121 ();
 sg13g2_decap_8 FILLER_31_1168 ();
 sg13g2_fill_1 FILLER_31_1175 ();
 sg13g2_decap_8 FILLER_31_1181 ();
 sg13g2_decap_8 FILLER_31_1188 ();
 sg13g2_fill_1 FILLER_31_1195 ();
 sg13g2_fill_1 FILLER_31_1218 ();
 sg13g2_fill_2 FILLER_31_1276 ();
 sg13g2_fill_1 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1306 ();
 sg13g2_decap_8 FILLER_31_1316 ();
 sg13g2_decap_8 FILLER_31_1323 ();
 sg13g2_fill_2 FILLER_31_1330 ();
 sg13g2_fill_1 FILLER_31_1332 ();
 sg13g2_decap_8 FILLER_31_1359 ();
 sg13g2_decap_8 FILLER_31_1366 ();
 sg13g2_decap_4 FILLER_31_1373 ();
 sg13g2_fill_2 FILLER_31_1381 ();
 sg13g2_fill_2 FILLER_31_1436 ();
 sg13g2_fill_2 FILLER_31_1454 ();
 sg13g2_fill_1 FILLER_31_1491 ();
 sg13g2_fill_1 FILLER_31_1519 ();
 sg13g2_fill_1 FILLER_31_1524 ();
 sg13g2_decap_8 FILLER_31_1573 ();
 sg13g2_fill_1 FILLER_31_1580 ();
 sg13g2_fill_1 FILLER_31_1586 ();
 sg13g2_decap_8 FILLER_31_1591 ();
 sg13g2_decap_4 FILLER_31_1598 ();
 sg13g2_decap_4 FILLER_31_1615 ();
 sg13g2_fill_1 FILLER_31_1619 ();
 sg13g2_fill_2 FILLER_31_1643 ();
 sg13g2_fill_1 FILLER_31_1645 ();
 sg13g2_decap_8 FILLER_31_1782 ();
 sg13g2_fill_2 FILLER_31_1789 ();
 sg13g2_fill_1 FILLER_31_1791 ();
 sg13g2_decap_4 FILLER_31_1832 ();
 sg13g2_fill_1 FILLER_31_1836 ();
 sg13g2_fill_2 FILLER_31_1887 ();
 sg13g2_fill_1 FILLER_31_1889 ();
 sg13g2_decap_4 FILLER_31_1900 ();
 sg13g2_fill_2 FILLER_31_1933 ();
 sg13g2_fill_2 FILLER_31_1938 ();
 sg13g2_fill_1 FILLER_31_1954 ();
 sg13g2_fill_1 FILLER_31_1981 ();
 sg13g2_fill_1 FILLER_31_1992 ();
 sg13g2_fill_1 FILLER_31_2019 ();
 sg13g2_fill_2 FILLER_31_2051 ();
 sg13g2_fill_1 FILLER_31_2084 ();
 sg13g2_fill_1 FILLER_31_2089 ();
 sg13g2_fill_2 FILLER_31_2106 ();
 sg13g2_fill_1 FILLER_31_2108 ();
 sg13g2_fill_1 FILLER_31_2139 ();
 sg13g2_decap_8 FILLER_31_2150 ();
 sg13g2_fill_1 FILLER_31_2157 ();
 sg13g2_decap_4 FILLER_31_2179 ();
 sg13g2_fill_2 FILLER_31_2220 ();
 sg13g2_decap_8 FILLER_31_2278 ();
 sg13g2_fill_1 FILLER_31_2285 ();
 sg13g2_decap_4 FILLER_31_2296 ();
 sg13g2_fill_1 FILLER_31_2300 ();
 sg13g2_decap_8 FILLER_31_2353 ();
 sg13g2_fill_2 FILLER_31_2360 ();
 sg13g2_decap_8 FILLER_31_2372 ();
 sg13g2_decap_8 FILLER_31_2379 ();
 sg13g2_decap_4 FILLER_31_2386 ();
 sg13g2_fill_2 FILLER_31_2390 ();
 sg13g2_fill_1 FILLER_31_2422 ();
 sg13g2_decap_8 FILLER_31_2449 ();
 sg13g2_decap_4 FILLER_31_2459 ();
 sg13g2_fill_2 FILLER_31_2463 ();
 sg13g2_decap_4 FILLER_31_2469 ();
 sg13g2_fill_2 FILLER_31_2481 ();
 sg13g2_fill_2 FILLER_31_2493 ();
 sg13g2_fill_1 FILLER_31_2495 ();
 sg13g2_decap_8 FILLER_31_2500 ();
 sg13g2_decap_4 FILLER_31_2507 ();
 sg13g2_fill_2 FILLER_31_2511 ();
 sg13g2_fill_2 FILLER_31_2519 ();
 sg13g2_fill_1 FILLER_31_2556 ();
 sg13g2_fill_1 FILLER_31_2565 ();
 sg13g2_fill_1 FILLER_31_2571 ();
 sg13g2_fill_1 FILLER_31_2607 ();
 sg13g2_fill_1 FILLER_31_2640 ();
 sg13g2_fill_1 FILLER_31_2645 ();
 sg13g2_fill_2 FILLER_31_2660 ();
 sg13g2_decap_4 FILLER_31_2666 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_fill_1 FILLER_32_82 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_fill_2 FILLER_32_417 ();
 sg13g2_fill_1 FILLER_32_419 ();
 sg13g2_fill_2 FILLER_32_436 ();
 sg13g2_fill_2 FILLER_32_443 ();
 sg13g2_fill_1 FILLER_32_445 ();
 sg13g2_fill_2 FILLER_32_472 ();
 sg13g2_fill_1 FILLER_32_479 ();
 sg13g2_fill_1 FILLER_32_492 ();
 sg13g2_fill_1 FILLER_32_498 ();
 sg13g2_fill_1 FILLER_32_519 ();
 sg13g2_fill_1 FILLER_32_530 ();
 sg13g2_fill_1 FILLER_32_541 ();
 sg13g2_decap_4 FILLER_32_546 ();
 sg13g2_fill_2 FILLER_32_550 ();
 sg13g2_fill_1 FILLER_32_582 ();
 sg13g2_fill_2 FILLER_32_592 ();
 sg13g2_fill_2 FILLER_32_619 ();
 sg13g2_fill_1 FILLER_32_640 ();
 sg13g2_fill_1 FILLER_32_645 ();
 sg13g2_fill_1 FILLER_32_672 ();
 sg13g2_fill_1 FILLER_32_682 ();
 sg13g2_fill_2 FILLER_32_691 ();
 sg13g2_fill_1 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_710 ();
 sg13g2_fill_1 FILLER_32_717 ();
 sg13g2_decap_4 FILLER_32_741 ();
 sg13g2_fill_1 FILLER_32_745 ();
 sg13g2_fill_2 FILLER_32_834 ();
 sg13g2_fill_1 FILLER_32_856 ();
 sg13g2_fill_2 FILLER_32_862 ();
 sg13g2_fill_1 FILLER_32_895 ();
 sg13g2_fill_2 FILLER_32_912 ();
 sg13g2_fill_2 FILLER_32_925 ();
 sg13g2_fill_1 FILLER_32_951 ();
 sg13g2_fill_1 FILLER_32_959 ();
 sg13g2_fill_2 FILLER_32_970 ();
 sg13g2_fill_2 FILLER_32_1052 ();
 sg13g2_fill_1 FILLER_32_1084 ();
 sg13g2_fill_2 FILLER_32_1092 ();
 sg13g2_decap_4 FILLER_32_1107 ();
 sg13g2_decap_8 FILLER_32_1114 ();
 sg13g2_fill_1 FILLER_32_1121 ();
 sg13g2_fill_1 FILLER_32_1125 ();
 sg13g2_fill_1 FILLER_32_1152 ();
 sg13g2_decap_8 FILLER_32_1159 ();
 sg13g2_fill_2 FILLER_32_1166 ();
 sg13g2_fill_1 FILLER_32_1168 ();
 sg13g2_decap_4 FILLER_32_1203 ();
 sg13g2_fill_1 FILLER_32_1233 ();
 sg13g2_fill_1 FILLER_32_1280 ();
 sg13g2_fill_1 FILLER_32_1291 ();
 sg13g2_fill_1 FILLER_32_1296 ();
 sg13g2_fill_2 FILLER_32_1333 ();
 sg13g2_fill_1 FILLER_32_1335 ();
 sg13g2_fill_2 FILLER_32_1343 ();
 sg13g2_fill_2 FILLER_32_1375 ();
 sg13g2_fill_2 FILLER_32_1381 ();
 sg13g2_fill_2 FILLER_32_1398 ();
 sg13g2_fill_1 FILLER_32_1452 ();
 sg13g2_fill_1 FILLER_32_1478 ();
 sg13g2_fill_1 FILLER_32_1489 ();
 sg13g2_fill_2 FILLER_32_1548 ();
 sg13g2_fill_2 FILLER_32_1612 ();
 sg13g2_fill_1 FILLER_32_1614 ();
 sg13g2_fill_2 FILLER_32_1619 ();
 sg13g2_fill_1 FILLER_32_1621 ();
 sg13g2_fill_2 FILLER_32_1653 ();
 sg13g2_fill_1 FILLER_32_1655 ();
 sg13g2_decap_4 FILLER_32_1662 ();
 sg13g2_fill_1 FILLER_32_1670 ();
 sg13g2_fill_2 FILLER_32_1680 ();
 sg13g2_fill_2 FILLER_32_1688 ();
 sg13g2_fill_2 FILLER_32_1714 ();
 sg13g2_fill_2 FILLER_32_1741 ();
 sg13g2_decap_4 FILLER_32_1778 ();
 sg13g2_fill_1 FILLER_32_1782 ();
 sg13g2_decap_4 FILLER_32_1791 ();
 sg13g2_fill_2 FILLER_32_1795 ();
 sg13g2_decap_8 FILLER_32_1827 ();
 sg13g2_decap_8 FILLER_32_1834 ();
 sg13g2_decap_8 FILLER_32_1841 ();
 sg13g2_fill_1 FILLER_32_1848 ();
 sg13g2_decap_4 FILLER_32_1875 ();
 sg13g2_fill_1 FILLER_32_1879 ();
 sg13g2_decap_8 FILLER_32_1893 ();
 sg13g2_decap_4 FILLER_32_1900 ();
 sg13g2_fill_2 FILLER_32_1904 ();
 sg13g2_fill_2 FILLER_32_1910 ();
 sg13g2_fill_2 FILLER_32_1916 ();
 sg13g2_fill_2 FILLER_32_2004 ();
 sg13g2_fill_1 FILLER_32_2010 ();
 sg13g2_fill_2 FILLER_32_2021 ();
 sg13g2_fill_2 FILLER_32_2049 ();
 sg13g2_fill_2 FILLER_32_2055 ();
 sg13g2_fill_1 FILLER_32_2083 ();
 sg13g2_fill_2 FILLER_32_2088 ();
 sg13g2_fill_1 FILLER_32_2090 ();
 sg13g2_fill_2 FILLER_32_2095 ();
 sg13g2_fill_1 FILLER_32_2097 ();
 sg13g2_fill_1 FILLER_32_2138 ();
 sg13g2_fill_2 FILLER_32_2169 ();
 sg13g2_fill_1 FILLER_32_2171 ();
 sg13g2_fill_1 FILLER_32_2219 ();
 sg13g2_fill_1 FILLER_32_2230 ();
 sg13g2_decap_4 FILLER_32_2241 ();
 sg13g2_fill_2 FILLER_32_2245 ();
 sg13g2_fill_2 FILLER_32_2272 ();
 sg13g2_fill_1 FILLER_32_2274 ();
 sg13g2_decap_4 FILLER_32_2357 ();
 sg13g2_fill_1 FILLER_32_2361 ();
 sg13g2_fill_2 FILLER_32_2407 ();
 sg13g2_fill_1 FILLER_32_2409 ();
 sg13g2_fill_2 FILLER_32_2441 ();
 sg13g2_fill_1 FILLER_32_2443 ();
 sg13g2_fill_2 FILLER_32_2456 ();
 sg13g2_fill_1 FILLER_32_2458 ();
 sg13g2_decap_4 FILLER_32_2497 ();
 sg13g2_fill_2 FILLER_32_2501 ();
 sg13g2_fill_2 FILLER_32_2514 ();
 sg13g2_fill_1 FILLER_32_2533 ();
 sg13g2_fill_2 FILLER_32_2668 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_decap_4 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_decap_4 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_244 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_decap_4 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_315 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_4 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_368 ();
 sg13g2_fill_2 FILLER_33_414 ();
 sg13g2_decap_4 FILLER_33_420 ();
 sg13g2_fill_1 FILLER_33_424 ();
 sg13g2_decap_4 FILLER_33_434 ();
 sg13g2_fill_1 FILLER_33_438 ();
 sg13g2_fill_1 FILLER_33_443 ();
 sg13g2_fill_2 FILLER_33_498 ();
 sg13g2_fill_1 FILLER_33_500 ();
 sg13g2_fill_2 FILLER_33_535 ();
 sg13g2_fill_1 FILLER_33_537 ();
 sg13g2_fill_1 FILLER_33_558 ();
 sg13g2_fill_1 FILLER_33_585 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_fill_2 FILLER_33_625 ();
 sg13g2_fill_2 FILLER_33_659 ();
 sg13g2_fill_2 FILLER_33_671 ();
 sg13g2_decap_4 FILLER_33_709 ();
 sg13g2_fill_1 FILLER_33_713 ();
 sg13g2_fill_2 FILLER_33_723 ();
 sg13g2_fill_1 FILLER_33_725 ();
 sg13g2_fill_1 FILLER_33_737 ();
 sg13g2_fill_1 FILLER_33_748 ();
 sg13g2_fill_1 FILLER_33_806 ();
 sg13g2_fill_1 FILLER_33_860 ();
 sg13g2_fill_1 FILLER_33_961 ();
 sg13g2_fill_1 FILLER_33_988 ();
 sg13g2_fill_2 FILLER_33_1032 ();
 sg13g2_fill_2 FILLER_33_1038 ();
 sg13g2_fill_2 FILLER_33_1043 ();
 sg13g2_fill_1 FILLER_33_1049 ();
 sg13g2_fill_1 FILLER_33_1057 ();
 sg13g2_fill_2 FILLER_33_1115 ();
 sg13g2_fill_1 FILLER_33_1117 ();
 sg13g2_decap_8 FILLER_33_1148 ();
 sg13g2_fill_1 FILLER_33_1155 ();
 sg13g2_decap_8 FILLER_33_1186 ();
 sg13g2_fill_1 FILLER_33_1193 ();
 sg13g2_fill_1 FILLER_33_1215 ();
 sg13g2_fill_2 FILLER_33_1242 ();
 sg13g2_fill_2 FILLER_33_1256 ();
 sg13g2_fill_2 FILLER_33_1270 ();
 sg13g2_fill_2 FILLER_33_1334 ();
 sg13g2_decap_8 FILLER_33_1346 ();
 sg13g2_fill_1 FILLER_33_1353 ();
 sg13g2_fill_2 FILLER_33_1427 ();
 sg13g2_fill_2 FILLER_33_1433 ();
 sg13g2_fill_2 FILLER_33_1448 ();
 sg13g2_fill_1 FILLER_33_1494 ();
 sg13g2_fill_2 FILLER_33_1524 ();
 sg13g2_fill_1 FILLER_33_1526 ();
 sg13g2_fill_1 FILLER_33_1540 ();
 sg13g2_decap_8 FILLER_33_1550 ();
 sg13g2_decap_8 FILLER_33_1557 ();
 sg13g2_fill_2 FILLER_33_1564 ();
 sg13g2_fill_2 FILLER_33_1571 ();
 sg13g2_decap_8 FILLER_33_1581 ();
 sg13g2_fill_2 FILLER_33_1588 ();
 sg13g2_fill_1 FILLER_33_1590 ();
 sg13g2_decap_8 FILLER_33_1596 ();
 sg13g2_fill_1 FILLER_33_1607 ();
 sg13g2_fill_1 FILLER_33_1687 ();
 sg13g2_fill_1 FILLER_33_1744 ();
 sg13g2_fill_2 FILLER_33_1785 ();
 sg13g2_decap_8 FILLER_33_1791 ();
 sg13g2_decap_4 FILLER_33_1798 ();
 sg13g2_decap_8 FILLER_33_1812 ();
 sg13g2_fill_2 FILLER_33_1852 ();
 sg13g2_fill_2 FILLER_33_1873 ();
 sg13g2_fill_2 FILLER_33_1883 ();
 sg13g2_decap_8 FILLER_33_1889 ();
 sg13g2_fill_2 FILLER_33_1896 ();
 sg13g2_fill_1 FILLER_33_1898 ();
 sg13g2_fill_1 FILLER_33_1994 ();
 sg13g2_fill_2 FILLER_33_2005 ();
 sg13g2_fill_2 FILLER_33_2046 ();
 sg13g2_fill_1 FILLER_33_2048 ();
 sg13g2_decap_8 FILLER_33_2062 ();
 sg13g2_decap_8 FILLER_33_2069 ();
 sg13g2_decap_8 FILLER_33_2076 ();
 sg13g2_fill_1 FILLER_33_2083 ();
 sg13g2_decap_8 FILLER_33_2089 ();
 sg13g2_decap_4 FILLER_33_2096 ();
 sg13g2_fill_2 FILLER_33_2100 ();
 sg13g2_fill_2 FILLER_33_2114 ();
 sg13g2_fill_1 FILLER_33_2120 ();
 sg13g2_fill_2 FILLER_33_2147 ();
 sg13g2_fill_2 FILLER_33_2170 ();
 sg13g2_fill_2 FILLER_33_2182 ();
 sg13g2_decap_8 FILLER_33_2236 ();
 sg13g2_decap_8 FILLER_33_2243 ();
 sg13g2_decap_8 FILLER_33_2250 ();
 sg13g2_fill_2 FILLER_33_2257 ();
 sg13g2_fill_1 FILLER_33_2259 ();
 sg13g2_fill_2 FILLER_33_2281 ();
 sg13g2_fill_2 FILLER_33_2309 ();
 sg13g2_fill_1 FILLER_33_2311 ();
 sg13g2_decap_4 FILLER_33_2316 ();
 sg13g2_fill_2 FILLER_33_2320 ();
 sg13g2_fill_2 FILLER_33_2335 ();
 sg13g2_fill_1 FILLER_33_2337 ();
 sg13g2_decap_8 FILLER_33_2342 ();
 sg13g2_decap_4 FILLER_33_2349 ();
 sg13g2_fill_1 FILLER_33_2353 ();
 sg13g2_fill_2 FILLER_33_2372 ();
 sg13g2_decap_4 FILLER_33_2400 ();
 sg13g2_fill_2 FILLER_33_2409 ();
 sg13g2_fill_2 FILLER_33_2419 ();
 sg13g2_fill_1 FILLER_33_2421 ();
 sg13g2_fill_2 FILLER_33_2461 ();
 sg13g2_fill_2 FILLER_33_2468 ();
 sg13g2_decap_4 FILLER_33_2479 ();
 sg13g2_fill_1 FILLER_33_2497 ();
 sg13g2_fill_1 FILLER_33_2534 ();
 sg13g2_fill_1 FILLER_33_2551 ();
 sg13g2_fill_2 FILLER_33_2579 ();
 sg13g2_fill_2 FILLER_33_2599 ();
 sg13g2_decap_8 FILLER_33_2663 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_36 ();
 sg13g2_decap_8 FILLER_34_41 ();
 sg13g2_decap_8 FILLER_34_48 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_62 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_80 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_132 ();
 sg13g2_decap_4 FILLER_34_139 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_decap_4 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_decap_4 FILLER_34_449 ();
 sg13g2_fill_1 FILLER_34_453 ();
 sg13g2_fill_1 FILLER_34_458 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_fill_2 FILLER_34_475 ();
 sg13g2_fill_1 FILLER_34_477 ();
 sg13g2_decap_8 FILLER_34_491 ();
 sg13g2_fill_2 FILLER_34_518 ();
 sg13g2_fill_1 FILLER_34_524 ();
 sg13g2_fill_2 FILLER_34_543 ();
 sg13g2_fill_1 FILLER_34_545 ();
 sg13g2_fill_2 FILLER_34_664 ();
 sg13g2_fill_2 FILLER_34_671 ();
 sg13g2_fill_1 FILLER_34_678 ();
 sg13g2_fill_1 FILLER_34_689 ();
 sg13g2_fill_2 FILLER_34_694 ();
 sg13g2_decap_8 FILLER_34_703 ();
 sg13g2_decap_8 FILLER_34_710 ();
 sg13g2_decap_4 FILLER_34_717 ();
 sg13g2_fill_1 FILLER_34_721 ();
 sg13g2_decap_4 FILLER_34_736 ();
 sg13g2_fill_2 FILLER_34_758 ();
 sg13g2_fill_2 FILLER_34_796 ();
 sg13g2_fill_2 FILLER_34_819 ();
 sg13g2_fill_2 FILLER_34_877 ();
 sg13g2_fill_2 FILLER_34_923 ();
 sg13g2_fill_2 FILLER_34_948 ();
 sg13g2_fill_2 FILLER_34_969 ();
 sg13g2_fill_1 FILLER_34_1019 ();
 sg13g2_fill_2 FILLER_34_1024 ();
 sg13g2_fill_1 FILLER_34_1033 ();
 sg13g2_fill_1 FILLER_34_1039 ();
 sg13g2_fill_2 FILLER_34_1071 ();
 sg13g2_fill_1 FILLER_34_1080 ();
 sg13g2_fill_2 FILLER_34_1098 ();
 sg13g2_fill_1 FILLER_34_1100 ();
 sg13g2_decap_8 FILLER_34_1131 ();
 sg13g2_decap_8 FILLER_34_1138 ();
 sg13g2_decap_8 FILLER_34_1145 ();
 sg13g2_decap_8 FILLER_34_1152 ();
 sg13g2_decap_8 FILLER_34_1159 ();
 sg13g2_fill_2 FILLER_34_1166 ();
 sg13g2_fill_2 FILLER_34_1172 ();
 sg13g2_fill_1 FILLER_34_1174 ();
 sg13g2_decap_8 FILLER_34_1184 ();
 sg13g2_fill_2 FILLER_34_1191 ();
 sg13g2_fill_1 FILLER_34_1325 ();
 sg13g2_decap_8 FILLER_34_1339 ();
 sg13g2_decap_8 FILLER_34_1346 ();
 sg13g2_decap_4 FILLER_34_1353 ();
 sg13g2_fill_2 FILLER_34_1416 ();
 sg13g2_fill_1 FILLER_34_1434 ();
 sg13g2_fill_2 FILLER_34_1445 ();
 sg13g2_fill_1 FILLER_34_1468 ();
 sg13g2_decap_8 FILLER_34_1508 ();
 sg13g2_fill_2 FILLER_34_1515 ();
 sg13g2_fill_1 FILLER_34_1517 ();
 sg13g2_decap_8 FILLER_34_1546 ();
 sg13g2_fill_2 FILLER_34_1553 ();
 sg13g2_fill_1 FILLER_34_1555 ();
 sg13g2_fill_2 FILLER_34_1581 ();
 sg13g2_fill_1 FILLER_34_1583 ();
 sg13g2_decap_8 FILLER_34_1589 ();
 sg13g2_fill_1 FILLER_34_1596 ();
 sg13g2_decap_8 FILLER_34_1607 ();
 sg13g2_decap_4 FILLER_34_1614 ();
 sg13g2_fill_1 FILLER_34_1618 ();
 sg13g2_fill_2 FILLER_34_1624 ();
 sg13g2_fill_2 FILLER_34_1630 ();
 sg13g2_fill_1 FILLER_34_1632 ();
 sg13g2_fill_2 FILLER_34_1638 ();
 sg13g2_fill_1 FILLER_34_1640 ();
 sg13g2_fill_2 FILLER_34_1645 ();
 sg13g2_fill_2 FILLER_34_1651 ();
 sg13g2_fill_2 FILLER_34_1674 ();
 sg13g2_fill_1 FILLER_34_1726 ();
 sg13g2_fill_1 FILLER_34_1736 ();
 sg13g2_fill_1 FILLER_34_1808 ();
 sg13g2_decap_8 FILLER_34_1814 ();
 sg13g2_decap_4 FILLER_34_1821 ();
 sg13g2_decap_4 FILLER_34_1829 ();
 sg13g2_fill_1 FILLER_34_1846 ();
 sg13g2_fill_1 FILLER_34_1856 ();
 sg13g2_fill_2 FILLER_34_1867 ();
 sg13g2_fill_2 FILLER_34_1954 ();
 sg13g2_fill_1 FILLER_34_1997 ();
 sg13g2_fill_2 FILLER_34_2095 ();
 sg13g2_fill_1 FILLER_34_2097 ();
 sg13g2_fill_1 FILLER_34_2103 ();
 sg13g2_decap_4 FILLER_34_2109 ();
 sg13g2_fill_1 FILLER_34_2113 ();
 sg13g2_fill_1 FILLER_34_2128 ();
 sg13g2_decap_8 FILLER_34_2133 ();
 sg13g2_decap_8 FILLER_34_2140 ();
 sg13g2_fill_1 FILLER_34_2194 ();
 sg13g2_fill_2 FILLER_34_2199 ();
 sg13g2_fill_1 FILLER_34_2201 ();
 sg13g2_fill_2 FILLER_34_2215 ();
 sg13g2_decap_8 FILLER_34_2221 ();
 sg13g2_decap_4 FILLER_34_2228 ();
 sg13g2_fill_1 FILLER_34_2232 ();
 sg13g2_fill_1 FILLER_34_2254 ();
 sg13g2_fill_2 FILLER_34_2312 ();
 sg13g2_decap_8 FILLER_34_2340 ();
 sg13g2_decap_4 FILLER_34_2347 ();
 sg13g2_fill_1 FILLER_34_2351 ();
 sg13g2_decap_4 FILLER_34_2404 ();
 sg13g2_fill_1 FILLER_34_2408 ();
 sg13g2_fill_1 FILLER_34_2440 ();
 sg13g2_fill_2 FILLER_34_2446 ();
 sg13g2_fill_1 FILLER_34_2448 ();
 sg13g2_decap_4 FILLER_34_2453 ();
 sg13g2_fill_2 FILLER_34_2475 ();
 sg13g2_fill_2 FILLER_34_2485 ();
 sg13g2_fill_2 FILLER_34_2493 ();
 sg13g2_fill_1 FILLER_34_2526 ();
 sg13g2_fill_1 FILLER_34_2608 ();
 sg13g2_fill_2 FILLER_34_2615 ();
 sg13g2_decap_8 FILLER_34_2646 ();
 sg13g2_decap_8 FILLER_34_2653 ();
 sg13g2_decap_8 FILLER_34_2660 ();
 sg13g2_fill_2 FILLER_34_2667 ();
 sg13g2_fill_1 FILLER_34_2669 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_22 ();
 sg13g2_decap_8 FILLER_35_29 ();
 sg13g2_fill_2 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_38 ();
 sg13g2_decap_8 FILLER_35_59 ();
 sg13g2_fill_2 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_4 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_255 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_396 ();
 sg13g2_fill_1 FILLER_35_415 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_fill_1 FILLER_35_456 ();
 sg13g2_decap_4 FILLER_35_489 ();
 sg13g2_fill_2 FILLER_35_493 ();
 sg13g2_decap_4 FILLER_35_504 ();
 sg13g2_fill_1 FILLER_35_508 ();
 sg13g2_decap_4 FILLER_35_543 ();
 sg13g2_fill_1 FILLER_35_613 ();
 sg13g2_fill_1 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_624 ();
 sg13g2_fill_1 FILLER_35_633 ();
 sg13g2_fill_2 FILLER_35_655 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_fill_1 FILLER_35_700 ();
 sg13g2_fill_2 FILLER_35_706 ();
 sg13g2_fill_1 FILLER_35_708 ();
 sg13g2_decap_8 FILLER_35_720 ();
 sg13g2_decap_8 FILLER_35_727 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_decap_8 FILLER_35_745 ();
 sg13g2_fill_2 FILLER_35_752 ();
 sg13g2_fill_1 FILLER_35_754 ();
 sg13g2_fill_2 FILLER_35_767 ();
 sg13g2_fill_1 FILLER_35_769 ();
 sg13g2_decap_4 FILLER_35_775 ();
 sg13g2_fill_1 FILLER_35_779 ();
 sg13g2_fill_2 FILLER_35_855 ();
 sg13g2_fill_2 FILLER_35_870 ();
 sg13g2_fill_2 FILLER_35_898 ();
 sg13g2_fill_1 FILLER_35_907 ();
 sg13g2_fill_1 FILLER_35_956 ();
 sg13g2_fill_2 FILLER_35_982 ();
 sg13g2_fill_1 FILLER_35_1005 ();
 sg13g2_fill_1 FILLER_35_1029 ();
 sg13g2_fill_1 FILLER_35_1049 ();
 sg13g2_fill_1 FILLER_35_1055 ();
 sg13g2_fill_1 FILLER_35_1098 ();
 sg13g2_fill_2 FILLER_35_1108 ();
 sg13g2_fill_2 FILLER_35_1136 ();
 sg13g2_fill_1 FILLER_35_1142 ();
 sg13g2_fill_2 FILLER_35_1183 ();
 sg13g2_fill_2 FILLER_35_1237 ();
 sg13g2_fill_2 FILLER_35_1265 ();
 sg13g2_fill_1 FILLER_35_1283 ();
 sg13g2_fill_2 FILLER_35_1320 ();
 sg13g2_fill_1 FILLER_35_1370 ();
 sg13g2_fill_1 FILLER_35_1402 ();
 sg13g2_fill_1 FILLER_35_1463 ();
 sg13g2_fill_1 FILLER_35_1478 ();
 sg13g2_fill_2 FILLER_35_1504 ();
 sg13g2_fill_1 FILLER_35_1506 ();
 sg13g2_fill_1 FILLER_35_1511 ();
 sg13g2_decap_4 FILLER_35_1516 ();
 sg13g2_fill_1 FILLER_35_1520 ();
 sg13g2_fill_2 FILLER_35_1546 ();
 sg13g2_fill_1 FILLER_35_1552 ();
 sg13g2_fill_2 FILLER_35_1563 ();
 sg13g2_fill_1 FILLER_35_1565 ();
 sg13g2_decap_8 FILLER_35_1597 ();
 sg13g2_decap_8 FILLER_35_1604 ();
 sg13g2_fill_1 FILLER_35_1646 ();
 sg13g2_fill_2 FILLER_35_1684 ();
 sg13g2_fill_1 FILLER_35_1686 ();
 sg13g2_fill_2 FILLER_35_1695 ();
 sg13g2_fill_2 FILLER_35_1700 ();
 sg13g2_decap_4 FILLER_35_1706 ();
 sg13g2_fill_1 FILLER_35_1710 ();
 sg13g2_decap_8 FILLER_35_1716 ();
 sg13g2_fill_1 FILLER_35_1723 ();
 sg13g2_fill_2 FILLER_35_1737 ();
 sg13g2_fill_2 FILLER_35_1757 ();
 sg13g2_fill_1 FILLER_35_1759 ();
 sg13g2_decap_8 FILLER_35_1772 ();
 sg13g2_decap_8 FILLER_35_1779 ();
 sg13g2_decap_4 FILLER_35_1786 ();
 sg13g2_fill_1 FILLER_35_1790 ();
 sg13g2_fill_1 FILLER_35_1868 ();
 sg13g2_fill_1 FILLER_35_1908 ();
 sg13g2_fill_2 FILLER_35_1998 ();
 sg13g2_fill_2 FILLER_35_2005 ();
 sg13g2_fill_1 FILLER_35_2033 ();
 sg13g2_fill_1 FILLER_35_2044 ();
 sg13g2_decap_4 FILLER_35_2096 ();
 sg13g2_decap_8 FILLER_35_2117 ();
 sg13g2_decap_8 FILLER_35_2124 ();
 sg13g2_decap_8 FILLER_35_2131 ();
 sg13g2_decap_4 FILLER_35_2138 ();
 sg13g2_fill_2 FILLER_35_2142 ();
 sg13g2_decap_8 FILLER_35_2184 ();
 sg13g2_decap_8 FILLER_35_2191 ();
 sg13g2_decap_8 FILLER_35_2198 ();
 sg13g2_decap_8 FILLER_35_2205 ();
 sg13g2_decap_4 FILLER_35_2222 ();
 sg13g2_fill_2 FILLER_35_2226 ();
 sg13g2_decap_8 FILLER_35_2257 ();
 sg13g2_decap_8 FILLER_35_2264 ();
 sg13g2_fill_2 FILLER_35_2271 ();
 sg13g2_decap_8 FILLER_35_2277 ();
 sg13g2_fill_2 FILLER_35_2284 ();
 sg13g2_decap_4 FILLER_35_2295 ();
 sg13g2_decap_4 FILLER_35_2303 ();
 sg13g2_fill_2 FILLER_35_2317 ();
 sg13g2_fill_1 FILLER_35_2319 ();
 sg13g2_decap_8 FILLER_35_2324 ();
 sg13g2_decap_8 FILLER_35_2331 ();
 sg13g2_fill_1 FILLER_35_2377 ();
 sg13g2_fill_2 FILLER_35_2416 ();
 sg13g2_decap_8 FILLER_35_2448 ();
 sg13g2_decap_8 FILLER_35_2455 ();
 sg13g2_decap_8 FILLER_35_2462 ();
 sg13g2_fill_2 FILLER_35_2469 ();
 sg13g2_fill_1 FILLER_35_2471 ();
 sg13g2_fill_1 FILLER_35_2513 ();
 sg13g2_fill_2 FILLER_35_2582 ();
 sg13g2_fill_1 FILLER_35_2615 ();
 sg13g2_decap_8 FILLER_35_2646 ();
 sg13g2_decap_8 FILLER_35_2653 ();
 sg13g2_decap_8 FILLER_35_2660 ();
 sg13g2_fill_2 FILLER_35_2667 ();
 sg13g2_fill_1 FILLER_35_2669 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_397 ();
 sg13g2_fill_1 FILLER_36_419 ();
 sg13g2_fill_2 FILLER_36_454 ();
 sg13g2_fill_1 FILLER_36_456 ();
 sg13g2_fill_2 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_512 ();
 sg13g2_decap_4 FILLER_36_519 ();
 sg13g2_fill_1 FILLER_36_523 ();
 sg13g2_decap_4 FILLER_36_528 ();
 sg13g2_fill_1 FILLER_36_532 ();
 sg13g2_fill_1 FILLER_36_582 ();
 sg13g2_fill_1 FILLER_36_628 ();
 sg13g2_fill_1 FILLER_36_642 ();
 sg13g2_fill_1 FILLER_36_648 ();
 sg13g2_fill_2 FILLER_36_786 ();
 sg13g2_fill_1 FILLER_36_798 ();
 sg13g2_fill_1 FILLER_36_808 ();
 sg13g2_fill_1 FILLER_36_849 ();
 sg13g2_fill_1 FILLER_36_879 ();
 sg13g2_fill_2 FILLER_36_955 ();
 sg13g2_fill_2 FILLER_36_985 ();
 sg13g2_fill_2 FILLER_36_1000 ();
 sg13g2_fill_1 FILLER_36_1025 ();
 sg13g2_fill_1 FILLER_36_1029 ();
 sg13g2_fill_1 FILLER_36_1055 ();
 sg13g2_fill_2 FILLER_36_1099 ();
 sg13g2_fill_1 FILLER_36_1101 ();
 sg13g2_decap_4 FILLER_36_1107 ();
 sg13g2_fill_2 FILLER_36_1111 ();
 sg13g2_decap_8 FILLER_36_1122 ();
 sg13g2_decap_8 FILLER_36_1129 ();
 sg13g2_decap_8 FILLER_36_1136 ();
 sg13g2_fill_1 FILLER_36_1173 ();
 sg13g2_fill_1 FILLER_36_1206 ();
 sg13g2_fill_1 FILLER_36_1211 ();
 sg13g2_fill_2 FILLER_36_1236 ();
 sg13g2_fill_1 FILLER_36_1251 ();
 sg13g2_fill_2 FILLER_36_1303 ();
 sg13g2_fill_1 FILLER_36_1341 ();
 sg13g2_fill_2 FILLER_36_1399 ();
 sg13g2_fill_1 FILLER_36_1427 ();
 sg13g2_fill_2 FILLER_36_1507 ();
 sg13g2_fill_2 FILLER_36_1513 ();
 sg13g2_fill_2 FILLER_36_1520 ();
 sg13g2_decap_4 FILLER_36_1526 ();
 sg13g2_fill_2 FILLER_36_1534 ();
 sg13g2_fill_1 FILLER_36_1644 ();
 sg13g2_fill_1 FILLER_36_1652 ();
 sg13g2_fill_1 FILLER_36_1656 ();
 sg13g2_fill_1 FILLER_36_1663 ();
 sg13g2_fill_2 FILLER_36_1674 ();
 sg13g2_decap_4 FILLER_36_1688 ();
 sg13g2_fill_2 FILLER_36_1692 ();
 sg13g2_fill_2 FILLER_36_1706 ();
 sg13g2_decap_4 FILLER_36_1712 ();
 sg13g2_decap_8 FILLER_36_1724 ();
 sg13g2_fill_1 FILLER_36_1739 ();
 sg13g2_decap_8 FILLER_36_1771 ();
 sg13g2_decap_8 FILLER_36_1778 ();
 sg13g2_decap_8 FILLER_36_1785 ();
 sg13g2_decap_8 FILLER_36_1792 ();
 sg13g2_decap_8 FILLER_36_1799 ();
 sg13g2_decap_4 FILLER_36_1810 ();
 sg13g2_fill_2 FILLER_36_1822 ();
 sg13g2_fill_2 FILLER_36_1880 ();
 sg13g2_decap_8 FILLER_36_1929 ();
 sg13g2_fill_1 FILLER_36_1936 ();
 sg13g2_fill_1 FILLER_36_1979 ();
 sg13g2_decap_8 FILLER_36_2007 ();
 sg13g2_decap_4 FILLER_36_2052 ();
 sg13g2_fill_2 FILLER_36_2056 ();
 sg13g2_fill_2 FILLER_36_2088 ();
 sg13g2_fill_1 FILLER_36_2090 ();
 sg13g2_fill_2 FILLER_36_2101 ();
 sg13g2_fill_1 FILLER_36_2103 ();
 sg13g2_decap_4 FILLER_36_2114 ();
 sg13g2_fill_1 FILLER_36_2118 ();
 sg13g2_decap_8 FILLER_36_2129 ();
 sg13g2_fill_1 FILLER_36_2136 ();
 sg13g2_fill_2 FILLER_36_2173 ();
 sg13g2_fill_1 FILLER_36_2175 ();
 sg13g2_decap_4 FILLER_36_2179 ();
 sg13g2_fill_1 FILLER_36_2211 ();
 sg13g2_fill_2 FILLER_36_2219 ();
 sg13g2_fill_1 FILLER_36_2234 ();
 sg13g2_decap_8 FILLER_36_2261 ();
 sg13g2_fill_2 FILLER_36_2268 ();
 sg13g2_fill_1 FILLER_36_2270 ();
 sg13g2_fill_1 FILLER_36_2288 ();
 sg13g2_decap_8 FILLER_36_2310 ();
 sg13g2_decap_8 FILLER_36_2317 ();
 sg13g2_decap_8 FILLER_36_2324 ();
 sg13g2_decap_8 FILLER_36_2331 ();
 sg13g2_decap_8 FILLER_36_2338 ();
 sg13g2_decap_4 FILLER_36_2358 ();
 sg13g2_fill_2 FILLER_36_2372 ();
 sg13g2_fill_2 FILLER_36_2378 ();
 sg13g2_fill_2 FILLER_36_2384 ();
 sg13g2_fill_1 FILLER_36_2390 ();
 sg13g2_fill_2 FILLER_36_2425 ();
 sg13g2_fill_1 FILLER_36_2448 ();
 sg13g2_decap_8 FILLER_36_2456 ();
 sg13g2_fill_1 FILLER_36_2474 ();
 sg13g2_fill_1 FILLER_36_2507 ();
 sg13g2_fill_2 FILLER_36_2573 ();
 sg13g2_fill_1 FILLER_36_2634 ();
 sg13g2_decap_8 FILLER_36_2661 ();
 sg13g2_fill_2 FILLER_36_2668 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_2 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_78 ();
 sg13g2_decap_8 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_decap_8 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_decap_4 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_1 FILLER_37_409 ();
 sg13g2_fill_1 FILLER_37_423 ();
 sg13g2_fill_2 FILLER_37_450 ();
 sg13g2_fill_2 FILLER_37_457 ();
 sg13g2_decap_4 FILLER_37_471 ();
 sg13g2_fill_2 FILLER_37_497 ();
 sg13g2_fill_2 FILLER_37_514 ();
 sg13g2_fill_1 FILLER_37_516 ();
 sg13g2_decap_8 FILLER_37_543 ();
 sg13g2_decap_4 FILLER_37_550 ();
 sg13g2_fill_2 FILLER_37_554 ();
 sg13g2_decap_4 FILLER_37_570 ();
 sg13g2_fill_1 FILLER_37_590 ();
 sg13g2_fill_2 FILLER_37_596 ();
 sg13g2_fill_1 FILLER_37_607 ();
 sg13g2_fill_2 FILLER_37_617 ();
 sg13g2_fill_2 FILLER_37_645 ();
 sg13g2_fill_1 FILLER_37_659 ();
 sg13g2_fill_1 FILLER_37_669 ();
 sg13g2_fill_1 FILLER_37_678 ();
 sg13g2_fill_2 FILLER_37_684 ();
 sg13g2_fill_1 FILLER_37_720 ();
 sg13g2_fill_2 FILLER_37_778 ();
 sg13g2_fill_1 FILLER_37_780 ();
 sg13g2_fill_1 FILLER_37_786 ();
 sg13g2_fill_2 FILLER_37_813 ();
 sg13g2_fill_2 FILLER_37_825 ();
 sg13g2_fill_1 FILLER_37_843 ();
 sg13g2_fill_1 FILLER_37_871 ();
 sg13g2_fill_2 FILLER_37_888 ();
 sg13g2_fill_2 FILLER_37_905 ();
 sg13g2_fill_1 FILLER_37_929 ();
 sg13g2_fill_2 FILLER_37_943 ();
 sg13g2_fill_1 FILLER_37_991 ();
 sg13g2_fill_1 FILLER_37_1033 ();
 sg13g2_decap_4 FILLER_37_1088 ();
 sg13g2_fill_1 FILLER_37_1092 ();
 sg13g2_decap_4 FILLER_37_1133 ();
 sg13g2_fill_1 FILLER_37_1137 ();
 sg13g2_fill_2 FILLER_37_1148 ();
 sg13g2_fill_2 FILLER_37_1185 ();
 sg13g2_fill_1 FILLER_37_1187 ();
 sg13g2_decap_8 FILLER_37_1192 ();
 sg13g2_fill_1 FILLER_37_1199 ();
 sg13g2_fill_2 FILLER_37_1293 ();
 sg13g2_fill_1 FILLER_37_1364 ();
 sg13g2_fill_2 FILLER_37_1391 ();
 sg13g2_fill_2 FILLER_37_1429 ();
 sg13g2_fill_1 FILLER_37_1438 ();
 sg13g2_fill_1 FILLER_37_1470 ();
 sg13g2_fill_2 FILLER_37_1491 ();
 sg13g2_fill_2 FILLER_37_1516 ();
 sg13g2_fill_2 FILLER_37_1533 ();
 sg13g2_decap_8 FILLER_37_1543 ();
 sg13g2_decap_4 FILLER_37_1550 ();
 sg13g2_fill_1 FILLER_37_1554 ();
 sg13g2_decap_4 FILLER_37_1574 ();
 sg13g2_fill_2 FILLER_37_1578 ();
 sg13g2_fill_1 FILLER_37_1589 ();
 sg13g2_decap_4 FILLER_37_1603 ();
 sg13g2_fill_1 FILLER_37_1607 ();
 sg13g2_fill_1 FILLER_37_1613 ();
 sg13g2_fill_1 FILLER_37_1618 ();
 sg13g2_fill_1 FILLER_37_1623 ();
 sg13g2_fill_2 FILLER_37_1629 ();
 sg13g2_fill_1 FILLER_37_1644 ();
 sg13g2_decap_4 FILLER_37_1677 ();
 sg13g2_decap_4 FILLER_37_1689 ();
 sg13g2_fill_2 FILLER_37_1703 ();
 sg13g2_fill_1 FILLER_37_1705 ();
 sg13g2_decap_8 FILLER_37_1766 ();
 sg13g2_decap_8 FILLER_37_1773 ();
 sg13g2_decap_8 FILLER_37_1780 ();
 sg13g2_fill_2 FILLER_37_1787 ();
 sg13g2_decap_8 FILLER_37_1820 ();
 sg13g2_decap_4 FILLER_37_1827 ();
 sg13g2_decap_4 FILLER_37_1835 ();
 sg13g2_fill_1 FILLER_37_1839 ();
 sg13g2_fill_1 FILLER_37_1880 ();
 sg13g2_fill_2 FILLER_37_1924 ();
 sg13g2_fill_1 FILLER_37_1983 ();
 sg13g2_decap_8 FILLER_37_2018 ();
 sg13g2_decap_4 FILLER_37_2046 ();
 sg13g2_fill_1 FILLER_37_2050 ();
 sg13g2_fill_2 FILLER_37_2098 ();
 sg13g2_fill_1 FILLER_37_2179 ();
 sg13g2_fill_1 FILLER_37_2187 ();
 sg13g2_fill_1 FILLER_37_2198 ();
 sg13g2_fill_1 FILLER_37_2232 ();
 sg13g2_decap_8 FILLER_37_2247 ();
 sg13g2_fill_2 FILLER_37_2254 ();
 sg13g2_fill_1 FILLER_37_2256 ();
 sg13g2_fill_1 FILLER_37_2293 ();
 sg13g2_decap_8 FILLER_37_2330 ();
 sg13g2_decap_8 FILLER_37_2337 ();
 sg13g2_decap_8 FILLER_37_2344 ();
 sg13g2_decap_4 FILLER_37_2351 ();
 sg13g2_fill_2 FILLER_37_2355 ();
 sg13g2_fill_1 FILLER_37_2362 ();
 sg13g2_decap_8 FILLER_37_2371 ();
 sg13g2_decap_8 FILLER_37_2383 ();
 sg13g2_fill_1 FILLER_37_2390 ();
 sg13g2_fill_1 FILLER_37_2481 ();
 sg13g2_fill_1 FILLER_37_2515 ();
 sg13g2_fill_1 FILLER_37_2547 ();
 sg13g2_fill_1 FILLER_37_2553 ();
 sg13g2_fill_1 FILLER_37_2558 ();
 sg13g2_fill_2 FILLER_37_2564 ();
 sg13g2_fill_1 FILLER_37_2571 ();
 sg13g2_fill_2 FILLER_37_2602 ();
 sg13g2_decap_8 FILLER_37_2639 ();
 sg13g2_decap_8 FILLER_37_2646 ();
 sg13g2_decap_8 FILLER_37_2653 ();
 sg13g2_decap_8 FILLER_37_2660 ();
 sg13g2_fill_2 FILLER_37_2667 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_13 ();
 sg13g2_fill_2 FILLER_38_41 ();
 sg13g2_fill_1 FILLER_38_43 ();
 sg13g2_fill_2 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_103 ();
 sg13g2_fill_1 FILLER_38_105 ();
 sg13g2_decap_4 FILLER_38_110 ();
 sg13g2_decap_8 FILLER_38_121 ();
 sg13g2_decap_8 FILLER_38_128 ();
 sg13g2_decap_4 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_decap_4 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_decap_4 FILLER_38_313 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_329 ();
 sg13g2_fill_2 FILLER_38_372 ();
 sg13g2_fill_1 FILLER_38_378 ();
 sg13g2_fill_2 FILLER_38_392 ();
 sg13g2_fill_2 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_465 ();
 sg13g2_fill_2 FILLER_38_480 ();
 sg13g2_fill_1 FILLER_38_482 ();
 sg13g2_decap_8 FILLER_38_512 ();
 sg13g2_fill_1 FILLER_38_519 ();
 sg13g2_fill_1 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_577 ();
 sg13g2_decap_4 FILLER_38_583 ();
 sg13g2_fill_1 FILLER_38_618 ();
 sg13g2_fill_2 FILLER_38_654 ();
 sg13g2_fill_2 FILLER_38_661 ();
 sg13g2_fill_1 FILLER_38_663 ();
 sg13g2_fill_1 FILLER_38_669 ();
 sg13g2_fill_1 FILLER_38_675 ();
 sg13g2_fill_1 FILLER_38_681 ();
 sg13g2_fill_2 FILLER_38_687 ();
 sg13g2_fill_2 FILLER_38_697 ();
 sg13g2_fill_1 FILLER_38_703 ();
 sg13g2_fill_1 FILLER_38_726 ();
 sg13g2_fill_2 FILLER_38_828 ();
 sg13g2_fill_1 FILLER_38_837 ();
 sg13g2_fill_1 FILLER_38_842 ();
 sg13g2_fill_1 FILLER_38_851 ();
 sg13g2_fill_2 FILLER_38_893 ();
 sg13g2_fill_1 FILLER_38_979 ();
 sg13g2_fill_1 FILLER_38_1001 ();
 sg13g2_fill_2 FILLER_38_1029 ();
 sg13g2_fill_1 FILLER_38_1047 ();
 sg13g2_fill_1 FILLER_38_1074 ();
 sg13g2_decap_8 FILLER_38_1088 ();
 sg13g2_decap_4 FILLER_38_1095 ();
 sg13g2_fill_1 FILLER_38_1099 ();
 sg13g2_decap_4 FILLER_38_1104 ();
 sg13g2_fill_2 FILLER_38_1108 ();
 sg13g2_decap_8 FILLER_38_1114 ();
 sg13g2_decap_4 FILLER_38_1121 ();
 sg13g2_fill_1 FILLER_38_1125 ();
 sg13g2_decap_4 FILLER_38_1156 ();
 sg13g2_fill_1 FILLER_38_1160 ();
 sg13g2_fill_2 FILLER_38_1174 ();
 sg13g2_fill_1 FILLER_38_1176 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_fill_2 FILLER_38_1187 ();
 sg13g2_fill_1 FILLER_38_1189 ();
 sg13g2_decap_4 FILLER_38_1200 ();
 sg13g2_fill_1 FILLER_38_1204 ();
 sg13g2_fill_2 FILLER_38_1215 ();
 sg13g2_fill_2 FILLER_38_1224 ();
 sg13g2_fill_1 FILLER_38_1239 ();
 sg13g2_fill_1 FILLER_38_1281 ();
 sg13g2_fill_2 FILLER_38_1311 ();
 sg13g2_fill_1 FILLER_38_1320 ();
 sg13g2_decap_4 FILLER_38_1365 ();
 sg13g2_fill_1 FILLER_38_1369 ();
 sg13g2_decap_8 FILLER_38_1374 ();
 sg13g2_decap_8 FILLER_38_1381 ();
 sg13g2_decap_4 FILLER_38_1388 ();
 sg13g2_fill_1 FILLER_38_1396 ();
 sg13g2_fill_1 FILLER_38_1458 ();
 sg13g2_fill_1 FILLER_38_1516 ();
 sg13g2_fill_1 FILLER_38_1522 ();
 sg13g2_fill_1 FILLER_38_1527 ();
 sg13g2_fill_1 FILLER_38_1532 ();
 sg13g2_fill_1 FILLER_38_1550 ();
 sg13g2_fill_1 FILLER_38_1555 ();
 sg13g2_decap_8 FILLER_38_1570 ();
 sg13g2_fill_1 FILLER_38_1577 ();
 sg13g2_decap_4 FILLER_38_1587 ();
 sg13g2_fill_1 FILLER_38_1591 ();
 sg13g2_decap_8 FILLER_38_1601 ();
 sg13g2_decap_8 FILLER_38_1608 ();
 sg13g2_fill_2 FILLER_38_1620 ();
 sg13g2_fill_1 FILLER_38_1622 ();
 sg13g2_decap_4 FILLER_38_1641 ();
 sg13g2_fill_2 FILLER_38_1681 ();
 sg13g2_fill_2 FILLER_38_1687 ();
 sg13g2_fill_1 FILLER_38_1693 ();
 sg13g2_fill_2 FILLER_38_1712 ();
 sg13g2_decap_4 FILLER_38_1719 ();
 sg13g2_fill_1 FILLER_38_1723 ();
 sg13g2_fill_1 FILLER_38_1732 ();
 sg13g2_fill_1 FILLER_38_1736 ();
 sg13g2_decap_4 FILLER_38_1741 ();
 sg13g2_fill_1 FILLER_38_1745 ();
 sg13g2_decap_4 FILLER_38_1750 ();
 sg13g2_decap_4 FILLER_38_1759 ();
 sg13g2_decap_4 FILLER_38_1766 ();
 sg13g2_decap_8 FILLER_38_1782 ();
 sg13g2_decap_8 FILLER_38_1789 ();
 sg13g2_fill_2 FILLER_38_1796 ();
 sg13g2_fill_2 FILLER_38_1802 ();
 sg13g2_fill_2 FILLER_38_1809 ();
 sg13g2_fill_1 FILLER_38_1811 ();
 sg13g2_decap_4 FILLER_38_1825 ();
 sg13g2_fill_1 FILLER_38_1829 ();
 sg13g2_decap_8 FILLER_38_1834 ();
 sg13g2_decap_8 FILLER_38_1841 ();
 sg13g2_fill_2 FILLER_38_1848 ();
 sg13g2_fill_2 FILLER_38_1883 ();
 sg13g2_fill_1 FILLER_38_1888 ();
 sg13g2_fill_1 FILLER_38_1923 ();
 sg13g2_fill_2 FILLER_38_1942 ();
 sg13g2_fill_1 FILLER_38_1944 ();
 sg13g2_decap_4 FILLER_38_2023 ();
 sg13g2_fill_2 FILLER_38_2037 ();
 sg13g2_fill_1 FILLER_38_2039 ();
 sg13g2_fill_2 FILLER_38_2106 ();
 sg13g2_fill_2 FILLER_38_2171 ();
 sg13g2_decap_8 FILLER_38_2220 ();
 sg13g2_fill_1 FILLER_38_2227 ();
 sg13g2_decap_8 FILLER_38_2231 ();
 sg13g2_decap_4 FILLER_38_2238 ();
 sg13g2_fill_2 FILLER_38_2242 ();
 sg13g2_fill_2 FILLER_38_2301 ();
 sg13g2_decap_8 FILLER_38_2339 ();
 sg13g2_decap_8 FILLER_38_2346 ();
 sg13g2_fill_1 FILLER_38_2353 ();
 sg13g2_fill_1 FILLER_38_2385 ();
 sg13g2_fill_2 FILLER_38_2427 ();
 sg13g2_fill_1 FILLER_38_2492 ();
 sg13g2_fill_2 FILLER_38_2513 ();
 sg13g2_fill_1 FILLER_38_2538 ();
 sg13g2_fill_1 FILLER_38_2544 ();
 sg13g2_fill_1 FILLER_38_2585 ();
 sg13g2_fill_1 FILLER_38_2625 ();
 sg13g2_fill_2 FILLER_38_2631 ();
 sg13g2_decap_8 FILLER_38_2637 ();
 sg13g2_decap_8 FILLER_38_2644 ();
 sg13g2_decap_8 FILLER_38_2651 ();
 sg13g2_decap_8 FILLER_38_2658 ();
 sg13g2_decap_4 FILLER_38_2665 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_decap_4 FILLER_39_60 ();
 sg13g2_fill_2 FILLER_39_64 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_126 ();
 sg13g2_decap_4 FILLER_39_231 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_decap_4 FILLER_39_254 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_1 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_285 ();
 sg13g2_fill_2 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_342 ();
 sg13g2_fill_1 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_413 ();
 sg13g2_fill_1 FILLER_39_446 ();
 sg13g2_decap_4 FILLER_39_456 ();
 sg13g2_fill_1 FILLER_39_460 ();
 sg13g2_fill_1 FILLER_39_472 ();
 sg13g2_decap_8 FILLER_39_499 ();
 sg13g2_fill_2 FILLER_39_506 ();
 sg13g2_fill_1 FILLER_39_508 ();
 sg13g2_fill_2 FILLER_39_571 ();
 sg13g2_fill_1 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_579 ();
 sg13g2_fill_2 FILLER_39_586 ();
 sg13g2_fill_2 FILLER_39_592 ();
 sg13g2_fill_1 FILLER_39_594 ();
 sg13g2_fill_1 FILLER_39_600 ();
 sg13g2_fill_2 FILLER_39_606 ();
 sg13g2_fill_2 FILLER_39_664 ();
 sg13g2_fill_1 FILLER_39_686 ();
 sg13g2_fill_1 FILLER_39_697 ();
 sg13g2_fill_1 FILLER_39_708 ();
 sg13g2_decap_4 FILLER_39_735 ();
 sg13g2_fill_2 FILLER_39_744 ();
 sg13g2_fill_1 FILLER_39_746 ();
 sg13g2_fill_1 FILLER_39_831 ();
 sg13g2_fill_2 FILLER_39_837 ();
 sg13g2_fill_1 FILLER_39_847 ();
 sg13g2_fill_1 FILLER_39_865 ();
 sg13g2_fill_1 FILLER_39_880 ();
 sg13g2_fill_1 FILLER_39_940 ();
 sg13g2_fill_1 FILLER_39_947 ();
 sg13g2_fill_2 FILLER_39_956 ();
 sg13g2_fill_1 FILLER_39_966 ();
 sg13g2_fill_1 FILLER_39_1046 ();
 sg13g2_fill_1 FILLER_39_1073 ();
 sg13g2_fill_1 FILLER_39_1078 ();
 sg13g2_fill_2 FILLER_39_1109 ();
 sg13g2_fill_1 FILLER_39_1111 ();
 sg13g2_fill_1 FILLER_39_1138 ();
 sg13g2_fill_2 FILLER_39_1205 ();
 sg13g2_fill_1 FILLER_39_1223 ();
 sg13g2_fill_2 FILLER_39_1250 ();
 sg13g2_fill_2 FILLER_39_1266 ();
 sg13g2_fill_1 FILLER_39_1268 ();
 sg13g2_fill_1 FILLER_39_1301 ();
 sg13g2_fill_2 FILLER_39_1311 ();
 sg13g2_fill_1 FILLER_39_1325 ();
 sg13g2_decap_8 FILLER_39_1347 ();
 sg13g2_decap_8 FILLER_39_1390 ();
 sg13g2_decap_8 FILLER_39_1401 ();
 sg13g2_decap_8 FILLER_39_1414 ();
 sg13g2_decap_4 FILLER_39_1421 ();
 sg13g2_fill_1 FILLER_39_1425 ();
 sg13g2_decap_4 FILLER_39_1432 ();
 sg13g2_decap_8 FILLER_39_1452 ();
 sg13g2_fill_1 FILLER_39_1459 ();
 sg13g2_decap_4 FILLER_39_1465 ();
 sg13g2_decap_8 FILLER_39_1499 ();
 sg13g2_fill_1 FILLER_39_1506 ();
 sg13g2_fill_1 FILLER_39_1510 ();
 sg13g2_fill_1 FILLER_39_1555 ();
 sg13g2_decap_4 FILLER_39_1567 ();
 sg13g2_fill_1 FILLER_39_1576 ();
 sg13g2_fill_1 FILLER_39_1581 ();
 sg13g2_decap_4 FILLER_39_1587 ();
 sg13g2_fill_1 FILLER_39_1591 ();
 sg13g2_fill_1 FILLER_39_1609 ();
 sg13g2_decap_4 FILLER_39_1615 ();
 sg13g2_fill_2 FILLER_39_1623 ();
 sg13g2_fill_1 FILLER_39_1625 ();
 sg13g2_fill_1 FILLER_39_1630 ();
 sg13g2_fill_1 FILLER_39_1640 ();
 sg13g2_decap_8 FILLER_39_1694 ();
 sg13g2_decap_8 FILLER_39_1713 ();
 sg13g2_decap_8 FILLER_39_1720 ();
 sg13g2_decap_4 FILLER_39_1727 ();
 sg13g2_decap_8 FILLER_39_1735 ();
 sg13g2_fill_2 FILLER_39_1780 ();
 sg13g2_fill_1 FILLER_39_1782 ();
 sg13g2_decap_4 FILLER_39_1817 ();
 sg13g2_fill_1 FILLER_39_1821 ();
 sg13g2_fill_1 FILLER_39_1848 ();
 sg13g2_fill_1 FILLER_39_1879 ();
 sg13g2_decap_4 FILLER_39_1899 ();
 sg13g2_fill_1 FILLER_39_1903 ();
 sg13g2_fill_1 FILLER_39_1916 ();
 sg13g2_fill_1 FILLER_39_1930 ();
 sg13g2_fill_2 FILLER_39_1935 ();
 sg13g2_fill_1 FILLER_39_2002 ();
 sg13g2_fill_1 FILLER_39_2007 ();
 sg13g2_fill_1 FILLER_39_2034 ();
 sg13g2_fill_1 FILLER_39_2061 ();
 sg13g2_fill_1 FILLER_39_2066 ();
 sg13g2_decap_8 FILLER_39_2126 ();
 sg13g2_fill_2 FILLER_39_2143 ();
 sg13g2_decap_4 FILLER_39_2158 ();
 sg13g2_fill_1 FILLER_39_2162 ();
 sg13g2_fill_1 FILLER_39_2167 ();
 sg13g2_fill_2 FILLER_39_2293 ();
 sg13g2_fill_2 FILLER_39_2309 ();
 sg13g2_fill_2 FILLER_39_2341 ();
 sg13g2_decap_4 FILLER_39_2369 ();
 sg13g2_fill_2 FILLER_39_2383 ();
 sg13g2_fill_2 FILLER_39_2495 ();
 sg13g2_fill_1 FILLER_39_2528 ();
 sg13g2_fill_1 FILLER_39_2555 ();
 sg13g2_fill_2 FILLER_39_2587 ();
 sg13g2_fill_2 FILLER_39_2595 ();
 sg13g2_fill_2 FILLER_39_2624 ();
 sg13g2_decap_8 FILLER_39_2652 ();
 sg13g2_decap_8 FILLER_39_2659 ();
 sg13g2_decap_4 FILLER_39_2666 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_12 ();
 sg13g2_fill_1 FILLER_40_23 ();
 sg13g2_fill_1 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_45 ();
 sg13g2_decap_8 FILLER_40_52 ();
 sg13g2_fill_2 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_fill_2 FILLER_40_93 ();
 sg13g2_fill_1 FILLER_40_100 ();
 sg13g2_fill_2 FILLER_40_105 ();
 sg13g2_decap_4 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_160 ();
 sg13g2_fill_1 FILLER_40_188 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_fill_2 FILLER_40_222 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_decap_4 FILLER_40_261 ();
 sg13g2_decap_4 FILLER_40_269 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_fill_2 FILLER_40_279 ();
 sg13g2_decap_4 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_320 ();
 sg13g2_decap_4 FILLER_40_328 ();
 sg13g2_fill_1 FILLER_40_332 ();
 sg13g2_fill_2 FILLER_40_393 ();
 sg13g2_fill_2 FILLER_40_433 ();
 sg13g2_fill_2 FILLER_40_443 ();
 sg13g2_fill_1 FILLER_40_445 ();
 sg13g2_fill_2 FILLER_40_474 ();
 sg13g2_fill_1 FILLER_40_476 ();
 sg13g2_decap_4 FILLER_40_502 ();
 sg13g2_fill_1 FILLER_40_516 ();
 sg13g2_decap_4 FILLER_40_532 ();
 sg13g2_fill_2 FILLER_40_536 ();
 sg13g2_fill_2 FILLER_40_543 ();
 sg13g2_fill_1 FILLER_40_545 ();
 sg13g2_decap_8 FILLER_40_556 ();
 sg13g2_fill_1 FILLER_40_563 ();
 sg13g2_fill_2 FILLER_40_582 ();
 sg13g2_fill_1 FILLER_40_584 ();
 sg13g2_fill_2 FILLER_40_590 ();
 sg13g2_fill_1 FILLER_40_596 ();
 sg13g2_fill_2 FILLER_40_602 ();
 sg13g2_fill_2 FILLER_40_612 ();
 sg13g2_decap_8 FILLER_40_619 ();
 sg13g2_decap_8 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_647 ();
 sg13g2_decap_8 FILLER_40_654 ();
 sg13g2_decap_8 FILLER_40_661 ();
 sg13g2_fill_2 FILLER_40_692 ();
 sg13g2_fill_2 FILLER_40_699 ();
 sg13g2_fill_2 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_727 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_fill_1 FILLER_40_736 ();
 sg13g2_fill_2 FILLER_40_755 ();
 sg13g2_fill_1 FILLER_40_757 ();
 sg13g2_fill_2 FILLER_40_780 ();
 sg13g2_fill_1 FILLER_40_782 ();
 sg13g2_fill_1 FILLER_40_801 ();
 sg13g2_decap_4 FILLER_40_806 ();
 sg13g2_fill_2 FILLER_40_818 ();
 sg13g2_fill_2 FILLER_40_875 ();
 sg13g2_fill_2 FILLER_40_922 ();
 sg13g2_fill_1 FILLER_40_936 ();
 sg13g2_fill_2 FILLER_40_978 ();
 sg13g2_fill_1 FILLER_40_985 ();
 sg13g2_fill_1 FILLER_40_1076 ();
 sg13g2_fill_1 FILLER_40_1107 ();
 sg13g2_fill_1 FILLER_40_1118 ();
 sg13g2_fill_1 FILLER_40_1123 ();
 sg13g2_decap_8 FILLER_40_1134 ();
 sg13g2_decap_8 FILLER_40_1141 ();
 sg13g2_fill_1 FILLER_40_1148 ();
 sg13g2_decap_8 FILLER_40_1153 ();
 sg13g2_decap_8 FILLER_40_1196 ();
 sg13g2_fill_1 FILLER_40_1203 ();
 sg13g2_decap_4 FILLER_40_1238 ();
 sg13g2_fill_1 FILLER_40_1247 ();
 sg13g2_decap_4 FILLER_40_1258 ();
 sg13g2_fill_2 FILLER_40_1274 ();
 sg13g2_fill_1 FILLER_40_1276 ();
 sg13g2_fill_2 FILLER_40_1284 ();
 sg13g2_fill_1 FILLER_40_1290 ();
 sg13g2_fill_1 FILLER_40_1301 ();
 sg13g2_fill_1 FILLER_40_1348 ();
 sg13g2_decap_4 FILLER_40_1363 ();
 sg13g2_decap_8 FILLER_40_1375 ();
 sg13g2_fill_2 FILLER_40_1382 ();
 sg13g2_fill_1 FILLER_40_1384 ();
 sg13g2_decap_8 FILLER_40_1390 ();
 sg13g2_fill_2 FILLER_40_1397 ();
 sg13g2_decap_8 FILLER_40_1420 ();
 sg13g2_decap_8 FILLER_40_1427 ();
 sg13g2_decap_4 FILLER_40_1434 ();
 sg13g2_decap_8 FILLER_40_1446 ();
 sg13g2_decap_8 FILLER_40_1453 ();
 sg13g2_fill_2 FILLER_40_1460 ();
 sg13g2_fill_2 FILLER_40_1502 ();
 sg13g2_fill_1 FILLER_40_1504 ();
 sg13g2_fill_2 FILLER_40_1508 ();
 sg13g2_fill_2 FILLER_40_1516 ();
 sg13g2_fill_2 FILLER_40_1527 ();
 sg13g2_fill_2 FILLER_40_1533 ();
 sg13g2_fill_2 FILLER_40_1561 ();
 sg13g2_fill_1 FILLER_40_1563 ();
 sg13g2_decap_4 FILLER_40_1572 ();
 sg13g2_fill_2 FILLER_40_1576 ();
 sg13g2_decap_4 FILLER_40_1595 ();
 sg13g2_fill_1 FILLER_40_1599 ();
 sg13g2_fill_2 FILLER_40_1623 ();
 sg13g2_fill_1 FILLER_40_1629 ();
 sg13g2_fill_1 FILLER_40_1635 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1719 ();
 sg13g2_decap_8 FILLER_40_1726 ();
 sg13g2_decap_8 FILLER_40_1733 ();
 sg13g2_decap_4 FILLER_40_1740 ();
 sg13g2_fill_2 FILLER_40_1744 ();
 sg13g2_fill_2 FILLER_40_1843 ();
 sg13g2_fill_1 FILLER_40_1845 ();
 sg13g2_decap_4 FILLER_40_1855 ();
 sg13g2_fill_2 FILLER_40_1859 ();
 sg13g2_decap_8 FILLER_40_1900 ();
 sg13g2_decap_8 FILLER_40_1907 ();
 sg13g2_decap_4 FILLER_40_1914 ();
 sg13g2_fill_2 FILLER_40_1930 ();
 sg13g2_decap_8 FILLER_40_1962 ();
 sg13g2_decap_8 FILLER_40_1969 ();
 sg13g2_fill_2 FILLER_40_1976 ();
 sg13g2_fill_1 FILLER_40_1978 ();
 sg13g2_fill_2 FILLER_40_1987 ();
 sg13g2_fill_1 FILLER_40_1989 ();
 sg13g2_decap_4 FILLER_40_1994 ();
 sg13g2_fill_2 FILLER_40_1998 ();
 sg13g2_decap_4 FILLER_40_2010 ();
 sg13g2_fill_2 FILLER_40_2014 ();
 sg13g2_decap_4 FILLER_40_2020 ();
 sg13g2_fill_1 FILLER_40_2034 ();
 sg13g2_decap_4 FILLER_40_2121 ();
 sg13g2_decap_8 FILLER_40_2130 ();
 sg13g2_decap_4 FILLER_40_2137 ();
 sg13g2_fill_1 FILLER_40_2141 ();
 sg13g2_fill_2 FILLER_40_2176 ();
 sg13g2_fill_2 FILLER_40_2184 ();
 sg13g2_fill_2 FILLER_40_2237 ();
 sg13g2_decap_4 FILLER_40_2333 ();
 sg13g2_fill_2 FILLER_40_2337 ();
 sg13g2_fill_1 FILLER_40_2365 ();
 sg13g2_fill_2 FILLER_40_2375 ();
 sg13g2_fill_1 FILLER_40_2377 ();
 sg13g2_fill_2 FILLER_40_2384 ();
 sg13g2_fill_2 FILLER_40_2412 ();
 sg13g2_fill_1 FILLER_40_2414 ();
 sg13g2_fill_1 FILLER_40_2432 ();
 sg13g2_fill_2 FILLER_40_2516 ();
 sg13g2_fill_1 FILLER_40_2518 ();
 sg13g2_fill_2 FILLER_40_2545 ();
 sg13g2_fill_2 FILLER_40_2550 ();
 sg13g2_fill_2 FILLER_40_2578 ();
 sg13g2_fill_1 FILLER_40_2584 ();
 sg13g2_decap_8 FILLER_40_2640 ();
 sg13g2_decap_8 FILLER_40_2647 ();
 sg13g2_decap_8 FILLER_40_2654 ();
 sg13g2_decap_8 FILLER_40_2661 ();
 sg13g2_fill_2 FILLER_40_2668 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_18 ();
 sg13g2_decap_8 FILLER_41_60 ();
 sg13g2_fill_2 FILLER_41_67 ();
 sg13g2_fill_1 FILLER_41_69 ();
 sg13g2_fill_2 FILLER_41_93 ();
 sg13g2_decap_4 FILLER_41_121 ();
 sg13g2_fill_1 FILLER_41_151 ();
 sg13g2_fill_1 FILLER_41_169 ();
 sg13g2_decap_4 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_234 ();
 sg13g2_decap_8 FILLER_41_241 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_250 ();
 sg13g2_fill_2 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_267 ();
 sg13g2_fill_1 FILLER_41_269 ();
 sg13g2_fill_2 FILLER_41_305 ();
 sg13g2_decap_8 FILLER_41_327 ();
 sg13g2_decap_4 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_342 ();
 sg13g2_fill_2 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_351 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_396 ();
 sg13g2_decap_8 FILLER_41_414 ();
 sg13g2_decap_4 FILLER_41_421 ();
 sg13g2_fill_1 FILLER_41_472 ();
 sg13g2_decap_8 FILLER_41_486 ();
 sg13g2_decap_4 FILLER_41_493 ();
 sg13g2_fill_1 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_528 ();
 sg13g2_fill_1 FILLER_41_539 ();
 sg13g2_fill_2 FILLER_41_544 ();
 sg13g2_fill_1 FILLER_41_556 ();
 sg13g2_fill_2 FILLER_41_567 ();
 sg13g2_fill_1 FILLER_41_569 ();
 sg13g2_decap_8 FILLER_41_584 ();
 sg13g2_fill_2 FILLER_41_591 ();
 sg13g2_fill_1 FILLER_41_593 ();
 sg13g2_fill_2 FILLER_41_603 ();
 sg13g2_fill_1 FILLER_41_605 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_4 FILLER_41_637 ();
 sg13g2_fill_1 FILLER_41_641 ();
 sg13g2_decap_8 FILLER_41_646 ();
 sg13g2_decap_4 FILLER_41_653 ();
 sg13g2_fill_1 FILLER_41_657 ();
 sg13g2_decap_4 FILLER_41_663 ();
 sg13g2_fill_1 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_673 ();
 sg13g2_decap_8 FILLER_41_680 ();
 sg13g2_decap_8 FILLER_41_692 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_8 FILLER_41_738 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_fill_2 FILLER_41_768 ();
 sg13g2_fill_1 FILLER_41_774 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_fill_2 FILLER_41_815 ();
 sg13g2_fill_2 FILLER_41_822 ();
 sg13g2_fill_2 FILLER_41_827 ();
 sg13g2_decap_4 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_879 ();
 sg13g2_fill_2 FILLER_41_894 ();
 sg13g2_fill_1 FILLER_41_904 ();
 sg13g2_fill_1 FILLER_41_915 ();
 sg13g2_fill_1 FILLER_41_950 ();
 sg13g2_fill_2 FILLER_41_986 ();
 sg13g2_fill_2 FILLER_41_1076 ();
 sg13g2_fill_1 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1099 ();
 sg13g2_decap_4 FILLER_41_1106 ();
 sg13g2_fill_1 FILLER_41_1110 ();
 sg13g2_fill_2 FILLER_41_1121 ();
 sg13g2_decap_8 FILLER_41_1159 ();
 sg13g2_decap_8 FILLER_41_1166 ();
 sg13g2_decap_4 FILLER_41_1173 ();
 sg13g2_decap_8 FILLER_41_1181 ();
 sg13g2_decap_4 FILLER_41_1196 ();
 sg13g2_fill_1 FILLER_41_1200 ();
 sg13g2_fill_1 FILLER_41_1216 ();
 sg13g2_fill_1 FILLER_41_1230 ();
 sg13g2_fill_2 FILLER_41_1254 ();
 sg13g2_fill_1 FILLER_41_1261 ();
 sg13g2_fill_2 FILLER_41_1272 ();
 sg13g2_fill_2 FILLER_41_1290 ();
 sg13g2_fill_2 FILLER_41_1317 ();
 sg13g2_decap_4 FILLER_41_1333 ();
 sg13g2_fill_1 FILLER_41_1337 ();
 sg13g2_fill_1 FILLER_41_1344 ();
 sg13g2_fill_2 FILLER_41_1354 ();
 sg13g2_fill_1 FILLER_41_1356 ();
 sg13g2_decap_8 FILLER_41_1387 ();
 sg13g2_decap_4 FILLER_41_1394 ();
 sg13g2_decap_8 FILLER_41_1408 ();
 sg13g2_decap_8 FILLER_41_1415 ();
 sg13g2_decap_8 FILLER_41_1422 ();
 sg13g2_fill_2 FILLER_41_1438 ();
 sg13g2_decap_8 FILLER_41_1444 ();
 sg13g2_fill_1 FILLER_41_1451 ();
 sg13g2_decap_4 FILLER_41_1459 ();
 sg13g2_fill_2 FILLER_41_1472 ();
 sg13g2_decap_4 FILLER_41_1505 ();
 sg13g2_fill_1 FILLER_41_1509 ();
 sg13g2_fill_2 FILLER_41_1514 ();
 sg13g2_fill_2 FILLER_41_1528 ();
 sg13g2_fill_1 FILLER_41_1530 ();
 sg13g2_decap_4 FILLER_41_1534 ();
 sg13g2_decap_4 FILLER_41_1610 ();
 sg13g2_fill_2 FILLER_41_1614 ();
 sg13g2_fill_1 FILLER_41_1620 ();
 sg13g2_fill_2 FILLER_41_1626 ();
 sg13g2_fill_2 FILLER_41_1633 ();
 sg13g2_fill_1 FILLER_41_1639 ();
 sg13g2_fill_1 FILLER_41_1659 ();
 sg13g2_fill_1 FILLER_41_1691 ();
 sg13g2_decap_8 FILLER_41_1718 ();
 sg13g2_decap_8 FILLER_41_1725 ();
 sg13g2_decap_8 FILLER_41_1732 ();
 sg13g2_fill_2 FILLER_41_1739 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_fill_2 FILLER_41_1781 ();
 sg13g2_fill_2 FILLER_41_1809 ();
 sg13g2_fill_1 FILLER_41_1811 ();
 sg13g2_fill_1 FILLER_41_1820 ();
 sg13g2_fill_2 FILLER_41_1825 ();
 sg13g2_fill_2 FILLER_41_1831 ();
 sg13g2_decap_8 FILLER_41_1838 ();
 sg13g2_decap_8 FILLER_41_1845 ();
 sg13g2_fill_2 FILLER_41_1852 ();
 sg13g2_fill_1 FILLER_41_1854 ();
 sg13g2_fill_2 FILLER_41_1870 ();
 sg13g2_fill_1 FILLER_41_1872 ();
 sg13g2_fill_2 FILLER_41_1878 ();
 sg13g2_fill_2 FILLER_41_1921 ();
 sg13g2_fill_2 FILLER_41_1936 ();
 sg13g2_fill_1 FILLER_41_1938 ();
 sg13g2_fill_2 FILLER_41_1950 ();
 sg13g2_decap_8 FILLER_41_1960 ();
 sg13g2_decap_8 FILLER_41_1967 ();
 sg13g2_decap_8 FILLER_41_1974 ();
 sg13g2_fill_1 FILLER_41_1981 ();
 sg13g2_decap_8 FILLER_41_2018 ();
 sg13g2_decap_8 FILLER_41_2025 ();
 sg13g2_decap_4 FILLER_41_2042 ();
 sg13g2_fill_1 FILLER_41_2050 ();
 sg13g2_fill_1 FILLER_41_2083 ();
 sg13g2_fill_1 FILLER_41_2107 ();
 sg13g2_decap_8 FILLER_41_2141 ();
 sg13g2_fill_1 FILLER_41_2148 ();
 sg13g2_decap_4 FILLER_41_2175 ();
 sg13g2_fill_2 FILLER_41_2179 ();
 sg13g2_decap_4 FILLER_41_2184 ();
 sg13g2_fill_2 FILLER_41_2188 ();
 sg13g2_fill_2 FILLER_41_2207 ();
 sg13g2_fill_1 FILLER_41_2215 ();
 sg13g2_decap_4 FILLER_41_2248 ();
 sg13g2_fill_1 FILLER_41_2252 ();
 sg13g2_fill_2 FILLER_41_2257 ();
 sg13g2_fill_2 FILLER_41_2270 ();
 sg13g2_decap_8 FILLER_41_2319 ();
 sg13g2_decap_4 FILLER_41_2326 ();
 sg13g2_fill_1 FILLER_41_2330 ();
 sg13g2_fill_2 FILLER_41_2372 ();
 sg13g2_fill_1 FILLER_41_2374 ();
 sg13g2_decap_4 FILLER_41_2380 ();
 sg13g2_fill_1 FILLER_41_2423 ();
 sg13g2_fill_1 FILLER_41_2433 ();
 sg13g2_fill_1 FILLER_41_2450 ();
 sg13g2_fill_2 FILLER_41_2470 ();
 sg13g2_fill_1 FILLER_41_2530 ();
 sg13g2_fill_2 FILLER_41_2535 ();
 sg13g2_fill_2 FILLER_41_2541 ();
 sg13g2_fill_1 FILLER_41_2543 ();
 sg13g2_fill_2 FILLER_41_2561 ();
 sg13g2_fill_1 FILLER_41_2563 ();
 sg13g2_fill_1 FILLER_41_2570 ();
 sg13g2_fill_1 FILLER_41_2600 ();
 sg13g2_decap_8 FILLER_41_2631 ();
 sg13g2_decap_8 FILLER_41_2638 ();
 sg13g2_decap_8 FILLER_41_2645 ();
 sg13g2_decap_8 FILLER_41_2652 ();
 sg13g2_decap_8 FILLER_41_2659 ();
 sg13g2_decap_4 FILLER_41_2666 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_30 ();
 sg13g2_fill_2 FILLER_42_92 ();
 sg13g2_fill_1 FILLER_42_94 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_fill_2 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_114 ();
 sg13g2_fill_2 FILLER_42_120 ();
 sg13g2_fill_1 FILLER_42_122 ();
 sg13g2_fill_2 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_133 ();
 sg13g2_fill_2 FILLER_42_140 ();
 sg13g2_fill_2 FILLER_42_160 ();
 sg13g2_fill_1 FILLER_42_162 ();
 sg13g2_fill_2 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_177 ();
 sg13g2_fill_2 FILLER_42_185 ();
 sg13g2_fill_1 FILLER_42_187 ();
 sg13g2_fill_2 FILLER_42_197 ();
 sg13g2_fill_1 FILLER_42_199 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_4 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_221 ();
 sg13g2_decap_8 FILLER_42_256 ();
 sg13g2_fill_2 FILLER_42_263 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_fill_1 FILLER_42_287 ();
 sg13g2_fill_2 FILLER_42_291 ();
 sg13g2_fill_2 FILLER_42_297 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_fill_1 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_341 ();
 sg13g2_decap_4 FILLER_42_348 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_fill_1 FILLER_42_389 ();
 sg13g2_fill_1 FILLER_42_426 ();
 sg13g2_fill_2 FILLER_42_432 ();
 sg13g2_fill_1 FILLER_42_434 ();
 sg13g2_fill_1 FILLER_42_461 ();
 sg13g2_fill_1 FILLER_42_499 ();
 sg13g2_decap_8 FILLER_42_585 ();
 sg13g2_decap_8 FILLER_42_592 ();
 sg13g2_decap_8 FILLER_42_599 ();
 sg13g2_fill_2 FILLER_42_606 ();
 sg13g2_fill_1 FILLER_42_608 ();
 sg13g2_decap_8 FILLER_42_617 ();
 sg13g2_decap_4 FILLER_42_624 ();
 sg13g2_fill_2 FILLER_42_633 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_8 FILLER_42_678 ();
 sg13g2_fill_1 FILLER_42_719 ();
 sg13g2_fill_2 FILLER_42_730 ();
 sg13g2_fill_1 FILLER_42_732 ();
 sg13g2_fill_2 FILLER_42_738 ();
 sg13g2_fill_1 FILLER_42_740 ();
 sg13g2_fill_1 FILLER_42_759 ();
 sg13g2_fill_2 FILLER_42_770 ();
 sg13g2_fill_1 FILLER_42_772 ();
 sg13g2_fill_1 FILLER_42_778 ();
 sg13g2_decap_4 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_824 ();
 sg13g2_decap_4 FILLER_42_831 ();
 sg13g2_fill_1 FILLER_42_835 ();
 sg13g2_decap_4 FILLER_42_844 ();
 sg13g2_fill_2 FILLER_42_848 ();
 sg13g2_fill_1 FILLER_42_864 ();
 sg13g2_fill_1 FILLER_42_955 ();
 sg13g2_fill_1 FILLER_42_960 ();
 sg13g2_fill_2 FILLER_42_971 ();
 sg13g2_fill_1 FILLER_42_1006 ();
 sg13g2_fill_1 FILLER_42_1038 ();
 sg13g2_decap_8 FILLER_42_1043 ();
 sg13g2_fill_2 FILLER_42_1050 ();
 sg13g2_decap_8 FILLER_42_1088 ();
 sg13g2_decap_8 FILLER_42_1095 ();
 sg13g2_decap_8 FILLER_42_1128 ();
 sg13g2_decap_8 FILLER_42_1161 ();
 sg13g2_fill_1 FILLER_42_1175 ();
 sg13g2_fill_2 FILLER_42_1189 ();
 sg13g2_fill_1 FILLER_42_1191 ();
 sg13g2_fill_1 FILLER_42_1228 ();
 sg13g2_fill_1 FILLER_42_1262 ();
 sg13g2_fill_1 FILLER_42_1267 ();
 sg13g2_fill_1 FILLER_42_1295 ();
 sg13g2_decap_8 FILLER_42_1340 ();
 sg13g2_fill_1 FILLER_42_1354 ();
 sg13g2_fill_2 FILLER_42_1366 ();
 sg13g2_decap_4 FILLER_42_1379 ();
 sg13g2_fill_1 FILLER_42_1383 ();
 sg13g2_fill_2 FILLER_42_1390 ();
 sg13g2_fill_1 FILLER_42_1392 ();
 sg13g2_fill_1 FILLER_42_1492 ();
 sg13g2_fill_2 FILLER_42_1534 ();
 sg13g2_fill_1 FILLER_42_1546 ();
 sg13g2_fill_2 FILLER_42_1556 ();
 sg13g2_fill_2 FILLER_42_1563 ();
 sg13g2_fill_1 FILLER_42_1565 ();
 sg13g2_fill_2 FILLER_42_1582 ();
 sg13g2_fill_1 FILLER_42_1597 ();
 sg13g2_fill_1 FILLER_42_1609 ();
 sg13g2_fill_1 FILLER_42_1615 ();
 sg13g2_fill_1 FILLER_42_1623 ();
 sg13g2_fill_1 FILLER_42_1628 ();
 sg13g2_fill_1 FILLER_42_1634 ();
 sg13g2_fill_1 FILLER_42_1640 ();
 sg13g2_fill_2 FILLER_42_1654 ();
 sg13g2_fill_1 FILLER_42_1656 ();
 sg13g2_decap_8 FILLER_42_1687 ();
 sg13g2_decap_4 FILLER_42_1694 ();
 sg13g2_decap_4 FILLER_42_1702 ();
 sg13g2_fill_2 FILLER_42_1712 ();
 sg13g2_fill_2 FILLER_42_1724 ();
 sg13g2_fill_1 FILLER_42_1726 ();
 sg13g2_decap_4 FILLER_42_1732 ();
 sg13g2_fill_2 FILLER_42_1744 ();
 sg13g2_fill_1 FILLER_42_1773 ();
 sg13g2_decap_4 FILLER_42_1787 ();
 sg13g2_fill_1 FILLER_42_1791 ();
 sg13g2_fill_2 FILLER_42_1796 ();
 sg13g2_fill_1 FILLER_42_1798 ();
 sg13g2_decap_4 FILLER_42_1803 ();
 sg13g2_fill_2 FILLER_42_1807 ();
 sg13g2_decap_4 FILLER_42_1843 ();
 sg13g2_decap_8 FILLER_42_1850 ();
 sg13g2_decap_8 FILLER_42_1861 ();
 sg13g2_fill_1 FILLER_42_1868 ();
 sg13g2_fill_2 FILLER_42_1880 ();
 sg13g2_fill_2 FILLER_42_1919 ();
 sg13g2_fill_1 FILLER_42_1921 ();
 sg13g2_fill_2 FILLER_42_1948 ();
 sg13g2_decap_4 FILLER_42_1980 ();
 sg13g2_fill_2 FILLER_42_1984 ();
 sg13g2_fill_2 FILLER_42_1996 ();
 sg13g2_fill_1 FILLER_42_1998 ();
 sg13g2_fill_2 FILLER_42_2003 ();
 sg13g2_fill_1 FILLER_42_2005 ();
 sg13g2_decap_8 FILLER_42_2010 ();
 sg13g2_decap_4 FILLER_42_2017 ();
 sg13g2_fill_1 FILLER_42_2021 ();
 sg13g2_decap_8 FILLER_42_2026 ();
 sg13g2_decap_4 FILLER_42_2033 ();
 sg13g2_fill_1 FILLER_42_2037 ();
 sg13g2_decap_4 FILLER_42_2052 ();
 sg13g2_fill_1 FILLER_42_2056 ();
 sg13g2_fill_1 FILLER_42_2096 ();
 sg13g2_fill_1 FILLER_42_2104 ();
 sg13g2_fill_1 FILLER_42_2141 ();
 sg13g2_fill_2 FILLER_42_2152 ();
 sg13g2_fill_2 FILLER_42_2158 ();
 sg13g2_decap_8 FILLER_42_2254 ();
 sg13g2_fill_1 FILLER_42_2261 ();
 sg13g2_fill_1 FILLER_42_2297 ();
 sg13g2_decap_8 FILLER_42_2336 ();
 sg13g2_decap_8 FILLER_42_2347 ();
 sg13g2_decap_4 FILLER_42_2358 ();
 sg13g2_fill_2 FILLER_42_2370 ();
 sg13g2_fill_1 FILLER_42_2372 ();
 sg13g2_decap_4 FILLER_42_2387 ();
 sg13g2_decap_4 FILLER_42_2395 ();
 sg13g2_fill_2 FILLER_42_2410 ();
 sg13g2_fill_1 FILLER_42_2449 ();
 sg13g2_fill_1 FILLER_42_2467 ();
 sg13g2_fill_2 FILLER_42_2473 ();
 sg13g2_fill_1 FILLER_42_2501 ();
 sg13g2_fill_2 FILLER_42_2507 ();
 sg13g2_decap_8 FILLER_42_2515 ();
 sg13g2_decap_8 FILLER_42_2532 ();
 sg13g2_decap_4 FILLER_42_2539 ();
 sg13g2_fill_2 FILLER_42_2561 ();
 sg13g2_fill_1 FILLER_42_2589 ();
 sg13g2_fill_2 FILLER_42_2595 ();
 sg13g2_decap_8 FILLER_42_2629 ();
 sg13g2_decap_8 FILLER_42_2636 ();
 sg13g2_decap_8 FILLER_42_2643 ();
 sg13g2_decap_8 FILLER_42_2650 ();
 sg13g2_decap_8 FILLER_42_2657 ();
 sg13g2_decap_4 FILLER_42_2664 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_4 ();
 sg13g2_fill_1 FILLER_43_10 ();
 sg13g2_fill_2 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_33 ();
 sg13g2_decap_8 FILLER_43_61 ();
 sg13g2_decap_8 FILLER_43_68 ();
 sg13g2_fill_2 FILLER_43_75 ();
 sg13g2_fill_2 FILLER_43_87 ();
 sg13g2_fill_1 FILLER_43_89 ();
 sg13g2_decap_4 FILLER_43_94 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_decap_4 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_235 ();
 sg13g2_fill_2 FILLER_43_243 ();
 sg13g2_decap_8 FILLER_43_253 ();
 sg13g2_decap_8 FILLER_43_260 ();
 sg13g2_decap_8 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_360 ();
 sg13g2_fill_1 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_367 ();
 sg13g2_fill_2 FILLER_43_374 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_2 FILLER_43_402 ();
 sg13g2_fill_1 FILLER_43_410 ();
 sg13g2_fill_1 FILLER_43_426 ();
 sg13g2_fill_2 FILLER_43_437 ();
 sg13g2_fill_1 FILLER_43_443 ();
 sg13g2_fill_1 FILLER_43_448 ();
 sg13g2_fill_1 FILLER_43_454 ();
 sg13g2_fill_1 FILLER_43_460 ();
 sg13g2_decap_8 FILLER_43_500 ();
 sg13g2_fill_2 FILLER_43_507 ();
 sg13g2_fill_1 FILLER_43_540 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_fill_2 FILLER_43_588 ();
 sg13g2_fill_2 FILLER_43_603 ();
 sg13g2_fill_1 FILLER_43_605 ();
 sg13g2_fill_1 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_627 ();
 sg13g2_fill_2 FILLER_43_685 ();
 sg13g2_fill_2 FILLER_43_724 ();
 sg13g2_fill_1 FILLER_43_736 ();
 sg13g2_fill_2 FILLER_43_780 ();
 sg13g2_fill_1 FILLER_43_805 ();
 sg13g2_fill_1 FILLER_43_836 ();
 sg13g2_fill_2 FILLER_43_863 ();
 sg13g2_fill_1 FILLER_43_869 ();
 sg13g2_fill_1 FILLER_43_880 ();
 sg13g2_fill_2 FILLER_43_889 ();
 sg13g2_fill_2 FILLER_43_895 ();
 sg13g2_fill_1 FILLER_43_901 ();
 sg13g2_fill_1 FILLER_43_928 ();
 sg13g2_fill_1 FILLER_43_978 ();
 sg13g2_fill_1 FILLER_43_1016 ();
 sg13g2_decap_8 FILLER_43_1027 ();
 sg13g2_decap_8 FILLER_43_1034 ();
 sg13g2_decap_8 FILLER_43_1041 ();
 sg13g2_decap_8 FILLER_43_1048 ();
 sg13g2_fill_2 FILLER_43_1055 ();
 sg13g2_fill_1 FILLER_43_1057 ();
 sg13g2_fill_1 FILLER_43_1068 ();
 sg13g2_decap_4 FILLER_43_1073 ();
 sg13g2_decap_8 FILLER_43_1113 ();
 sg13g2_decap_4 FILLER_43_1124 ();
 sg13g2_fill_1 FILLER_43_1128 ();
 sg13g2_fill_1 FILLER_43_1139 ();
 sg13g2_decap_8 FILLER_43_1148 ();
 sg13g2_decap_4 FILLER_43_1195 ();
 sg13g2_decap_4 FILLER_43_1203 ();
 sg13g2_fill_2 FILLER_43_1212 ();
 sg13g2_decap_4 FILLER_43_1218 ();
 sg13g2_fill_2 FILLER_43_1242 ();
 sg13g2_fill_1 FILLER_43_1280 ();
 sg13g2_decap_4 FILLER_43_1340 ();
 sg13g2_fill_1 FILLER_43_1359 ();
 sg13g2_fill_2 FILLER_43_1370 ();
 sg13g2_fill_1 FILLER_43_1387 ();
 sg13g2_fill_2 FILLER_43_1398 ();
 sg13g2_fill_1 FILLER_43_1400 ();
 sg13g2_fill_2 FILLER_43_1469 ();
 sg13g2_fill_1 FILLER_43_1488 ();
 sg13g2_fill_1 FILLER_43_1525 ();
 sg13g2_decap_8 FILLER_43_1572 ();
 sg13g2_decap_8 FILLER_43_1628 ();
 sg13g2_decap_4 FILLER_43_1635 ();
 sg13g2_fill_2 FILLER_43_1639 ();
 sg13g2_decap_8 FILLER_43_1645 ();
 sg13g2_decap_8 FILLER_43_1652 ();
 sg13g2_decap_8 FILLER_43_1659 ();
 sg13g2_decap_8 FILLER_43_1666 ();
 sg13g2_decap_8 FILLER_43_1681 ();
 sg13g2_decap_8 FILLER_43_1688 ();
 sg13g2_decap_8 FILLER_43_1695 ();
 sg13g2_decap_8 FILLER_43_1702 ();
 sg13g2_fill_2 FILLER_43_1709 ();
 sg13g2_fill_1 FILLER_43_1711 ();
 sg13g2_fill_2 FILLER_43_1720 ();
 sg13g2_fill_1 FILLER_43_1756 ();
 sg13g2_decap_8 FILLER_43_1797 ();
 sg13g2_decap_8 FILLER_43_1804 ();
 sg13g2_decap_8 FILLER_43_1811 ();
 sg13g2_decap_8 FILLER_43_1818 ();
 sg13g2_decap_8 FILLER_43_1829 ();
 sg13g2_decap_8 FILLER_43_1836 ();
 sg13g2_fill_2 FILLER_43_1843 ();
 sg13g2_decap_8 FILLER_43_1850 ();
 sg13g2_decap_4 FILLER_43_1857 ();
 sg13g2_fill_1 FILLER_43_1861 ();
 sg13g2_fill_2 FILLER_43_1871 ();
 sg13g2_fill_1 FILLER_43_1873 ();
 sg13g2_decap_4 FILLER_43_1879 ();
 sg13g2_fill_1 FILLER_43_1913 ();
 sg13g2_fill_1 FILLER_43_1918 ();
 sg13g2_fill_2 FILLER_43_1923 ();
 sg13g2_fill_2 FILLER_43_1951 ();
 sg13g2_fill_1 FILLER_43_1953 ();
 sg13g2_fill_1 FILLER_43_1964 ();
 sg13g2_fill_1 FILLER_43_1978 ();
 sg13g2_fill_1 FILLER_43_2041 ();
 sg13g2_fill_1 FILLER_43_2063 ();
 sg13g2_fill_2 FILLER_43_2103 ();
 sg13g2_fill_2 FILLER_43_2135 ();
 sg13g2_fill_1 FILLER_43_2137 ();
 sg13g2_decap_4 FILLER_43_2178 ();
 sg13g2_fill_1 FILLER_43_2182 ();
 sg13g2_decap_8 FILLER_43_2248 ();
 sg13g2_fill_1 FILLER_43_2267 ();
 sg13g2_fill_2 FILLER_43_2274 ();
 sg13g2_fill_2 FILLER_43_2286 ();
 sg13g2_decap_4 FILLER_43_2291 ();
 sg13g2_fill_1 FILLER_43_2295 ();
 sg13g2_decap_8 FILLER_43_2326 ();
 sg13g2_decap_8 FILLER_43_2333 ();
 sg13g2_decap_8 FILLER_43_2340 ();
 sg13g2_fill_1 FILLER_43_2347 ();
 sg13g2_fill_1 FILLER_43_2352 ();
 sg13g2_fill_2 FILLER_43_2388 ();
 sg13g2_fill_1 FILLER_43_2390 ();
 sg13g2_fill_1 FILLER_43_2436 ();
 sg13g2_fill_2 FILLER_43_2443 ();
 sg13g2_fill_1 FILLER_43_2452 ();
 sg13g2_fill_2 FILLER_43_2481 ();
 sg13g2_fill_2 FILLER_43_2509 ();
 sg13g2_fill_2 FILLER_43_2531 ();
 sg13g2_fill_2 FILLER_43_2537 ();
 sg13g2_fill_1 FILLER_43_2539 ();
 sg13g2_fill_2 FILLER_43_2544 ();
 sg13g2_fill_1 FILLER_43_2546 ();
 sg13g2_fill_2 FILLER_43_2585 ();
 sg13g2_fill_1 FILLER_43_2596 ();
 sg13g2_decap_8 FILLER_43_2601 ();
 sg13g2_fill_2 FILLER_43_2608 ();
 sg13g2_decap_8 FILLER_43_2618 ();
 sg13g2_decap_8 FILLER_43_2625 ();
 sg13g2_decap_8 FILLER_43_2632 ();
 sg13g2_decap_8 FILLER_43_2639 ();
 sg13g2_decap_8 FILLER_43_2646 ();
 sg13g2_decap_8 FILLER_43_2653 ();
 sg13g2_decap_8 FILLER_43_2660 ();
 sg13g2_fill_2 FILLER_43_2667 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_fill_1 FILLER_44_78 ();
 sg13g2_decap_4 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_118 ();
 sg13g2_decap_4 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_129 ();
 sg13g2_decap_8 FILLER_44_186 ();
 sg13g2_fill_2 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_fill_2 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_254 ();
 sg13g2_fill_2 FILLER_44_261 ();
 sg13g2_decap_4 FILLER_44_268 ();
 sg13g2_fill_1 FILLER_44_276 ();
 sg13g2_fill_1 FILLER_44_300 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_fill_1 FILLER_44_328 ();
 sg13g2_fill_1 FILLER_44_338 ();
 sg13g2_decap_4 FILLER_44_349 ();
 sg13g2_decap_4 FILLER_44_357 ();
 sg13g2_fill_1 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_44_416 ();
 sg13g2_fill_1 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_44_446 ();
 sg13g2_decap_8 FILLER_44_453 ();
 sg13g2_decap_8 FILLER_44_460 ();
 sg13g2_fill_2 FILLER_44_467 ();
 sg13g2_fill_1 FILLER_44_488 ();
 sg13g2_decap_8 FILLER_44_500 ();
 sg13g2_fill_1 FILLER_44_507 ();
 sg13g2_fill_1 FILLER_44_525 ();
 sg13g2_decap_8 FILLER_44_540 ();
 sg13g2_decap_8 FILLER_44_547 ();
 sg13g2_fill_1 FILLER_44_554 ();
 sg13g2_fill_2 FILLER_44_582 ();
 sg13g2_fill_1 FILLER_44_588 ();
 sg13g2_fill_1 FILLER_44_619 ();
 sg13g2_decap_4 FILLER_44_656 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_4 FILLER_44_686 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_fill_2 FILLER_44_700 ();
 sg13g2_decap_4 FILLER_44_766 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_4 FILLER_44_782 ();
 sg13g2_fill_2 FILLER_44_795 ();
 sg13g2_fill_1 FILLER_44_797 ();
 sg13g2_fill_2 FILLER_44_849 ();
 sg13g2_fill_2 FILLER_44_877 ();
 sg13g2_fill_1 FILLER_44_879 ();
 sg13g2_fill_1 FILLER_44_890 ();
 sg13g2_fill_1 FILLER_44_908 ();
 sg13g2_fill_2 FILLER_44_926 ();
 sg13g2_fill_1 FILLER_44_938 ();
 sg13g2_fill_2 FILLER_44_947 ();
 sg13g2_fill_2 FILLER_44_964 ();
 sg13g2_fill_1 FILLER_44_1016 ();
 sg13g2_decap_8 FILLER_44_1034 ();
 sg13g2_decap_8 FILLER_44_1041 ();
 sg13g2_decap_8 FILLER_44_1048 ();
 sg13g2_decap_8 FILLER_44_1055 ();
 sg13g2_decap_8 FILLER_44_1062 ();
 sg13g2_fill_2 FILLER_44_1069 ();
 sg13g2_fill_2 FILLER_44_1078 ();
 sg13g2_fill_1 FILLER_44_1080 ();
 sg13g2_fill_2 FILLER_44_1098 ();
 sg13g2_fill_1 FILLER_44_1100 ();
 sg13g2_fill_2 FILLER_44_1111 ();
 sg13g2_decap_4 FILLER_44_1139 ();
 sg13g2_fill_2 FILLER_44_1143 ();
 sg13g2_decap_8 FILLER_44_1149 ();
 sg13g2_fill_2 FILLER_44_1156 ();
 sg13g2_decap_8 FILLER_44_1162 ();
 sg13g2_decap_4 FILLER_44_1169 ();
 sg13g2_fill_1 FILLER_44_1173 ();
 sg13g2_fill_1 FILLER_44_1203 ();
 sg13g2_decap_8 FILLER_44_1208 ();
 sg13g2_decap_4 FILLER_44_1215 ();
 sg13g2_fill_2 FILLER_44_1219 ();
 sg13g2_fill_2 FILLER_44_1269 ();
 sg13g2_fill_1 FILLER_44_1271 ();
 sg13g2_fill_1 FILLER_44_1304 ();
 sg13g2_fill_2 FILLER_44_1318 ();
 sg13g2_decap_8 FILLER_44_1332 ();
 sg13g2_fill_1 FILLER_44_1339 ();
 sg13g2_fill_1 FILLER_44_1354 ();
 sg13g2_fill_1 FILLER_44_1360 ();
 sg13g2_decap_4 FILLER_44_1370 ();
 sg13g2_fill_2 FILLER_44_1374 ();
 sg13g2_fill_2 FILLER_44_1381 ();
 sg13g2_fill_1 FILLER_44_1383 ();
 sg13g2_fill_1 FILLER_44_1395 ();
 sg13g2_fill_2 FILLER_44_1414 ();
 sg13g2_decap_4 FILLER_44_1429 ();
 sg13g2_decap_4 FILLER_44_1437 ();
 sg13g2_fill_1 FILLER_44_1441 ();
 sg13g2_fill_2 FILLER_44_1450 ();
 sg13g2_fill_2 FILLER_44_1456 ();
 sg13g2_fill_1 FILLER_44_1462 ();
 sg13g2_fill_1 FILLER_44_1468 ();
 sg13g2_fill_1 FILLER_44_1478 ();
 sg13g2_fill_2 FILLER_44_1499 ();
 sg13g2_fill_2 FILLER_44_1529 ();
 sg13g2_fill_1 FILLER_44_1546 ();
 sg13g2_decap_4 FILLER_44_1568 ();
 sg13g2_fill_2 FILLER_44_1572 ();
 sg13g2_decap_4 FILLER_44_1608 ();
 sg13g2_fill_1 FILLER_44_1612 ();
 sg13g2_fill_2 FILLER_44_1617 ();
 sg13g2_fill_1 FILLER_44_1619 ();
 sg13g2_fill_2 FILLER_44_1624 ();
 sg13g2_fill_1 FILLER_44_1626 ();
 sg13g2_fill_1 FILLER_44_1660 ();
 sg13g2_decap_8 FILLER_44_1680 ();
 sg13g2_decap_8 FILLER_44_1687 ();
 sg13g2_decap_4 FILLER_44_1694 ();
 sg13g2_fill_2 FILLER_44_1698 ();
 sg13g2_fill_2 FILLER_44_1710 ();
 sg13g2_fill_1 FILLER_44_1712 ();
 sg13g2_fill_1 FILLER_44_1755 ();
 sg13g2_fill_2 FILLER_44_1761 ();
 sg13g2_fill_1 FILLER_44_1763 ();
 sg13g2_decap_4 FILLER_44_1797 ();
 sg13g2_fill_2 FILLER_44_1806 ();
 sg13g2_decap_4 FILLER_44_1812 ();
 sg13g2_decap_8 FILLER_44_1830 ();
 sg13g2_decap_8 FILLER_44_1837 ();
 sg13g2_fill_1 FILLER_44_1844 ();
 sg13g2_decap_4 FILLER_44_1850 ();
 sg13g2_fill_1 FILLER_44_1854 ();
 sg13g2_decap_4 FILLER_44_1899 ();
 sg13g2_fill_2 FILLER_44_1903 ();
 sg13g2_fill_2 FILLER_44_1935 ();
 sg13g2_fill_1 FILLER_44_1937 ();
 sg13g2_decap_4 FILLER_44_1945 ();
 sg13g2_fill_1 FILLER_44_1949 ();
 sg13g2_fill_2 FILLER_44_1981 ();
 sg13g2_fill_1 FILLER_44_1994 ();
 sg13g2_decap_4 FILLER_44_2021 ();
 sg13g2_fill_2 FILLER_44_2025 ();
 sg13g2_fill_1 FILLER_44_2053 ();
 sg13g2_fill_2 FILLER_44_2080 ();
 sg13g2_fill_2 FILLER_44_2086 ();
 sg13g2_fill_2 FILLER_44_2113 ();
 sg13g2_fill_2 FILLER_44_2131 ();
 sg13g2_fill_1 FILLER_44_2133 ();
 sg13g2_decap_4 FILLER_44_2138 ();
 sg13g2_fill_2 FILLER_44_2142 ();
 sg13g2_fill_2 FILLER_44_2171 ();
 sg13g2_fill_1 FILLER_44_2183 ();
 sg13g2_fill_1 FILLER_44_2192 ();
 sg13g2_fill_2 FILLER_44_2222 ();
 sg13g2_fill_1 FILLER_44_2224 ();
 sg13g2_fill_1 FILLER_44_2231 ();
 sg13g2_fill_2 FILLER_44_2301 ();
 sg13g2_fill_1 FILLER_44_2303 ();
 sg13g2_fill_2 FILLER_44_2338 ();
 sg13g2_fill_1 FILLER_44_2432 ();
 sg13g2_fill_1 FILLER_44_2456 ();
 sg13g2_fill_1 FILLER_44_2468 ();
 sg13g2_fill_1 FILLER_44_2479 ();
 sg13g2_fill_2 FILLER_44_2495 ();
 sg13g2_fill_1 FILLER_44_2497 ();
 sg13g2_decap_8 FILLER_44_2503 ();
 sg13g2_fill_1 FILLER_44_2510 ();
 sg13g2_fill_2 FILLER_44_2551 ();
 sg13g2_decap_4 FILLER_44_2557 ();
 sg13g2_decap_8 FILLER_44_2590 ();
 sg13g2_decap_8 FILLER_44_2597 ();
 sg13g2_decap_8 FILLER_44_2610 ();
 sg13g2_decap_8 FILLER_44_2617 ();
 sg13g2_decap_8 FILLER_44_2624 ();
 sg13g2_decap_8 FILLER_44_2631 ();
 sg13g2_decap_8 FILLER_44_2638 ();
 sg13g2_decap_8 FILLER_44_2645 ();
 sg13g2_decap_8 FILLER_44_2652 ();
 sg13g2_decap_8 FILLER_44_2659 ();
 sg13g2_decap_4 FILLER_44_2666 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_4 ();
 sg13g2_fill_1 FILLER_45_20 ();
 sg13g2_fill_2 FILLER_45_25 ();
 sg13g2_fill_2 FILLER_45_37 ();
 sg13g2_decap_4 FILLER_45_43 ();
 sg13g2_fill_2 FILLER_45_55 ();
 sg13g2_decap_8 FILLER_45_96 ();
 sg13g2_decap_8 FILLER_45_108 ();
 sg13g2_fill_2 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_122 ();
 sg13g2_fill_1 FILLER_45_201 ();
 sg13g2_fill_2 FILLER_45_212 ();
 sg13g2_fill_1 FILLER_45_219 ();
 sg13g2_fill_1 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_234 ();
 sg13g2_fill_2 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_250 ();
 sg13g2_decap_4 FILLER_45_262 ();
 sg13g2_fill_2 FILLER_45_284 ();
 sg13g2_fill_1 FILLER_45_316 ();
 sg13g2_fill_1 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_fill_1 FILLER_45_357 ();
 sg13g2_fill_2 FILLER_45_361 ();
 sg13g2_decap_4 FILLER_45_399 ();
 sg13g2_fill_1 FILLER_45_412 ();
 sg13g2_decap_4 FILLER_45_443 ();
 sg13g2_fill_1 FILLER_45_447 ();
 sg13g2_fill_1 FILLER_45_457 ();
 sg13g2_decap_8 FILLER_45_471 ();
 sg13g2_decap_4 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_498 ();
 sg13g2_fill_1 FILLER_45_505 ();
 sg13g2_decap_4 FILLER_45_541 ();
 sg13g2_fill_1 FILLER_45_545 ();
 sg13g2_fill_1 FILLER_45_568 ();
 sg13g2_fill_2 FILLER_45_613 ();
 sg13g2_fill_1 FILLER_45_615 ();
 sg13g2_decap_8 FILLER_45_657 ();
 sg13g2_decap_8 FILLER_45_673 ();
 sg13g2_fill_1 FILLER_45_680 ();
 sg13g2_fill_2 FILLER_45_710 ();
 sg13g2_decap_4 FILLER_45_756 ();
 sg13g2_decap_4 FILLER_45_768 ();
 sg13g2_fill_1 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_fill_2 FILLER_45_795 ();
 sg13g2_fill_1 FILLER_45_797 ();
 sg13g2_fill_2 FILLER_45_803 ();
 sg13g2_fill_1 FILLER_45_805 ();
 sg13g2_decap_4 FILLER_45_840 ();
 sg13g2_fill_2 FILLER_45_854 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_fill_1 FILLER_45_862 ();
 sg13g2_fill_2 FILLER_45_966 ();
 sg13g2_fill_1 FILLER_45_979 ();
 sg13g2_fill_1 FILLER_45_984 ();
 sg13g2_fill_1 FILLER_45_990 ();
 sg13g2_fill_1 FILLER_45_995 ();
 sg13g2_decap_4 FILLER_45_1032 ();
 sg13g2_fill_1 FILLER_45_1036 ();
 sg13g2_fill_2 FILLER_45_1047 ();
 sg13g2_decap_8 FILLER_45_1075 ();
 sg13g2_decap_8 FILLER_45_1082 ();
 sg13g2_decap_8 FILLER_45_1089 ();
 sg13g2_decap_8 FILLER_45_1096 ();
 sg13g2_decap_4 FILLER_45_1103 ();
 sg13g2_decap_8 FILLER_45_1111 ();
 sg13g2_fill_2 FILLER_45_1118 ();
 sg13g2_decap_4 FILLER_45_1130 ();
 sg13g2_fill_2 FILLER_45_1134 ();
 sg13g2_decap_8 FILLER_45_1162 ();
 sg13g2_decap_4 FILLER_45_1169 ();
 sg13g2_fill_1 FILLER_45_1173 ();
 sg13g2_decap_8 FILLER_45_1184 ();
 sg13g2_decap_4 FILLER_45_1191 ();
 sg13g2_fill_1 FILLER_45_1195 ();
 sg13g2_decap_8 FILLER_45_1222 ();
 sg13g2_decap_4 FILLER_45_1229 ();
 sg13g2_fill_2 FILLER_45_1233 ();
 sg13g2_fill_2 FILLER_45_1240 ();
 sg13g2_fill_2 FILLER_45_1256 ();
 sg13g2_decap_4 FILLER_45_1269 ();
 sg13g2_fill_1 FILLER_45_1297 ();
 sg13g2_fill_1 FILLER_45_1303 ();
 sg13g2_fill_1 FILLER_45_1308 ();
 sg13g2_fill_1 FILLER_45_1314 ();
 sg13g2_fill_1 FILLER_45_1320 ();
 sg13g2_decap_4 FILLER_45_1336 ();
 sg13g2_fill_1 FILLER_45_1340 ();
 sg13g2_fill_1 FILLER_45_1353 ();
 sg13g2_decap_8 FILLER_45_1364 ();
 sg13g2_fill_1 FILLER_45_1371 ();
 sg13g2_decap_8 FILLER_45_1390 ();
 sg13g2_decap_8 FILLER_45_1397 ();
 sg13g2_decap_8 FILLER_45_1404 ();
 sg13g2_decap_4 FILLER_45_1411 ();
 sg13g2_fill_2 FILLER_45_1420 ();
 sg13g2_decap_8 FILLER_45_1429 ();
 sg13g2_decap_4 FILLER_45_1436 ();
 sg13g2_decap_8 FILLER_45_1444 ();
 sg13g2_decap_4 FILLER_45_1451 ();
 sg13g2_fill_1 FILLER_45_1455 ();
 sg13g2_fill_2 FILLER_45_1465 ();
 sg13g2_decap_8 FILLER_45_1471 ();
 sg13g2_decap_4 FILLER_45_1478 ();
 sg13g2_fill_1 FILLER_45_1482 ();
 sg13g2_fill_1 FILLER_45_1516 ();
 sg13g2_fill_1 FILLER_45_1521 ();
 sg13g2_decap_4 FILLER_45_1554 ();
 sg13g2_fill_2 FILLER_45_1558 ();
 sg13g2_fill_1 FILLER_45_1565 ();
 sg13g2_fill_2 FILLER_45_1570 ();
 sg13g2_decap_4 FILLER_45_1577 ();
 sg13g2_decap_8 FILLER_45_1585 ();
 sg13g2_fill_2 FILLER_45_1592 ();
 sg13g2_decap_8 FILLER_45_1604 ();
 sg13g2_fill_1 FILLER_45_1611 ();
 sg13g2_decap_8 FILLER_45_1617 ();
 sg13g2_decap_8 FILLER_45_1624 ();
 sg13g2_decap_8 FILLER_45_1631 ();
 sg13g2_decap_4 FILLER_45_1638 ();
 sg13g2_decap_8 FILLER_45_1647 ();
 sg13g2_decap_8 FILLER_45_1689 ();
 sg13g2_decap_8 FILLER_45_1699 ();
 sg13g2_decap_8 FILLER_45_1706 ();
 sg13g2_fill_1 FILLER_45_1718 ();
 sg13g2_decap_8 FILLER_45_1726 ();
 sg13g2_fill_2 FILLER_45_1766 ();
 sg13g2_fill_1 FILLER_45_1778 ();
 sg13g2_fill_2 FILLER_45_1788 ();
 sg13g2_fill_1 FILLER_45_1799 ();
 sg13g2_fill_2 FILLER_45_1808 ();
 sg13g2_fill_1 FILLER_45_1810 ();
 sg13g2_fill_1 FILLER_45_1828 ();
 sg13g2_fill_2 FILLER_45_1854 ();
 sg13g2_fill_1 FILLER_45_1856 ();
 sg13g2_decap_8 FILLER_45_1883 ();
 sg13g2_fill_1 FILLER_45_1890 ();
 sg13g2_decap_8 FILLER_45_1896 ();
 sg13g2_decap_8 FILLER_45_1903 ();
 sg13g2_decap_8 FILLER_45_1920 ();
 sg13g2_decap_4 FILLER_45_1927 ();
 sg13g2_decap_8 FILLER_45_1946 ();
 sg13g2_decap_4 FILLER_45_1953 ();
 sg13g2_fill_1 FILLER_45_1957 ();
 sg13g2_fill_1 FILLER_45_1962 ();
 sg13g2_fill_2 FILLER_45_1973 ();
 sg13g2_fill_1 FILLER_45_1975 ();
 sg13g2_decap_8 FILLER_45_2003 ();
 sg13g2_decap_8 FILLER_45_2010 ();
 sg13g2_fill_2 FILLER_45_2017 ();
 sg13g2_fill_1 FILLER_45_2019 ();
 sg13g2_fill_2 FILLER_45_2056 ();
 sg13g2_fill_1 FILLER_45_2114 ();
 sg13g2_fill_1 FILLER_45_2127 ();
 sg13g2_decap_4 FILLER_45_2138 ();
 sg13g2_fill_2 FILLER_45_2142 ();
 sg13g2_decap_8 FILLER_45_2169 ();
 sg13g2_decap_8 FILLER_45_2176 ();
 sg13g2_decap_8 FILLER_45_2183 ();
 sg13g2_fill_1 FILLER_45_2194 ();
 sg13g2_fill_1 FILLER_45_2205 ();
 sg13g2_decap_4 FILLER_45_2209 ();
 sg13g2_fill_1 FILLER_45_2261 ();
 sg13g2_fill_2 FILLER_45_2289 ();
 sg13g2_decap_8 FILLER_45_2311 ();
 sg13g2_decap_8 FILLER_45_2318 ();
 sg13g2_decap_4 FILLER_45_2325 ();
 sg13g2_fill_1 FILLER_45_2329 ();
 sg13g2_fill_2 FILLER_45_2334 ();
 sg13g2_fill_1 FILLER_45_2336 ();
 sg13g2_fill_1 FILLER_45_2400 ();
 sg13g2_fill_2 FILLER_45_2424 ();
 sg13g2_fill_1 FILLER_45_2431 ();
 sg13g2_fill_1 FILLER_45_2436 ();
 sg13g2_fill_1 FILLER_45_2471 ();
 sg13g2_fill_2 FILLER_45_2502 ();
 sg13g2_fill_1 FILLER_45_2504 ();
 sg13g2_fill_2 FILLER_45_2535 ();
 sg13g2_decap_8 FILLER_45_2541 ();
 sg13g2_fill_1 FILLER_45_2548 ();
 sg13g2_fill_2 FILLER_45_2589 ();
 sg13g2_fill_1 FILLER_45_2591 ();
 sg13g2_decap_8 FILLER_45_2596 ();
 sg13g2_decap_4 FILLER_45_2624 ();
 sg13g2_fill_1 FILLER_45_2628 ();
 sg13g2_decap_8 FILLER_45_2655 ();
 sg13g2_decap_8 FILLER_45_2662 ();
 sg13g2_fill_1 FILLER_45_2669 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_11 ();
 sg13g2_decap_8 FILLER_46_38 ();
 sg13g2_decap_8 FILLER_46_45 ();
 sg13g2_decap_8 FILLER_46_52 ();
 sg13g2_decap_8 FILLER_46_59 ();
 sg13g2_fill_2 FILLER_46_66 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_decap_4 FILLER_46_102 ();
 sg13g2_decap_8 FILLER_46_110 ();
 sg13g2_decap_4 FILLER_46_117 ();
 sg13g2_fill_2 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_170 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_decap_4 FILLER_46_202 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_fill_1 FILLER_46_219 ();
 sg13g2_decap_4 FILLER_46_261 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_fill_2 FILLER_46_275 ();
 sg13g2_decap_8 FILLER_46_345 ();
 sg13g2_fill_2 FILLER_46_352 ();
 sg13g2_fill_1 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_fill_2 FILLER_46_402 ();
 sg13g2_fill_1 FILLER_46_410 ();
 sg13g2_fill_2 FILLER_46_416 ();
 sg13g2_fill_1 FILLER_46_422 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_fill_1 FILLER_46_437 ();
 sg13g2_decap_4 FILLER_46_458 ();
 sg13g2_fill_2 FILLER_46_462 ();
 sg13g2_fill_1 FILLER_46_509 ();
 sg13g2_fill_1 FILLER_46_520 ();
 sg13g2_fill_2 FILLER_46_531 ();
 sg13g2_fill_1 FILLER_46_537 ();
 sg13g2_fill_1 FILLER_46_579 ();
 sg13g2_fill_2 FILLER_46_640 ();
 sg13g2_decap_8 FILLER_46_671 ();
 sg13g2_fill_1 FILLER_46_678 ();
 sg13g2_fill_1 FILLER_46_736 ();
 sg13g2_decap_4 FILLER_46_771 ();
 sg13g2_fill_1 FILLER_46_775 ();
 sg13g2_decap_8 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_4 FILLER_46_799 ();
 sg13g2_fill_2 FILLER_46_803 ();
 sg13g2_decap_4 FILLER_46_827 ();
 sg13g2_fill_2 FILLER_46_867 ();
 sg13g2_decap_4 FILLER_46_875 ();
 sg13g2_fill_2 FILLER_46_879 ();
 sg13g2_decap_4 FILLER_46_885 ();
 sg13g2_fill_2 FILLER_46_889 ();
 sg13g2_fill_2 FILLER_46_909 ();
 sg13g2_fill_1 FILLER_46_917 ();
 sg13g2_fill_2 FILLER_46_960 ();
 sg13g2_fill_1 FILLER_46_967 ();
 sg13g2_fill_1 FILLER_46_1011 ();
 sg13g2_fill_1 FILLER_46_1022 ();
 sg13g2_fill_1 FILLER_46_1049 ();
 sg13g2_fill_1 FILLER_46_1076 ();
 sg13g2_decap_8 FILLER_46_1081 ();
 sg13g2_fill_2 FILLER_46_1088 ();
 sg13g2_fill_1 FILLER_46_1134 ();
 sg13g2_fill_2 FILLER_46_1161 ();
 sg13g2_fill_2 FILLER_46_1189 ();
 sg13g2_decap_4 FILLER_46_1217 ();
 sg13g2_decap_8 FILLER_46_1231 ();
 sg13g2_fill_1 FILLER_46_1238 ();
 sg13g2_decap_8 FILLER_46_1247 ();
 sg13g2_fill_1 FILLER_46_1254 ();
 sg13g2_decap_4 FILLER_46_1270 ();
 sg13g2_fill_1 FILLER_46_1274 ();
 sg13g2_fill_2 FILLER_46_1280 ();
 sg13g2_decap_8 FILLER_46_1286 ();
 sg13g2_decap_8 FILLER_46_1293 ();
 sg13g2_fill_2 FILLER_46_1300 ();
 sg13g2_fill_1 FILLER_46_1307 ();
 sg13g2_decap_4 FILLER_46_1323 ();
 sg13g2_fill_2 FILLER_46_1327 ();
 sg13g2_decap_4 FILLER_46_1335 ();
 sg13g2_fill_1 FILLER_46_1345 ();
 sg13g2_decap_8 FILLER_46_1355 ();
 sg13g2_fill_2 FILLER_46_1362 ();
 sg13g2_fill_1 FILLER_46_1391 ();
 sg13g2_decap_8 FILLER_46_1397 ();
 sg13g2_decap_8 FILLER_46_1404 ();
 sg13g2_fill_2 FILLER_46_1411 ();
 sg13g2_fill_1 FILLER_46_1413 ();
 sg13g2_fill_1 FILLER_46_1450 ();
 sg13g2_decap_4 FILLER_46_1487 ();
 sg13g2_fill_2 FILLER_46_1524 ();
 sg13g2_fill_1 FILLER_46_1529 ();
 sg13g2_fill_2 FILLER_46_1535 ();
 sg13g2_fill_2 FILLER_46_1551 ();
 sg13g2_fill_1 FILLER_46_1553 ();
 sg13g2_decap_8 FILLER_46_1563 ();
 sg13g2_fill_2 FILLER_46_1570 ();
 sg13g2_fill_1 FILLER_46_1572 ();
 sg13g2_decap_8 FILLER_46_1578 ();
 sg13g2_fill_1 FILLER_46_1589 ();
 sg13g2_fill_2 FILLER_46_1620 ();
 sg13g2_fill_1 FILLER_46_1622 ();
 sg13g2_fill_1 FILLER_46_1637 ();
 sg13g2_fill_1 FILLER_46_1646 ();
 sg13g2_fill_1 FILLER_46_1652 ();
 sg13g2_fill_2 FILLER_46_1658 ();
 sg13g2_fill_2 FILLER_46_1668 ();
 sg13g2_fill_1 FILLER_46_1685 ();
 sg13g2_fill_2 FILLER_46_1690 ();
 sg13g2_decap_4 FILLER_46_1717 ();
 sg13g2_fill_2 FILLER_46_1726 ();
 sg13g2_fill_2 FILLER_46_1738 ();
 sg13g2_fill_1 FILLER_46_1748 ();
 sg13g2_fill_2 FILLER_46_1752 ();
 sg13g2_fill_2 FILLER_46_1798 ();
 sg13g2_fill_1 FILLER_46_1800 ();
 sg13g2_fill_1 FILLER_46_1821 ();
 sg13g2_fill_2 FILLER_46_1826 ();
 sg13g2_fill_1 FILLER_46_1833 ();
 sg13g2_decap_8 FILLER_46_1843 ();
 sg13g2_fill_1 FILLER_46_1850 ();
 sg13g2_decap_8 FILLER_46_1856 ();
 sg13g2_fill_2 FILLER_46_1863 ();
 sg13g2_decap_4 FILLER_46_1873 ();
 sg13g2_fill_1 FILLER_46_1903 ();
 sg13g2_fill_1 FILLER_46_1930 ();
 sg13g2_fill_1 FILLER_46_1961 ();
 sg13g2_decap_8 FILLER_46_1974 ();
 sg13g2_fill_2 FILLER_46_1981 ();
 sg13g2_decap_4 FILLER_46_2009 ();
 sg13g2_fill_2 FILLER_46_2013 ();
 sg13g2_decap_4 FILLER_46_2019 ();
 sg13g2_decap_8 FILLER_46_2037 ();
 sg13g2_fill_2 FILLER_46_2044 ();
 sg13g2_fill_1 FILLER_46_2046 ();
 sg13g2_decap_8 FILLER_46_2154 ();
 sg13g2_fill_1 FILLER_46_2161 ();
 sg13g2_decap_4 FILLER_46_2192 ();
 sg13g2_decap_4 FILLER_46_2216 ();
 sg13g2_fill_2 FILLER_46_2220 ();
 sg13g2_fill_2 FILLER_46_2229 ();
 sg13g2_fill_2 FILLER_46_2234 ();
 sg13g2_fill_1 FILLER_46_2278 ();
 sg13g2_fill_2 FILLER_46_2305 ();
 sg13g2_fill_1 FILLER_46_2307 ();
 sg13g2_decap_4 FILLER_46_2312 ();
 sg13g2_decap_4 FILLER_46_2330 ();
 sg13g2_fill_1 FILLER_46_2334 ();
 sg13g2_fill_2 FILLER_46_2340 ();
 sg13g2_fill_1 FILLER_46_2342 ();
 sg13g2_decap_4 FILLER_46_2350 ();
 sg13g2_fill_1 FILLER_46_2373 ();
 sg13g2_fill_1 FILLER_46_2378 ();
 sg13g2_fill_1 FILLER_46_2391 ();
 sg13g2_fill_1 FILLER_46_2412 ();
 sg13g2_fill_1 FILLER_46_2434 ();
 sg13g2_decap_8 FILLER_46_2500 ();
 sg13g2_fill_1 FILLER_46_2507 ();
 sg13g2_fill_2 FILLER_46_2546 ();
 sg13g2_fill_1 FILLER_46_2548 ();
 sg13g2_decap_8 FILLER_46_2553 ();
 sg13g2_fill_1 FILLER_46_2603 ();
 sg13g2_fill_2 FILLER_46_2633 ();
 sg13g2_fill_1 FILLER_46_2635 ();
 sg13g2_decap_8 FILLER_46_2640 ();
 sg13g2_decap_8 FILLER_46_2647 ();
 sg13g2_decap_8 FILLER_46_2654 ();
 sg13g2_decap_8 FILLER_46_2661 ();
 sg13g2_fill_2 FILLER_46_2668 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_26 ();
 sg13g2_decap_8 FILLER_47_33 ();
 sg13g2_decap_8 FILLER_47_40 ();
 sg13g2_decap_8 FILLER_47_47 ();
 sg13g2_decap_8 FILLER_47_54 ();
 sg13g2_decap_8 FILLER_47_61 ();
 sg13g2_decap_4 FILLER_47_68 ();
 sg13g2_fill_2 FILLER_47_72 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_1 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_fill_1 FILLER_47_156 ();
 sg13g2_decap_4 FILLER_47_177 ();
 sg13g2_fill_2 FILLER_47_181 ();
 sg13g2_decap_4 FILLER_47_196 ();
 sg13g2_fill_1 FILLER_47_205 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_decap_8 FILLER_47_235 ();
 sg13g2_fill_1 FILLER_47_242 ();
 sg13g2_fill_2 FILLER_47_252 ();
 sg13g2_fill_1 FILLER_47_254 ();
 sg13g2_fill_2 FILLER_47_260 ();
 sg13g2_fill_2 FILLER_47_271 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_326 ();
 sg13g2_fill_2 FILLER_47_333 ();
 sg13g2_fill_2 FILLER_47_339 ();
 sg13g2_fill_1 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_347 ();
 sg13g2_fill_1 FILLER_47_362 ();
 sg13g2_fill_2 FILLER_47_368 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_47_379 ();
 sg13g2_fill_1 FILLER_47_383 ();
 sg13g2_decap_4 FILLER_47_399 ();
 sg13g2_decap_4 FILLER_47_412 ();
 sg13g2_fill_1 FILLER_47_416 ();
 sg13g2_fill_2 FILLER_47_470 ();
 sg13g2_fill_1 FILLER_47_472 ();
 sg13g2_fill_2 FILLER_47_516 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_fill_2 FILLER_47_577 ();
 sg13g2_fill_1 FILLER_47_591 ();
 sg13g2_fill_2 FILLER_47_599 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_fill_1 FILLER_47_722 ();
 sg13g2_fill_1 FILLER_47_769 ();
 sg13g2_fill_2 FILLER_47_774 ();
 sg13g2_fill_1 FILLER_47_836 ();
 sg13g2_fill_1 FILLER_47_845 ();
 sg13g2_fill_1 FILLER_47_890 ();
 sg13g2_fill_2 FILLER_47_921 ();
 sg13g2_fill_1 FILLER_47_965 ();
 sg13g2_fill_1 FILLER_47_987 ();
 sg13g2_fill_2 FILLER_47_1011 ();
 sg13g2_fill_2 FILLER_47_1021 ();
 sg13g2_fill_1 FILLER_47_1023 ();
 sg13g2_fill_1 FILLER_47_1030 ();
 sg13g2_decap_8 FILLER_47_1077 ();
 sg13g2_fill_1 FILLER_47_1084 ();
 sg13g2_fill_2 FILLER_47_1094 ();
 sg13g2_decap_4 FILLER_47_1122 ();
 sg13g2_fill_1 FILLER_47_1126 ();
 sg13g2_fill_2 FILLER_47_1137 ();
 sg13g2_fill_2 FILLER_47_1176 ();
 sg13g2_fill_2 FILLER_47_1181 ();
 sg13g2_fill_1 FILLER_47_1183 ();
 sg13g2_fill_2 FILLER_47_1214 ();
 sg13g2_decap_8 FILLER_47_1253 ();
 sg13g2_decap_8 FILLER_47_1260 ();
 sg13g2_decap_4 FILLER_47_1283 ();
 sg13g2_fill_2 FILLER_47_1287 ();
 sg13g2_fill_1 FILLER_47_1312 ();
 sg13g2_fill_2 FILLER_47_1317 ();
 sg13g2_decap_8 FILLER_47_1333 ();
 sg13g2_decap_4 FILLER_47_1340 ();
 sg13g2_fill_2 FILLER_47_1344 ();
 sg13g2_fill_2 FILLER_47_1367 ();
 sg13g2_fill_2 FILLER_47_1413 ();
 sg13g2_fill_2 FILLER_47_1420 ();
 sg13g2_fill_1 FILLER_47_1429 ();
 sg13g2_fill_1 FILLER_47_1456 ();
 sg13g2_decap_4 FILLER_47_1483 ();
 sg13g2_fill_2 FILLER_47_1548 ();
 sg13g2_fill_2 FILLER_47_1562 ();
 sg13g2_decap_8 FILLER_47_1569 ();
 sg13g2_fill_1 FILLER_47_1576 ();
 sg13g2_fill_2 FILLER_47_1585 ();
 sg13g2_fill_2 FILLER_47_1619 ();
 sg13g2_fill_1 FILLER_47_1621 ();
 sg13g2_fill_1 FILLER_47_1631 ();
 sg13g2_fill_1 FILLER_47_1646 ();
 sg13g2_fill_1 FILLER_47_1651 ();
 sg13g2_fill_2 FILLER_47_1657 ();
 sg13g2_fill_1 FILLER_47_1659 ();
 sg13g2_fill_1 FILLER_47_1665 ();
 sg13g2_fill_2 FILLER_47_1671 ();
 sg13g2_fill_1 FILLER_47_1673 ();
 sg13g2_fill_1 FILLER_47_1696 ();
 sg13g2_decap_4 FILLER_47_1716 ();
 sg13g2_decap_8 FILLER_47_1724 ();
 sg13g2_fill_2 FILLER_47_1731 ();
 sg13g2_fill_1 FILLER_47_1733 ();
 sg13g2_fill_1 FILLER_47_1744 ();
 sg13g2_fill_2 FILLER_47_1754 ();
 sg13g2_fill_2 FILLER_47_1761 ();
 sg13g2_fill_2 FILLER_47_1806 ();
 sg13g2_decap_4 FILLER_47_1818 ();
 sg13g2_fill_2 FILLER_47_1827 ();
 sg13g2_fill_2 FILLER_47_1843 ();
 sg13g2_fill_1 FILLER_47_1845 ();
 sg13g2_decap_8 FILLER_47_1850 ();
 sg13g2_decap_8 FILLER_47_1868 ();
 sg13g2_fill_1 FILLER_47_1875 ();
 sg13g2_decap_8 FILLER_47_1887 ();
 sg13g2_decap_8 FILLER_47_1894 ();
 sg13g2_decap_4 FILLER_47_1901 ();
 sg13g2_fill_1 FILLER_47_1949 ();
 sg13g2_fill_1 FILLER_47_2002 ();
 sg13g2_fill_2 FILLER_47_2039 ();
 sg13g2_fill_1 FILLER_47_2041 ();
 sg13g2_fill_2 FILLER_47_2090 ();
 sg13g2_fill_1 FILLER_47_2096 ();
 sg13g2_decap_8 FILLER_47_2166 ();
 sg13g2_fill_1 FILLER_47_2173 ();
 sg13g2_fill_2 FILLER_47_2178 ();
 sg13g2_fill_1 FILLER_47_2245 ();
 sg13g2_fill_1 FILLER_47_2315 ();
 sg13g2_fill_1 FILLER_47_2320 ();
 sg13g2_fill_2 FILLER_47_2326 ();
 sg13g2_decap_4 FILLER_47_2367 ();
 sg13g2_fill_1 FILLER_47_2371 ();
 sg13g2_fill_2 FILLER_47_2379 ();
 sg13g2_fill_2 FILLER_47_2413 ();
 sg13g2_fill_2 FILLER_47_2441 ();
 sg13g2_fill_2 FILLER_47_2478 ();
 sg13g2_fill_1 FILLER_47_2499 ();
 sg13g2_decap_8 FILLER_47_2505 ();
 sg13g2_decap_8 FILLER_47_2512 ();
 sg13g2_fill_1 FILLER_47_2532 ();
 sg13g2_decap_8 FILLER_47_2537 ();
 sg13g2_decap_8 FILLER_47_2544 ();
 sg13g2_decap_8 FILLER_47_2551 ();
 sg13g2_decap_4 FILLER_47_2558 ();
 sg13g2_fill_2 FILLER_47_2562 ();
 sg13g2_decap_4 FILLER_47_2576 ();
 sg13g2_decap_8 FILLER_47_2632 ();
 sg13g2_decap_8 FILLER_47_2639 ();
 sg13g2_decap_8 FILLER_47_2646 ();
 sg13g2_decap_8 FILLER_47_2653 ();
 sg13g2_decap_8 FILLER_47_2660 ();
 sg13g2_fill_2 FILLER_47_2667 ();
 sg13g2_fill_1 FILLER_47_2669 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_28 ();
 sg13g2_fill_1 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_50 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_decap_8 FILLER_48_104 ();
 sg13g2_fill_2 FILLER_48_111 ();
 sg13g2_fill_1 FILLER_48_113 ();
 sg13g2_decap_8 FILLER_48_118 ();
 sg13g2_decap_4 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_139 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_168 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_178 ();
 sg13g2_fill_2 FILLER_48_197 ();
 sg13g2_decap_4 FILLER_48_249 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_323 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_fill_2 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_367 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_2 FILLER_48_418 ();
 sg13g2_fill_2 FILLER_48_426 ();
 sg13g2_fill_1 FILLER_48_428 ();
 sg13g2_decap_8 FILLER_48_459 ();
 sg13g2_decap_8 FILLER_48_466 ();
 sg13g2_decap_4 FILLER_48_482 ();
 sg13g2_fill_2 FILLER_48_530 ();
 sg13g2_fill_1 FILLER_48_549 ();
 sg13g2_fill_1 FILLER_48_554 ();
 sg13g2_fill_2 FILLER_48_582 ();
 sg13g2_fill_2 FILLER_48_588 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_fill_2 FILLER_48_623 ();
 sg13g2_fill_2 FILLER_48_635 ();
 sg13g2_fill_1 FILLER_48_653 ();
 sg13g2_decap_8 FILLER_48_678 ();
 sg13g2_fill_2 FILLER_48_685 ();
 sg13g2_fill_1 FILLER_48_692 ();
 sg13g2_fill_1 FILLER_48_697 ();
 sg13g2_fill_1 FILLER_48_721 ();
 sg13g2_fill_2 FILLER_48_726 ();
 sg13g2_fill_2 FILLER_48_763 ();
 sg13g2_fill_1 FILLER_48_765 ();
 sg13g2_decap_4 FILLER_48_770 ();
 sg13g2_fill_1 FILLER_48_778 ();
 sg13g2_fill_2 FILLER_48_783 ();
 sg13g2_fill_1 FILLER_48_789 ();
 sg13g2_fill_2 FILLER_48_816 ();
 sg13g2_fill_2 FILLER_48_853 ();
 sg13g2_decap_4 FILLER_48_863 ();
 sg13g2_decap_4 FILLER_48_885 ();
 sg13g2_fill_2 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_894 ();
 sg13g2_fill_1 FILLER_48_905 ();
 sg13g2_fill_2 FILLER_48_924 ();
 sg13g2_fill_2 FILLER_48_992 ();
 sg13g2_fill_1 FILLER_48_1042 ();
 sg13g2_fill_2 FILLER_48_1061 ();
 sg13g2_fill_2 FILLER_48_1082 ();
 sg13g2_decap_8 FILLER_48_1144 ();
 sg13g2_decap_8 FILLER_48_1151 ();
 sg13g2_decap_8 FILLER_48_1158 ();
 sg13g2_decap_8 FILLER_48_1165 ();
 sg13g2_fill_2 FILLER_48_1172 ();
 sg13g2_fill_2 FILLER_48_1188 ();
 sg13g2_fill_2 FILLER_48_1203 ();
 sg13g2_decap_4 FILLER_48_1232 ();
 sg13g2_fill_1 FILLER_48_1236 ();
 sg13g2_fill_2 FILLER_48_1246 ();
 sg13g2_decap_8 FILLER_48_1253 ();
 sg13g2_fill_2 FILLER_48_1264 ();
 sg13g2_decap_8 FILLER_48_1271 ();
 sg13g2_fill_2 FILLER_48_1278 ();
 sg13g2_fill_2 FILLER_48_1296 ();
 sg13g2_decap_8 FILLER_48_1321 ();
 sg13g2_decap_4 FILLER_48_1328 ();
 sg13g2_fill_2 FILLER_48_1332 ();
 sg13g2_decap_4 FILLER_48_1338 ();
 sg13g2_fill_2 FILLER_48_1372 ();
 sg13g2_fill_1 FILLER_48_1378 ();
 sg13g2_fill_1 FILLER_48_1385 ();
 sg13g2_fill_1 FILLER_48_1391 ();
 sg13g2_fill_2 FILLER_48_1403 ();
 sg13g2_fill_1 FILLER_48_1405 ();
 sg13g2_fill_2 FILLER_48_1419 ();
 sg13g2_fill_1 FILLER_48_1421 ();
 sg13g2_fill_2 FILLER_48_1431 ();
 sg13g2_fill_1 FILLER_48_1433 ();
 sg13g2_decap_4 FILLER_48_1443 ();
 sg13g2_decap_4 FILLER_48_1465 ();
 sg13g2_fill_1 FILLER_48_1482 ();
 sg13g2_fill_2 FILLER_48_1498 ();
 sg13g2_fill_2 FILLER_48_1514 ();
 sg13g2_fill_1 FILLER_48_1520 ();
 sg13g2_fill_1 FILLER_48_1524 ();
 sg13g2_decap_4 FILLER_48_1543 ();
 sg13g2_decap_4 FILLER_48_1577 ();
 sg13g2_fill_2 FILLER_48_1585 ();
 sg13g2_fill_1 FILLER_48_1587 ();
 sg13g2_decap_4 FILLER_48_1593 ();
 sg13g2_fill_1 FILLER_48_1597 ();
 sg13g2_decap_8 FILLER_48_1602 ();
 sg13g2_fill_1 FILLER_48_1619 ();
 sg13g2_decap_8 FILLER_48_1624 ();
 sg13g2_decap_4 FILLER_48_1631 ();
 sg13g2_fill_1 FILLER_48_1639 ();
 sg13g2_fill_1 FILLER_48_1644 ();
 sg13g2_decap_4 FILLER_48_1657 ();
 sg13g2_fill_1 FILLER_48_1710 ();
 sg13g2_decap_4 FILLER_48_1739 ();
 sg13g2_fill_1 FILLER_48_1743 ();
 sg13g2_fill_2 FILLER_48_1749 ();
 sg13g2_fill_2 FILLER_48_1756 ();
 sg13g2_fill_1 FILLER_48_1758 ();
 sg13g2_fill_2 FILLER_48_1764 ();
 sg13g2_fill_1 FILLER_48_1774 ();
 sg13g2_fill_1 FILLER_48_1785 ();
 sg13g2_fill_1 FILLER_48_1800 ();
 sg13g2_decap_4 FILLER_48_1805 ();
 sg13g2_fill_2 FILLER_48_1813 ();
 sg13g2_fill_2 FILLER_48_1820 ();
 sg13g2_fill_1 FILLER_48_1822 ();
 sg13g2_fill_2 FILLER_48_1837 ();
 sg13g2_decap_8 FILLER_48_1847 ();
 sg13g2_decap_8 FILLER_48_1854 ();
 sg13g2_decap_8 FILLER_48_1861 ();
 sg13g2_decap_8 FILLER_48_1868 ();
 sg13g2_decap_8 FILLER_48_1875 ();
 sg13g2_fill_2 FILLER_48_1882 ();
 sg13g2_decap_8 FILLER_48_1888 ();
 sg13g2_decap_8 FILLER_48_1895 ();
 sg13g2_decap_8 FILLER_48_1902 ();
 sg13g2_fill_2 FILLER_48_1909 ();
 sg13g2_fill_1 FILLER_48_1911 ();
 sg13g2_decap_8 FILLER_48_1916 ();
 sg13g2_decap_8 FILLER_48_1923 ();
 sg13g2_fill_2 FILLER_48_2054 ();
 sg13g2_fill_1 FILLER_48_2126 ();
 sg13g2_fill_1 FILLER_48_2139 ();
 sg13g2_fill_1 FILLER_48_2144 ();
 sg13g2_fill_1 FILLER_48_2155 ();
 sg13g2_fill_1 FILLER_48_2182 ();
 sg13g2_decap_8 FILLER_48_2213 ();
 sg13g2_fill_2 FILLER_48_2220 ();
 sg13g2_fill_1 FILLER_48_2222 ();
 sg13g2_decap_8 FILLER_48_2244 ();
 sg13g2_fill_2 FILLER_48_2291 ();
 sg13g2_fill_1 FILLER_48_2363 ();
 sg13g2_fill_1 FILLER_48_2377 ();
 sg13g2_decap_8 FILLER_48_2450 ();
 sg13g2_decap_8 FILLER_48_2457 ();
 sg13g2_fill_1 FILLER_48_2464 ();
 sg13g2_fill_1 FILLER_48_2499 ();
 sg13g2_fill_1 FILLER_48_2531 ();
 sg13g2_decap_8 FILLER_48_2550 ();
 sg13g2_decap_8 FILLER_48_2557 ();
 sg13g2_decap_4 FILLER_48_2564 ();
 sg13g2_fill_1 FILLER_48_2568 ();
 sg13g2_decap_8 FILLER_48_2574 ();
 sg13g2_decap_8 FILLER_48_2581 ();
 sg13g2_decap_8 FILLER_48_2588 ();
 sg13g2_fill_2 FILLER_48_2595 ();
 sg13g2_fill_1 FILLER_48_2597 ();
 sg13g2_decap_8 FILLER_48_2627 ();
 sg13g2_decap_8 FILLER_48_2634 ();
 sg13g2_decap_8 FILLER_48_2641 ();
 sg13g2_decap_8 FILLER_48_2648 ();
 sg13g2_decap_8 FILLER_48_2655 ();
 sg13g2_decap_8 FILLER_48_2662 ();
 sg13g2_fill_1 FILLER_48_2669 ();
 sg13g2_fill_2 FILLER_49_4 ();
 sg13g2_fill_1 FILLER_49_6 ();
 sg13g2_decap_4 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_131 ();
 sg13g2_fill_2 FILLER_49_142 ();
 sg13g2_fill_1 FILLER_49_144 ();
 sg13g2_fill_2 FILLER_49_154 ();
 sg13g2_fill_1 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_160 ();
 sg13g2_fill_2 FILLER_49_176 ();
 sg13g2_fill_1 FILLER_49_178 ();
 sg13g2_fill_2 FILLER_49_224 ();
 sg13g2_fill_1 FILLER_49_226 ();
 sg13g2_fill_1 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_fill_1 FILLER_49_254 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_4 FILLER_49_271 ();
 sg13g2_fill_1 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_328 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_fill_1 FILLER_49_398 ();
 sg13g2_fill_2 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_412 ();
 sg13g2_decap_4 FILLER_49_418 ();
 sg13g2_decap_4 FILLER_49_430 ();
 sg13g2_fill_2 FILLER_49_447 ();
 sg13g2_fill_1 FILLER_49_449 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_463 ();
 sg13g2_fill_1 FILLER_49_478 ();
 sg13g2_fill_1 FILLER_49_531 ();
 sg13g2_fill_1 FILLER_49_537 ();
 sg13g2_fill_2 FILLER_49_543 ();
 sg13g2_fill_1 FILLER_49_558 ();
 sg13g2_fill_1 FILLER_49_603 ();
 sg13g2_fill_2 FILLER_49_630 ();
 sg13g2_fill_2 FILLER_49_635 ();
 sg13g2_fill_1 FILLER_49_649 ();
 sg13g2_fill_2 FILLER_49_654 ();
 sg13g2_fill_2 FILLER_49_661 ();
 sg13g2_decap_4 FILLER_49_670 ();
 sg13g2_fill_2 FILLER_49_674 ();
 sg13g2_decap_8 FILLER_49_702 ();
 sg13g2_fill_2 FILLER_49_733 ();
 sg13g2_fill_2 FILLER_49_746 ();
 sg13g2_decap_4 FILLER_49_755 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_4 FILLER_49_770 ();
 sg13g2_fill_1 FILLER_49_774 ();
 sg13g2_fill_2 FILLER_49_780 ();
 sg13g2_fill_2 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_966 ();
 sg13g2_fill_2 FILLER_49_997 ();
 sg13g2_fill_1 FILLER_49_1004 ();
 sg13g2_fill_1 FILLER_49_1014 ();
 sg13g2_fill_1 FILLER_49_1056 ();
 sg13g2_decap_8 FILLER_49_1061 ();
 sg13g2_decap_8 FILLER_49_1068 ();
 sg13g2_decap_4 FILLER_49_1075 ();
 sg13g2_fill_1 FILLER_49_1084 ();
 sg13g2_fill_1 FILLER_49_1114 ();
 sg13g2_decap_8 FILLER_49_1141 ();
 sg13g2_decap_8 FILLER_49_1174 ();
 sg13g2_fill_1 FILLER_49_1181 ();
 sg13g2_fill_1 FILLER_49_1204 ();
 sg13g2_fill_1 FILLER_49_1210 ();
 sg13g2_decap_8 FILLER_49_1255 ();
 sg13g2_fill_2 FILLER_49_1262 ();
 sg13g2_fill_2 FILLER_49_1279 ();
 sg13g2_fill_1 FILLER_49_1281 ();
 sg13g2_decap_4 FILLER_49_1297 ();
 sg13g2_decap_4 FILLER_49_1308 ();
 sg13g2_fill_2 FILLER_49_1312 ();
 sg13g2_decap_8 FILLER_49_1319 ();
 sg13g2_fill_1 FILLER_49_1330 ();
 sg13g2_fill_2 FILLER_49_1340 ();
 sg13g2_fill_1 FILLER_49_1342 ();
 sg13g2_fill_1 FILLER_49_1349 ();
 sg13g2_fill_1 FILLER_49_1371 ();
 sg13g2_fill_1 FILLER_49_1382 ();
 sg13g2_fill_1 FILLER_49_1389 ();
 sg13g2_fill_1 FILLER_49_1401 ();
 sg13g2_fill_1 FILLER_49_1428 ();
 sg13g2_decap_4 FILLER_49_1434 ();
 sg13g2_fill_1 FILLER_49_1438 ();
 sg13g2_decap_4 FILLER_49_1500 ();
 sg13g2_decap_8 FILLER_49_1517 ();
 sg13g2_fill_2 FILLER_49_1535 ();
 sg13g2_decap_8 FILLER_49_1542 ();
 sg13g2_fill_1 FILLER_49_1549 ();
 sg13g2_decap_4 FILLER_49_1583 ();
 sg13g2_decap_4 FILLER_49_1591 ();
 sg13g2_fill_2 FILLER_49_1595 ();
 sg13g2_fill_2 FILLER_49_1602 ();
 sg13g2_fill_1 FILLER_49_1604 ();
 sg13g2_fill_1 FILLER_49_1655 ();
 sg13g2_fill_2 FILLER_49_1661 ();
 sg13g2_fill_2 FILLER_49_1667 ();
 sg13g2_fill_1 FILLER_49_1669 ();
 sg13g2_fill_1 FILLER_49_1689 ();
 sg13g2_fill_2 FILLER_49_1731 ();
 sg13g2_fill_2 FILLER_49_1738 ();
 sg13g2_fill_1 FILLER_49_1745 ();
 sg13g2_fill_2 FILLER_49_1756 ();
 sg13g2_fill_2 FILLER_49_1763 ();
 sg13g2_fill_1 FILLER_49_1789 ();
 sg13g2_decap_8 FILLER_49_1795 ();
 sg13g2_decap_8 FILLER_49_1802 ();
 sg13g2_decap_8 FILLER_49_1809 ();
 sg13g2_fill_2 FILLER_49_1816 ();
 sg13g2_fill_1 FILLER_49_1818 ();
 sg13g2_decap_4 FILLER_49_1828 ();
 sg13g2_fill_1 FILLER_49_1832 ();
 sg13g2_fill_2 FILLER_49_1841 ();
 sg13g2_decap_4 FILLER_49_1851 ();
 sg13g2_fill_1 FILLER_49_1860 ();
 sg13g2_fill_1 FILLER_49_1865 ();
 sg13g2_fill_1 FILLER_49_1871 ();
 sg13g2_decap_4 FILLER_49_1886 ();
 sg13g2_fill_1 FILLER_49_1890 ();
 sg13g2_decap_8 FILLER_49_1903 ();
 sg13g2_decap_4 FILLER_49_1910 ();
 sg13g2_fill_2 FILLER_49_1914 ();
 sg13g2_decap_8 FILLER_49_1958 ();
 sg13g2_fill_2 FILLER_49_1965 ();
 sg13g2_fill_1 FILLER_49_1976 ();
 sg13g2_decap_4 FILLER_49_1986 ();
 sg13g2_fill_1 FILLER_49_1990 ();
 sg13g2_fill_1 FILLER_49_1999 ();
 sg13g2_decap_8 FILLER_49_2004 ();
 sg13g2_fill_1 FILLER_49_2011 ();
 sg13g2_fill_1 FILLER_49_2095 ();
 sg13g2_fill_2 FILLER_49_2135 ();
 sg13g2_fill_1 FILLER_49_2137 ();
 sg13g2_decap_4 FILLER_49_2169 ();
 sg13g2_fill_1 FILLER_49_2177 ();
 sg13g2_decap_8 FILLER_49_2183 ();
 sg13g2_fill_2 FILLER_49_2255 ();
 sg13g2_fill_1 FILLER_49_2257 ();
 sg13g2_decap_4 FILLER_49_2264 ();
 sg13g2_fill_2 FILLER_49_2278 ();
 sg13g2_fill_1 FILLER_49_2280 ();
 sg13g2_fill_2 FILLER_49_2291 ();
 sg13g2_decap_4 FILLER_49_2302 ();
 sg13g2_fill_2 FILLER_49_2316 ();
 sg13g2_fill_1 FILLER_49_2323 ();
 sg13g2_decap_8 FILLER_49_2328 ();
 sg13g2_fill_2 FILLER_49_2335 ();
 sg13g2_fill_1 FILLER_49_2337 ();
 sg13g2_fill_1 FILLER_49_2381 ();
 sg13g2_fill_1 FILLER_49_2404 ();
 sg13g2_fill_2 FILLER_49_2409 ();
 sg13g2_decap_8 FILLER_49_2424 ();
 sg13g2_fill_2 FILLER_49_2431 ();
 sg13g2_decap_8 FILLER_49_2437 ();
 sg13g2_decap_4 FILLER_49_2444 ();
 sg13g2_fill_1 FILLER_49_2488 ();
 sg13g2_fill_1 FILLER_49_2554 ();
 sg13g2_fill_2 FILLER_49_2560 ();
 sg13g2_fill_1 FILLER_49_2562 ();
 sg13g2_decap_8 FILLER_49_2568 ();
 sg13g2_decap_8 FILLER_49_2575 ();
 sg13g2_decap_8 FILLER_49_2582 ();
 sg13g2_decap_8 FILLER_49_2589 ();
 sg13g2_decap_8 FILLER_49_2596 ();
 sg13g2_decap_4 FILLER_49_2607 ();
 sg13g2_fill_2 FILLER_49_2611 ();
 sg13g2_decap_8 FILLER_49_2617 ();
 sg13g2_decap_8 FILLER_49_2624 ();
 sg13g2_decap_8 FILLER_49_2631 ();
 sg13g2_decap_8 FILLER_49_2638 ();
 sg13g2_decap_8 FILLER_49_2645 ();
 sg13g2_decap_8 FILLER_49_2652 ();
 sg13g2_decap_8 FILLER_49_2659 ();
 sg13g2_decap_4 FILLER_49_2666 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_1 FILLER_50_18 ();
 sg13g2_fill_1 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_78 ();
 sg13g2_fill_1 FILLER_50_84 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_fill_1 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_124 ();
 sg13g2_fill_2 FILLER_50_211 ();
 sg13g2_fill_1 FILLER_50_213 ();
 sg13g2_decap_4 FILLER_50_218 ();
 sg13g2_fill_2 FILLER_50_222 ();
 sg13g2_decap_4 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_267 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_301 ();
 sg13g2_fill_2 FILLER_50_324 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_fill_2 FILLER_50_354 ();
 sg13g2_fill_1 FILLER_50_359 ();
 sg13g2_fill_1 FILLER_50_375 ();
 sg13g2_fill_1 FILLER_50_381 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_fill_2 FILLER_50_420 ();
 sg13g2_fill_1 FILLER_50_427 ();
 sg13g2_fill_1 FILLER_50_455 ();
 sg13g2_fill_2 FILLER_50_493 ();
 sg13g2_fill_2 FILLER_50_502 ();
 sg13g2_fill_1 FILLER_50_578 ();
 sg13g2_fill_1 FILLER_50_585 ();
 sg13g2_fill_1 FILLER_50_600 ();
 sg13g2_decap_8 FILLER_50_645 ();
 sg13g2_decap_8 FILLER_50_652 ();
 sg13g2_decap_8 FILLER_50_659 ();
 sg13g2_decap_8 FILLER_50_666 ();
 sg13g2_decap_4 FILLER_50_673 ();
 sg13g2_fill_1 FILLER_50_708 ();
 sg13g2_fill_1 FILLER_50_728 ();
 sg13g2_fill_1 FILLER_50_733 ();
 sg13g2_fill_2 FILLER_50_760 ();
 sg13g2_fill_1 FILLER_50_762 ();
 sg13g2_fill_2 FILLER_50_771 ();
 sg13g2_fill_1 FILLER_50_773 ();
 sg13g2_fill_2 FILLER_50_782 ();
 sg13g2_fill_1 FILLER_50_784 ();
 sg13g2_fill_2 FILLER_50_790 ();
 sg13g2_fill_1 FILLER_50_792 ();
 sg13g2_fill_1 FILLER_50_801 ();
 sg13g2_fill_2 FILLER_50_836 ();
 sg13g2_decap_4 FILLER_50_854 ();
 sg13g2_fill_1 FILLER_50_868 ();
 sg13g2_decap_4 FILLER_50_895 ();
 sg13g2_fill_2 FILLER_50_899 ();
 sg13g2_fill_1 FILLER_50_927 ();
 sg13g2_fill_1 FILLER_50_970 ();
 sg13g2_fill_2 FILLER_50_991 ();
 sg13g2_decap_4 FILLER_50_1027 ();
 sg13g2_decap_4 FILLER_50_1038 ();
 sg13g2_decap_4 FILLER_50_1076 ();
 sg13g2_fill_2 FILLER_50_1123 ();
 sg13g2_fill_2 FILLER_50_1151 ();
 sg13g2_fill_2 FILLER_50_1219 ();
 sg13g2_fill_1 FILLER_50_1221 ();
 sg13g2_fill_2 FILLER_50_1232 ();
 sg13g2_fill_1 FILLER_50_1234 ();
 sg13g2_decap_8 FILLER_50_1255 ();
 sg13g2_fill_2 FILLER_50_1262 ();
 sg13g2_fill_2 FILLER_50_1268 ();
 sg13g2_fill_1 FILLER_50_1270 ();
 sg13g2_fill_2 FILLER_50_1307 ();
 sg13g2_decap_8 FILLER_50_1314 ();
 sg13g2_decap_8 FILLER_50_1321 ();
 sg13g2_decap_4 FILLER_50_1328 ();
 sg13g2_decap_4 FILLER_50_1349 ();
 sg13g2_fill_2 FILLER_50_1353 ();
 sg13g2_decap_4 FILLER_50_1360 ();
 sg13g2_fill_1 FILLER_50_1364 ();
 sg13g2_decap_4 FILLER_50_1370 ();
 sg13g2_fill_1 FILLER_50_1374 ();
 sg13g2_decap_4 FILLER_50_1381 ();
 sg13g2_decap_4 FILLER_50_1421 ();
 sg13g2_fill_2 FILLER_50_1429 ();
 sg13g2_fill_1 FILLER_50_1431 ();
 sg13g2_fill_1 FILLER_50_1450 ();
 sg13g2_fill_2 FILLER_50_1459 ();
 sg13g2_fill_2 FILLER_50_1465 ();
 sg13g2_fill_2 FILLER_50_1489 ();
 sg13g2_fill_1 FILLER_50_1491 ();
 sg13g2_decap_8 FILLER_50_1522 ();
 sg13g2_decap_8 FILLER_50_1539 ();
 sg13g2_decap_8 FILLER_50_1546 ();
 sg13g2_fill_1 FILLER_50_1553 ();
 sg13g2_fill_1 FILLER_50_1558 ();
 sg13g2_decap_4 FILLER_50_1571 ();
 sg13g2_fill_2 FILLER_50_1575 ();
 sg13g2_fill_2 FILLER_50_1586 ();
 sg13g2_fill_2 FILLER_50_1612 ();
 sg13g2_fill_1 FILLER_50_1614 ();
 sg13g2_fill_2 FILLER_50_1620 ();
 sg13g2_fill_1 FILLER_50_1627 ();
 sg13g2_decap_4 FILLER_50_1643 ();
 sg13g2_fill_2 FILLER_50_1647 ();
 sg13g2_decap_8 FILLER_50_1673 ();
 sg13g2_decap_4 FILLER_50_1680 ();
 sg13g2_decap_4 FILLER_50_1715 ();
 sg13g2_fill_1 FILLER_50_1719 ();
 sg13g2_decap_4 FILLER_50_1728 ();
 sg13g2_fill_2 FILLER_50_1751 ();
 sg13g2_fill_2 FILLER_50_1757 ();
 sg13g2_decap_8 FILLER_50_1764 ();
 sg13g2_decap_8 FILLER_50_1771 ();
 sg13g2_decap_4 FILLER_50_1778 ();
 sg13g2_fill_1 FILLER_50_1782 ();
 sg13g2_fill_1 FILLER_50_1796 ();
 sg13g2_fill_1 FILLER_50_1802 ();
 sg13g2_fill_1 FILLER_50_1807 ();
 sg13g2_decap_4 FILLER_50_1817 ();
 sg13g2_fill_1 FILLER_50_1821 ();
 sg13g2_decap_4 FILLER_50_1826 ();
 sg13g2_fill_1 FILLER_50_1849 ();
 sg13g2_fill_1 FILLER_50_1854 ();
 sg13g2_fill_2 FILLER_50_1882 ();
 sg13g2_decap_8 FILLER_50_1915 ();
 sg13g2_fill_2 FILLER_50_1922 ();
 sg13g2_fill_1 FILLER_50_1924 ();
 sg13g2_decap_8 FILLER_50_1981 ();
 sg13g2_fill_2 FILLER_50_1988 ();
 sg13g2_fill_1 FILLER_50_1990 ();
 sg13g2_decap_8 FILLER_50_1996 ();
 sg13g2_decap_8 FILLER_50_2003 ();
 sg13g2_decap_4 FILLER_50_2010 ();
 sg13g2_fill_1 FILLER_50_2014 ();
 sg13g2_decap_8 FILLER_50_2029 ();
 sg13g2_decap_8 FILLER_50_2036 ();
 sg13g2_fill_2 FILLER_50_2079 ();
 sg13g2_fill_2 FILLER_50_2085 ();
 sg13g2_fill_1 FILLER_50_2123 ();
 sg13g2_fill_1 FILLER_50_2128 ();
 sg13g2_decap_8 FILLER_50_2191 ();
 sg13g2_decap_4 FILLER_50_2198 ();
 sg13g2_fill_1 FILLER_50_2202 ();
 sg13g2_decap_4 FILLER_50_2207 ();
 sg13g2_decap_4 FILLER_50_2228 ();
 sg13g2_decap_8 FILLER_50_2236 ();
 sg13g2_decap_8 FILLER_50_2243 ();
 sg13g2_decap_8 FILLER_50_2250 ();
 sg13g2_decap_8 FILLER_50_2267 ();
 sg13g2_fill_2 FILLER_50_2274 ();
 sg13g2_decap_8 FILLER_50_2312 ();
 sg13g2_decap_8 FILLER_50_2319 ();
 sg13g2_decap_8 FILLER_50_2326 ();
 sg13g2_fill_2 FILLER_50_2333 ();
 sg13g2_fill_1 FILLER_50_2335 ();
 sg13g2_decap_8 FILLER_50_2340 ();
 sg13g2_decap_4 FILLER_50_2347 ();
 sg13g2_fill_1 FILLER_50_2351 ();
 sg13g2_fill_1 FILLER_50_2381 ();
 sg13g2_decap_8 FILLER_50_2425 ();
 sg13g2_fill_2 FILLER_50_2432 ();
 sg13g2_fill_1 FILLER_50_2448 ();
 sg13g2_decap_4 FILLER_50_2457 ();
 sg13g2_fill_2 FILLER_50_2461 ();
 sg13g2_fill_2 FILLER_50_2473 ();
 sg13g2_fill_1 FILLER_50_2475 ();
 sg13g2_fill_1 FILLER_50_2509 ();
 sg13g2_fill_2 FILLER_50_2515 ();
 sg13g2_fill_2 FILLER_50_2566 ();
 sg13g2_decap_8 FILLER_50_2572 ();
 sg13g2_decap_8 FILLER_50_2579 ();
 sg13g2_fill_2 FILLER_50_2586 ();
 sg13g2_decap_8 FILLER_50_2630 ();
 sg13g2_decap_8 FILLER_50_2637 ();
 sg13g2_decap_8 FILLER_50_2644 ();
 sg13g2_decap_8 FILLER_50_2651 ();
 sg13g2_decap_8 FILLER_50_2658 ();
 sg13g2_decap_4 FILLER_50_2665 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_fill_1 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_33 ();
 sg13g2_fill_1 FILLER_51_43 ();
 sg13g2_fill_1 FILLER_51_49 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_fill_2 FILLER_51_100 ();
 sg13g2_fill_2 FILLER_51_128 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_153 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_decap_4 FILLER_51_228 ();
 sg13g2_fill_2 FILLER_51_232 ();
 sg13g2_fill_1 FILLER_51_244 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_1 FILLER_51_252 ();
 sg13g2_fill_2 FILLER_51_279 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_336 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_374 ();
 sg13g2_decap_8 FILLER_51_451 ();
 sg13g2_decap_4 FILLER_51_464 ();
 sg13g2_fill_1 FILLER_51_468 ();
 sg13g2_decap_4 FILLER_51_477 ();
 sg13g2_fill_1 FILLER_51_481 ();
 sg13g2_fill_2 FILLER_51_498 ();
 sg13g2_fill_2 FILLER_51_509 ();
 sg13g2_fill_1 FILLER_51_518 ();
 sg13g2_fill_2 FILLER_51_596 ();
 sg13g2_fill_2 FILLER_51_602 ();
 sg13g2_fill_1 FILLER_51_609 ();
 sg13g2_fill_2 FILLER_51_621 ();
 sg13g2_decap_4 FILLER_51_638 ();
 sg13g2_decap_8 FILLER_51_646 ();
 sg13g2_fill_2 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_660 ();
 sg13g2_decap_4 FILLER_51_667 ();
 sg13g2_fill_2 FILLER_51_671 ();
 sg13g2_fill_1 FILLER_51_692 ();
 sg13g2_fill_1 FILLER_51_777 ();
 sg13g2_fill_1 FILLER_51_803 ();
 sg13g2_fill_2 FILLER_51_809 ();
 sg13g2_fill_1 FILLER_51_811 ();
 sg13g2_fill_2 FILLER_51_816 ();
 sg13g2_fill_1 FILLER_51_818 ();
 sg13g2_fill_2 FILLER_51_823 ();
 sg13g2_fill_1 FILLER_51_829 ();
 sg13g2_decap_8 FILLER_51_834 ();
 sg13g2_decap_4 FILLER_51_841 ();
 sg13g2_fill_1 FILLER_51_866 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_fill_2 FILLER_51_884 ();
 sg13g2_decap_8 FILLER_51_890 ();
 sg13g2_decap_8 FILLER_51_897 ();
 sg13g2_fill_2 FILLER_51_904 ();
 sg13g2_fill_1 FILLER_51_906 ();
 sg13g2_fill_2 FILLER_51_911 ();
 sg13g2_decap_8 FILLER_51_937 ();
 sg13g2_fill_1 FILLER_51_944 ();
 sg13g2_decap_8 FILLER_51_948 ();
 sg13g2_fill_2 FILLER_51_955 ();
 sg13g2_fill_1 FILLER_51_963 ();
 sg13g2_fill_2 FILLER_51_993 ();
 sg13g2_fill_2 FILLER_51_1007 ();
 sg13g2_fill_2 FILLER_51_1017 ();
 sg13g2_fill_2 FILLER_51_1024 ();
 sg13g2_fill_1 FILLER_51_1030 ();
 sg13g2_fill_1 FILLER_51_1067 ();
 sg13g2_fill_2 FILLER_51_1104 ();
 sg13g2_fill_1 FILLER_51_1106 ();
 sg13g2_decap_4 FILLER_51_1117 ();
 sg13g2_fill_1 FILLER_51_1125 ();
 sg13g2_decap_8 FILLER_51_1140 ();
 sg13g2_fill_2 FILLER_51_1147 ();
 sg13g2_fill_1 FILLER_51_1169 ();
 sg13g2_decap_8 FILLER_51_1174 ();
 sg13g2_decap_8 FILLER_51_1181 ();
 sg13g2_fill_2 FILLER_51_1188 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_fill_1 FILLER_51_1201 ();
 sg13g2_fill_1 FILLER_51_1206 ();
 sg13g2_fill_1 FILLER_51_1223 ();
 sg13g2_fill_2 FILLER_51_1237 ();
 sg13g2_fill_1 FILLER_51_1248 ();
 sg13g2_fill_1 FILLER_51_1258 ();
 sg13g2_fill_2 FILLER_51_1282 ();
 sg13g2_fill_1 FILLER_51_1284 ();
 sg13g2_fill_2 FILLER_51_1291 ();
 sg13g2_fill_2 FILLER_51_1299 ();
 sg13g2_decap_4 FILLER_51_1317 ();
 sg13g2_fill_1 FILLER_51_1321 ();
 sg13g2_fill_1 FILLER_51_1334 ();
 sg13g2_fill_2 FILLER_51_1350 ();
 sg13g2_fill_1 FILLER_51_1352 ();
 sg13g2_decap_8 FILLER_51_1363 ();
 sg13g2_decap_8 FILLER_51_1370 ();
 sg13g2_decap_8 FILLER_51_1377 ();
 sg13g2_fill_1 FILLER_51_1384 ();
 sg13g2_decap_4 FILLER_51_1388 ();
 sg13g2_decap_4 FILLER_51_1396 ();
 sg13g2_fill_2 FILLER_51_1400 ();
 sg13g2_fill_2 FILLER_51_1432 ();
 sg13g2_decap_4 FILLER_51_1438 ();
 sg13g2_fill_1 FILLER_51_1459 ();
 sg13g2_fill_1 FILLER_51_1475 ();
 sg13g2_decap_4 FILLER_51_1481 ();
 sg13g2_fill_2 FILLER_51_1489 ();
 sg13g2_decap_8 FILLER_51_1500 ();
 sg13g2_decap_8 FILLER_51_1511 ();
 sg13g2_fill_1 FILLER_51_1518 ();
 sg13g2_fill_1 FILLER_51_1523 ();
 sg13g2_fill_2 FILLER_51_1528 ();
 sg13g2_fill_1 FILLER_51_1530 ();
 sg13g2_fill_2 FILLER_51_1536 ();
 sg13g2_fill_1 FILLER_51_1551 ();
 sg13g2_fill_1 FILLER_51_1557 ();
 sg13g2_fill_2 FILLER_51_1562 ();
 sg13g2_fill_2 FILLER_51_1569 ();
 sg13g2_fill_2 FILLER_51_1575 ();
 sg13g2_fill_1 FILLER_51_1586 ();
 sg13g2_fill_1 FILLER_51_1636 ();
 sg13g2_decap_4 FILLER_51_1641 ();
 sg13g2_fill_1 FILLER_51_1653 ();
 sg13g2_fill_1 FILLER_51_1671 ();
 sg13g2_decap_8 FILLER_51_1693 ();
 sg13g2_decap_8 FILLER_51_1700 ();
 sg13g2_decap_8 FILLER_51_1707 ();
 sg13g2_decap_4 FILLER_51_1714 ();
 sg13g2_fill_1 FILLER_51_1727 ();
 sg13g2_fill_2 FILLER_51_1735 ();
 sg13g2_fill_2 FILLER_51_1749 ();
 sg13g2_decap_4 FILLER_51_1755 ();
 sg13g2_fill_2 FILLER_51_1759 ();
 sg13g2_decap_8 FILLER_51_1765 ();
 sg13g2_decap_8 FILLER_51_1772 ();
 sg13g2_decap_8 FILLER_51_1779 ();
 sg13g2_decap_4 FILLER_51_1786 ();
 sg13g2_fill_2 FILLER_51_1790 ();
 sg13g2_fill_2 FILLER_51_1801 ();
 sg13g2_fill_1 FILLER_51_1803 ();
 sg13g2_fill_1 FILLER_51_1818 ();
 sg13g2_fill_2 FILLER_51_1828 ();
 sg13g2_fill_1 FILLER_51_1847 ();
 sg13g2_fill_2 FILLER_51_1865 ();
 sg13g2_fill_2 FILLER_51_1872 ();
 sg13g2_fill_1 FILLER_51_1888 ();
 sg13g2_fill_2 FILLER_51_1910 ();
 sg13g2_decap_4 FILLER_51_1916 ();
 sg13g2_decap_8 FILLER_51_1924 ();
 sg13g2_decap_8 FILLER_51_1931 ();
 sg13g2_decap_4 FILLER_51_1942 ();
 sg13g2_decap_4 FILLER_51_1958 ();
 sg13g2_fill_2 FILLER_51_1962 ();
 sg13g2_decap_8 FILLER_51_1968 ();
 sg13g2_decap_4 FILLER_51_1975 ();
 sg13g2_decap_8 FILLER_51_1984 ();
 sg13g2_decap_8 FILLER_51_1991 ();
 sg13g2_decap_8 FILLER_51_1998 ();
 sg13g2_decap_8 FILLER_51_2005 ();
 sg13g2_fill_2 FILLER_51_2081 ();
 sg13g2_decap_8 FILLER_51_2123 ();
 sg13g2_fill_2 FILLER_51_2130 ();
 sg13g2_fill_1 FILLER_51_2132 ();
 sg13g2_decap_8 FILLER_51_2173 ();
 sg13g2_decap_4 FILLER_51_2180 ();
 sg13g2_fill_2 FILLER_51_2184 ();
 sg13g2_decap_8 FILLER_51_2190 ();
 sg13g2_fill_2 FILLER_51_2197 ();
 sg13g2_fill_1 FILLER_51_2199 ();
 sg13g2_fill_2 FILLER_51_2234 ();
 sg13g2_fill_1 FILLER_51_2236 ();
 sg13g2_fill_2 FILLER_51_2267 ();
 sg13g2_decap_4 FILLER_51_2275 ();
 sg13g2_fill_1 FILLER_51_2279 ();
 sg13g2_decap_8 FILLER_51_2294 ();
 sg13g2_fill_2 FILLER_51_2301 ();
 sg13g2_decap_8 FILLER_51_2309 ();
 sg13g2_fill_2 FILLER_51_2372 ();
 sg13g2_fill_2 FILLER_51_2404 ();
 sg13g2_decap_4 FILLER_51_2412 ();
 sg13g2_decap_4 FILLER_51_2426 ();
 sg13g2_fill_2 FILLER_51_2430 ();
 sg13g2_decap_8 FILLER_51_2463 ();
 sg13g2_fill_2 FILLER_51_2470 ();
 sg13g2_fill_1 FILLER_51_2472 ();
 sg13g2_decap_8 FILLER_51_2479 ();
 sg13g2_fill_2 FILLER_51_2492 ();
 sg13g2_fill_1 FILLER_51_2507 ();
 sg13g2_fill_2 FILLER_51_2512 ();
 sg13g2_fill_1 FILLER_51_2519 ();
 sg13g2_decap_8 FILLER_51_2577 ();
 sg13g2_decap_4 FILLER_51_2584 ();
 sg13g2_fill_2 FILLER_51_2588 ();
 sg13g2_decap_8 FILLER_51_2626 ();
 sg13g2_decap_8 FILLER_51_2637 ();
 sg13g2_decap_8 FILLER_51_2644 ();
 sg13g2_decap_8 FILLER_51_2651 ();
 sg13g2_decap_8 FILLER_51_2658 ();
 sg13g2_decap_4 FILLER_51_2665 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_17 ();
 sg13g2_fill_1 FILLER_52_22 ();
 sg13g2_fill_2 FILLER_52_43 ();
 sg13g2_fill_1 FILLER_52_67 ();
 sg13g2_fill_1 FILLER_52_73 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_fill_1 FILLER_52_137 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_fill_2 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_167 ();
 sg13g2_decap_8 FILLER_52_174 ();
 sg13g2_fill_2 FILLER_52_181 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_fill_2 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_fill_1 FILLER_52_274 ();
 sg13g2_fill_2 FILLER_52_280 ();
 sg13g2_fill_1 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_fill_2 FILLER_52_334 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_fill_2 FILLER_52_364 ();
 sg13g2_fill_1 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_394 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_decap_8 FILLER_52_415 ();
 sg13g2_fill_2 FILLER_52_426 ();
 sg13g2_fill_1 FILLER_52_428 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_8 FILLER_52_457 ();
 sg13g2_decap_4 FILLER_52_464 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_decap_8 FILLER_52_474 ();
 sg13g2_decap_8 FILLER_52_481 ();
 sg13g2_decap_4 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_492 ();
 sg13g2_fill_2 FILLER_52_503 ();
 sg13g2_fill_2 FILLER_52_534 ();
 sg13g2_fill_1 FILLER_52_552 ();
 sg13g2_fill_1 FILLER_52_593 ();
 sg13g2_fill_1 FILLER_52_598 ();
 sg13g2_fill_1 FILLER_52_629 ();
 sg13g2_fill_2 FILLER_52_660 ();
 sg13g2_fill_1 FILLER_52_668 ();
 sg13g2_fill_1 FILLER_52_682 ();
 sg13g2_fill_2 FILLER_52_707 ();
 sg13g2_fill_1 FILLER_52_709 ();
 sg13g2_fill_2 FILLER_52_719 ();
 sg13g2_fill_1 FILLER_52_727 ();
 sg13g2_fill_1 FILLER_52_734 ();
 sg13g2_fill_1 FILLER_52_745 ();
 sg13g2_decap_4 FILLER_52_750 ();
 sg13g2_decap_4 FILLER_52_764 ();
 sg13g2_fill_1 FILLER_52_768 ();
 sg13g2_decap_8 FILLER_52_803 ();
 sg13g2_decap_8 FILLER_52_810 ();
 sg13g2_decap_8 FILLER_52_817 ();
 sg13g2_fill_1 FILLER_52_824 ();
 sg13g2_fill_1 FILLER_52_865 ();
 sg13g2_fill_1 FILLER_52_871 ();
 sg13g2_fill_1 FILLER_52_876 ();
 sg13g2_decap_8 FILLER_52_882 ();
 sg13g2_fill_2 FILLER_52_903 ();
 sg13g2_decap_8 FILLER_52_911 ();
 sg13g2_decap_8 FILLER_52_918 ();
 sg13g2_decap_8 FILLER_52_925 ();
 sg13g2_fill_2 FILLER_52_932 ();
 sg13g2_fill_1 FILLER_52_934 ();
 sg13g2_decap_8 FILLER_52_955 ();
 sg13g2_fill_1 FILLER_52_962 ();
 sg13g2_fill_2 FILLER_52_997 ();
 sg13g2_fill_2 FILLER_52_1029 ();
 sg13g2_decap_8 FILLER_52_1037 ();
 sg13g2_decap_4 FILLER_52_1044 ();
 sg13g2_decap_8 FILLER_52_1056 ();
 sg13g2_decap_4 FILLER_52_1063 ();
 sg13g2_fill_2 FILLER_52_1077 ();
 sg13g2_decap_4 FILLER_52_1105 ();
 sg13g2_fill_2 FILLER_52_1139 ();
 sg13g2_decap_8 FILLER_52_1207 ();
 sg13g2_decap_4 FILLER_52_1214 ();
 sg13g2_fill_1 FILLER_52_1228 ();
 sg13g2_decap_8 FILLER_52_1238 ();
 sg13g2_fill_2 FILLER_52_1245 ();
 sg13g2_fill_1 FILLER_52_1247 ();
 sg13g2_fill_1 FILLER_52_1253 ();
 sg13g2_fill_2 FILLER_52_1258 ();
 sg13g2_fill_1 FILLER_52_1260 ();
 sg13g2_decap_4 FILLER_52_1282 ();
 sg13g2_decap_8 FILLER_52_1291 ();
 sg13g2_decap_8 FILLER_52_1298 ();
 sg13g2_decap_4 FILLER_52_1305 ();
 sg13g2_fill_1 FILLER_52_1309 ();
 sg13g2_fill_2 FILLER_52_1345 ();
 sg13g2_fill_1 FILLER_52_1347 ();
 sg13g2_fill_1 FILLER_52_1381 ();
 sg13g2_fill_1 FILLER_52_1401 ();
 sg13g2_decap_8 FILLER_52_1419 ();
 sg13g2_decap_8 FILLER_52_1426 ();
 sg13g2_decap_4 FILLER_52_1433 ();
 sg13g2_fill_2 FILLER_52_1437 ();
 sg13g2_decap_4 FILLER_52_1444 ();
 sg13g2_fill_1 FILLER_52_1448 ();
 sg13g2_fill_2 FILLER_52_1476 ();
 sg13g2_decap_4 FILLER_52_1486 ();
 sg13g2_fill_2 FILLER_52_1490 ();
 sg13g2_decap_8 FILLER_52_1505 ();
 sg13g2_decap_8 FILLER_52_1512 ();
 sg13g2_decap_8 FILLER_52_1519 ();
 sg13g2_decap_8 FILLER_52_1526 ();
 sg13g2_decap_8 FILLER_52_1533 ();
 sg13g2_decap_8 FILLER_52_1540 ();
 sg13g2_fill_2 FILLER_52_1562 ();
 sg13g2_fill_2 FILLER_52_1584 ();
 sg13g2_decap_8 FILLER_52_1596 ();
 sg13g2_fill_2 FILLER_52_1603 ();
 sg13g2_fill_1 FILLER_52_1605 ();
 sg13g2_fill_2 FILLER_52_1623 ();
 sg13g2_decap_4 FILLER_52_1632 ();
 sg13g2_decap_4 FILLER_52_1640 ();
 sg13g2_fill_2 FILLER_52_1644 ();
 sg13g2_decap_8 FILLER_52_1665 ();
 sg13g2_decap_4 FILLER_52_1672 ();
 sg13g2_decap_8 FILLER_52_1685 ();
 sg13g2_decap_8 FILLER_52_1692 ();
 sg13g2_decap_8 FILLER_52_1699 ();
 sg13g2_decap_8 FILLER_52_1706 ();
 sg13g2_fill_1 FILLER_52_1713 ();
 sg13g2_fill_2 FILLER_52_1733 ();
 sg13g2_fill_2 FILLER_52_1740 ();
 sg13g2_decap_8 FILLER_52_1757 ();
 sg13g2_decap_8 FILLER_52_1764 ();
 sg13g2_decap_4 FILLER_52_1771 ();
 sg13g2_fill_1 FILLER_52_1775 ();
 sg13g2_fill_2 FILLER_52_1780 ();
 sg13g2_fill_1 FILLER_52_1782 ();
 sg13g2_fill_1 FILLER_52_1798 ();
 sg13g2_decap_4 FILLER_52_1825 ();
 sg13g2_fill_1 FILLER_52_1833 ();
 sg13g2_fill_2 FILLER_52_1840 ();
 sg13g2_fill_1 FILLER_52_1842 ();
 sg13g2_fill_2 FILLER_52_1848 ();
 sg13g2_fill_1 FILLER_52_1854 ();
 sg13g2_fill_2 FILLER_52_1866 ();
 sg13g2_fill_2 FILLER_52_1891 ();
 sg13g2_fill_1 FILLER_52_1893 ();
 sg13g2_decap_8 FILLER_52_1923 ();
 sg13g2_fill_1 FILLER_52_1930 ();
 sg13g2_decap_4 FILLER_52_1960 ();
 sg13g2_fill_1 FILLER_52_1964 ();
 sg13g2_decap_4 FILLER_52_1971 ();
 sg13g2_decap_8 FILLER_52_2013 ();
 sg13g2_decap_8 FILLER_52_2020 ();
 sg13g2_fill_2 FILLER_52_2027 ();
 sg13g2_fill_1 FILLER_52_2029 ();
 sg13g2_decap_8 FILLER_52_2034 ();
 sg13g2_decap_4 FILLER_52_2041 ();
 sg13g2_fill_2 FILLER_52_2045 ();
 sg13g2_fill_2 FILLER_52_2087 ();
 sg13g2_fill_1 FILLER_52_2089 ();
 sg13g2_decap_4 FILLER_52_2126 ();
 sg13g2_fill_2 FILLER_52_2130 ();
 sg13g2_decap_8 FILLER_52_2162 ();
 sg13g2_fill_2 FILLER_52_2169 ();
 sg13g2_fill_1 FILLER_52_2171 ();
 sg13g2_fill_2 FILLER_52_2284 ();
 sg13g2_decap_4 FILLER_52_2338 ();
 sg13g2_fill_2 FILLER_52_2342 ();
 sg13g2_decap_8 FILLER_52_2419 ();
 sg13g2_fill_2 FILLER_52_2426 ();
 sg13g2_fill_1 FILLER_52_2428 ();
 sg13g2_decap_8 FILLER_52_2468 ();
 sg13g2_decap_8 FILLER_52_2475 ();
 sg13g2_decap_4 FILLER_52_2482 ();
 sg13g2_fill_1 FILLER_52_2531 ();
 sg13g2_fill_2 FILLER_52_2589 ();
 sg13g2_fill_1 FILLER_52_2591 ();
 sg13g2_fill_2 FILLER_52_2626 ();
 sg13g2_decap_8 FILLER_52_2654 ();
 sg13g2_decap_8 FILLER_52_2661 ();
 sg13g2_fill_2 FILLER_52_2668 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_39 ();
 sg13g2_decap_4 FILLER_53_46 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_fill_2 FILLER_53_60 ();
 sg13g2_fill_2 FILLER_53_76 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_83 ();
 sg13g2_decap_4 FILLER_53_99 ();
 sg13g2_fill_2 FILLER_53_113 ();
 sg13g2_fill_1 FILLER_53_115 ();
 sg13g2_decap_8 FILLER_53_151 ();
 sg13g2_decap_8 FILLER_53_158 ();
 sg13g2_fill_2 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_231 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_fill_2 FILLER_53_242 ();
 sg13g2_fill_2 FILLER_53_248 ();
 sg13g2_fill_1 FILLER_53_250 ();
 sg13g2_fill_2 FILLER_53_255 ();
 sg13g2_fill_2 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_decap_4 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_286 ();
 sg13g2_fill_1 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_349 ();
 sg13g2_decap_8 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_363 ();
 sg13g2_fill_2 FILLER_53_370 ();
 sg13g2_fill_2 FILLER_53_381 ();
 sg13g2_fill_1 FILLER_53_387 ();
 sg13g2_decap_4 FILLER_53_392 ();
 sg13g2_fill_1 FILLER_53_396 ();
 sg13g2_fill_1 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_410 ();
 sg13g2_fill_2 FILLER_53_417 ();
 sg13g2_fill_1 FILLER_53_419 ();
 sg13g2_decap_8 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_432 ();
 sg13g2_fill_2 FILLER_53_438 ();
 sg13g2_fill_2 FILLER_53_445 ();
 sg13g2_fill_1 FILLER_53_451 ();
 sg13g2_fill_1 FILLER_53_462 ();
 sg13g2_fill_1 FILLER_53_469 ();
 sg13g2_fill_1 FILLER_53_476 ();
 sg13g2_fill_2 FILLER_53_503 ();
 sg13g2_fill_1 FILLER_53_511 ();
 sg13g2_decap_8 FILLER_53_518 ();
 sg13g2_fill_1 FILLER_53_525 ();
 sg13g2_decap_4 FILLER_53_530 ();
 sg13g2_fill_1 FILLER_53_559 ();
 sg13g2_fill_2 FILLER_53_572 ();
 sg13g2_fill_1 FILLER_53_615 ();
 sg13g2_fill_1 FILLER_53_626 ();
 sg13g2_fill_1 FILLER_53_636 ();
 sg13g2_decap_8 FILLER_53_673 ();
 sg13g2_decap_4 FILLER_53_680 ();
 sg13g2_fill_2 FILLER_53_688 ();
 sg13g2_fill_2 FILLER_53_694 ();
 sg13g2_fill_2 FILLER_53_701 ();
 sg13g2_fill_1 FILLER_53_703 ();
 sg13g2_fill_1 FILLER_53_712 ();
 sg13g2_fill_2 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_720 ();
 sg13g2_fill_1 FILLER_53_732 ();
 sg13g2_fill_1 FILLER_53_741 ();
 sg13g2_decap_4 FILLER_53_746 ();
 sg13g2_fill_2 FILLER_53_750 ();
 sg13g2_decap_4 FILLER_53_757 ();
 sg13g2_fill_2 FILLER_53_761 ();
 sg13g2_fill_2 FILLER_53_825 ();
 sg13g2_decap_4 FILLER_53_841 ();
 sg13g2_decap_8 FILLER_53_865 ();
 sg13g2_decap_8 FILLER_53_872 ();
 sg13g2_decap_4 FILLER_53_879 ();
 sg13g2_fill_2 FILLER_53_883 ();
 sg13g2_decap_8 FILLER_53_917 ();
 sg13g2_fill_1 FILLER_53_924 ();
 sg13g2_fill_2 FILLER_53_935 ();
 sg13g2_fill_2 FILLER_53_963 ();
 sg13g2_fill_1 FILLER_53_1025 ();
 sg13g2_decap_8 FILLER_53_1062 ();
 sg13g2_decap_4 FILLER_53_1069 ();
 sg13g2_fill_1 FILLER_53_1073 ();
 sg13g2_decap_8 FILLER_53_1092 ();
 sg13g2_fill_2 FILLER_53_1099 ();
 sg13g2_fill_1 FILLER_53_1101 ();
 sg13g2_decap_4 FILLER_53_1112 ();
 sg13g2_fill_1 FILLER_53_1116 ();
 sg13g2_fill_1 FILLER_53_1121 ();
 sg13g2_fill_1 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1170 ();
 sg13g2_fill_2 FILLER_53_1187 ();
 sg13g2_fill_1 FILLER_53_1219 ();
 sg13g2_decap_4 FILLER_53_1226 ();
 sg13g2_fill_2 FILLER_53_1230 ();
 sg13g2_fill_1 FILLER_53_1242 ();
 sg13g2_fill_1 FILLER_53_1273 ();
 sg13g2_fill_2 FILLER_53_1277 ();
 sg13g2_decap_8 FILLER_53_1297 ();
 sg13g2_fill_2 FILLER_53_1304 ();
 sg13g2_fill_1 FILLER_53_1306 ();
 sg13g2_fill_2 FILLER_53_1329 ();
 sg13g2_decap_8 FILLER_53_1406 ();
 sg13g2_fill_2 FILLER_53_1413 ();
 sg13g2_decap_4 FILLER_53_1442 ();
 sg13g2_fill_1 FILLER_53_1450 ();
 sg13g2_fill_2 FILLER_53_1467 ();
 sg13g2_fill_1 FILLER_53_1469 ();
 sg13g2_decap_8 FILLER_53_1507 ();
 sg13g2_decap_8 FILLER_53_1514 ();
 sg13g2_decap_8 FILLER_53_1521 ();
 sg13g2_decap_8 FILLER_53_1532 ();
 sg13g2_fill_1 FILLER_53_1539 ();
 sg13g2_decap_4 FILLER_53_1566 ();
 sg13g2_fill_1 FILLER_53_1570 ();
 sg13g2_fill_2 FILLER_53_1585 ();
 sg13g2_fill_1 FILLER_53_1592 ();
 sg13g2_fill_2 FILLER_53_1630 ();
 sg13g2_fill_1 FILLER_53_1632 ();
 sg13g2_decap_8 FILLER_53_1663 ();
 sg13g2_fill_1 FILLER_53_1670 ();
 sg13g2_decap_8 FILLER_53_1705 ();
 sg13g2_decap_8 FILLER_53_1712 ();
 sg13g2_fill_1 FILLER_53_1719 ();
 sg13g2_decap_8 FILLER_53_1724 ();
 sg13g2_fill_1 FILLER_53_1762 ();
 sg13g2_fill_1 FILLER_53_1771 ();
 sg13g2_decap_4 FILLER_53_1780 ();
 sg13g2_fill_1 FILLER_53_1784 ();
 sg13g2_decap_4 FILLER_53_1794 ();
 sg13g2_decap_8 FILLER_53_1803 ();
 sg13g2_fill_2 FILLER_53_1810 ();
 sg13g2_fill_1 FILLER_53_1812 ();
 sg13g2_decap_4 FILLER_53_1817 ();
 sg13g2_fill_1 FILLER_53_1821 ();
 sg13g2_fill_2 FILLER_53_1827 ();
 sg13g2_decap_8 FILLER_53_1833 ();
 sg13g2_fill_1 FILLER_53_1840 ();
 sg13g2_fill_1 FILLER_53_1873 ();
 sg13g2_decap_4 FILLER_53_1880 ();
 sg13g2_fill_1 FILLER_53_1890 ();
 sg13g2_decap_4 FILLER_53_1927 ();
 sg13g2_fill_2 FILLER_53_1931 ();
 sg13g2_decap_4 FILLER_53_1943 ();
 sg13g2_fill_2 FILLER_53_1947 ();
 sg13g2_fill_1 FILLER_53_2006 ();
 sg13g2_decap_8 FILLER_53_2012 ();
 sg13g2_decap_4 FILLER_53_2019 ();
 sg13g2_fill_1 FILLER_53_2023 ();
 sg13g2_decap_4 FILLER_53_2028 ();
 sg13g2_decap_4 FILLER_53_2035 ();
 sg13g2_fill_2 FILLER_53_2039 ();
 sg13g2_decap_8 FILLER_53_2049 ();
 sg13g2_decap_8 FILLER_53_2056 ();
 sg13g2_decap_4 FILLER_53_2063 ();
 sg13g2_fill_1 FILLER_53_2067 ();
 sg13g2_decap_8 FILLER_53_2072 ();
 sg13g2_decap_4 FILLER_53_2079 ();
 sg13g2_fill_2 FILLER_53_2083 ();
 sg13g2_decap_8 FILLER_53_2112 ();
 sg13g2_decap_8 FILLER_53_2119 ();
 sg13g2_decap_4 FILLER_53_2136 ();
 sg13g2_fill_2 FILLER_53_2144 ();
 sg13g2_fill_1 FILLER_53_2150 ();
 sg13g2_decap_8 FILLER_53_2154 ();
 sg13g2_decap_8 FILLER_53_2161 ();
 sg13g2_decap_8 FILLER_53_2168 ();
 sg13g2_decap_4 FILLER_53_2175 ();
 sg13g2_fill_1 FILLER_53_2179 ();
 sg13g2_fill_1 FILLER_53_2228 ();
 sg13g2_decap_8 FILLER_53_2245 ();
 sg13g2_decap_8 FILLER_53_2252 ();
 sg13g2_decap_8 FILLER_53_2259 ();
 sg13g2_fill_1 FILLER_53_2315 ();
 sg13g2_fill_1 FILLER_53_2326 ();
 sg13g2_fill_2 FILLER_53_2376 ();
 sg13g2_fill_1 FILLER_53_2381 ();
 sg13g2_fill_1 FILLER_53_2395 ();
 sg13g2_fill_2 FILLER_53_2426 ();
 sg13g2_fill_1 FILLER_53_2434 ();
 sg13g2_fill_2 FILLER_53_2449 ();
 sg13g2_fill_1 FILLER_53_2451 ();
 sg13g2_fill_2 FILLER_53_2478 ();
 sg13g2_fill_2 FILLER_53_2506 ();
 sg13g2_fill_2 FILLER_53_2543 ();
 sg13g2_fill_1 FILLER_53_2545 ();
 sg13g2_decap_8 FILLER_53_2597 ();
 sg13g2_decap_8 FILLER_53_2604 ();
 sg13g2_decap_8 FILLER_53_2611 ();
 sg13g2_decap_8 FILLER_53_2618 ();
 sg13g2_decap_8 FILLER_53_2625 ();
 sg13g2_decap_8 FILLER_53_2632 ();
 sg13g2_decap_8 FILLER_53_2639 ();
 sg13g2_decap_8 FILLER_53_2646 ();
 sg13g2_decap_8 FILLER_53_2653 ();
 sg13g2_decap_8 FILLER_53_2660 ();
 sg13g2_fill_2 FILLER_53_2667 ();
 sg13g2_fill_1 FILLER_53_2669 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_13 ();
 sg13g2_fill_1 FILLER_54_15 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_52 ();
 sg13g2_decap_8 FILLER_54_78 ();
 sg13g2_fill_2 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_87 ();
 sg13g2_decap_4 FILLER_54_118 ();
 sg13g2_fill_1 FILLER_54_135 ();
 sg13g2_fill_2 FILLER_54_148 ();
 sg13g2_fill_1 FILLER_54_155 ();
 sg13g2_fill_2 FILLER_54_177 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_2 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_368 ();
 sg13g2_decap_8 FILLER_54_375 ();
 sg13g2_fill_2 FILLER_54_417 ();
 sg13g2_fill_1 FILLER_54_419 ();
 sg13g2_decap_4 FILLER_54_425 ();
 sg13g2_fill_2 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_54_466 ();
 sg13g2_fill_1 FILLER_54_508 ();
 sg13g2_decap_4 FILLER_54_519 ();
 sg13g2_fill_2 FILLER_54_523 ();
 sg13g2_decap_4 FILLER_54_529 ();
 sg13g2_fill_1 FILLER_54_533 ();
 sg13g2_fill_2 FILLER_54_552 ();
 sg13g2_fill_1 FILLER_54_559 ();
 sg13g2_fill_2 FILLER_54_621 ();
 sg13g2_decap_4 FILLER_54_627 ();
 sg13g2_fill_2 FILLER_54_636 ();
 sg13g2_fill_1 FILLER_54_638 ();
 sg13g2_fill_2 FILLER_54_657 ();
 sg13g2_fill_1 FILLER_54_675 ();
 sg13g2_fill_2 FILLER_54_721 ();
 sg13g2_fill_1 FILLER_54_723 ();
 sg13g2_fill_2 FILLER_54_750 ();
 sg13g2_fill_1 FILLER_54_752 ();
 sg13g2_fill_2 FILLER_54_757 ();
 sg13g2_fill_2 FILLER_54_769 ();
 sg13g2_fill_1 FILLER_54_789 ();
 sg13g2_fill_2 FILLER_54_794 ();
 sg13g2_decap_8 FILLER_54_810 ();
 sg13g2_fill_2 FILLER_54_817 ();
 sg13g2_fill_2 FILLER_54_855 ();
 sg13g2_fill_1 FILLER_54_857 ();
 sg13g2_fill_1 FILLER_54_866 ();
 sg13g2_decap_8 FILLER_54_883 ();
 sg13g2_fill_1 FILLER_54_920 ();
 sg13g2_decap_4 FILLER_54_931 ();
 sg13g2_fill_2 FILLER_54_938 ();
 sg13g2_fill_1 FILLER_54_975 ();
 sg13g2_fill_2 FILLER_54_1008 ();
 sg13g2_decap_8 FILLER_54_1054 ();
 sg13g2_decap_8 FILLER_54_1061 ();
 sg13g2_decap_8 FILLER_54_1068 ();
 sg13g2_decap_8 FILLER_54_1075 ();
 sg13g2_decap_8 FILLER_54_1082 ();
 sg13g2_decap_8 FILLER_54_1089 ();
 sg13g2_decap_4 FILLER_54_1096 ();
 sg13g2_fill_2 FILLER_54_1100 ();
 sg13g2_fill_1 FILLER_54_1184 ();
 sg13g2_decap_8 FILLER_54_1189 ();
 sg13g2_fill_2 FILLER_54_1196 ();
 sg13g2_fill_2 FILLER_54_1207 ();
 sg13g2_fill_1 FILLER_54_1209 ();
 sg13g2_decap_4 FILLER_54_1220 ();
 sg13g2_fill_1 FILLER_54_1224 ();
 sg13g2_decap_8 FILLER_54_1230 ();
 sg13g2_fill_1 FILLER_54_1237 ();
 sg13g2_fill_1 FILLER_54_1243 ();
 sg13g2_fill_2 FILLER_54_1248 ();
 sg13g2_fill_1 FILLER_54_1250 ();
 sg13g2_fill_1 FILLER_54_1261 ();
 sg13g2_fill_1 FILLER_54_1292 ();
 sg13g2_fill_2 FILLER_54_1298 ();
 sg13g2_fill_1 FILLER_54_1307 ();
 sg13g2_fill_1 FILLER_54_1315 ();
 sg13g2_fill_1 FILLER_54_1326 ();
 sg13g2_decap_8 FILLER_54_1373 ();
 sg13g2_decap_4 FILLER_54_1384 ();
 sg13g2_fill_1 FILLER_54_1388 ();
 sg13g2_decap_8 FILLER_54_1394 ();
 sg13g2_decap_8 FILLER_54_1401 ();
 sg13g2_decap_8 FILLER_54_1408 ();
 sg13g2_decap_8 FILLER_54_1415 ();
 sg13g2_decap_8 FILLER_54_1422 ();
 sg13g2_decap_4 FILLER_54_1429 ();
 sg13g2_fill_2 FILLER_54_1433 ();
 sg13g2_decap_8 FILLER_54_1493 ();
 sg13g2_decap_4 FILLER_54_1500 ();
 sg13g2_fill_1 FILLER_54_1504 ();
 sg13g2_fill_2 FILLER_54_1509 ();
 sg13g2_fill_1 FILLER_54_1511 ();
 sg13g2_fill_2 FILLER_54_1519 ();
 sg13g2_decap_8 FILLER_54_1547 ();
 sg13g2_decap_4 FILLER_54_1554 ();
 sg13g2_fill_2 FILLER_54_1558 ();
 sg13g2_decap_8 FILLER_54_1588 ();
 sg13g2_decap_8 FILLER_54_1595 ();
 sg13g2_fill_1 FILLER_54_1602 ();
 sg13g2_fill_1 FILLER_54_1612 ();
 sg13g2_decap_8 FILLER_54_1623 ();
 sg13g2_decap_4 FILLER_54_1630 ();
 sg13g2_fill_2 FILLER_54_1634 ();
 sg13g2_fill_2 FILLER_54_1639 ();
 sg13g2_fill_1 FILLER_54_1641 ();
 sg13g2_decap_4 FILLER_54_1668 ();
 sg13g2_fill_1 FILLER_54_1672 ();
 sg13g2_decap_4 FILLER_54_1681 ();
 sg13g2_fill_2 FILLER_54_1685 ();
 sg13g2_fill_1 FILLER_54_1705 ();
 sg13g2_decap_8 FILLER_54_1710 ();
 sg13g2_decap_4 FILLER_54_1717 ();
 sg13g2_fill_2 FILLER_54_1721 ();
 sg13g2_fill_2 FILLER_54_1727 ();
 sg13g2_fill_2 FILLER_54_1739 ();
 sg13g2_fill_2 FILLER_54_1778 ();
 sg13g2_fill_1 FILLER_54_1794 ();
 sg13g2_fill_2 FILLER_54_1803 ();
 sg13g2_fill_1 FILLER_54_1805 ();
 sg13g2_decap_8 FILLER_54_1819 ();
 sg13g2_fill_2 FILLER_54_1826 ();
 sg13g2_fill_1 FILLER_54_1828 ();
 sg13g2_fill_2 FILLER_54_1834 ();
 sg13g2_fill_1 FILLER_54_1836 ();
 sg13g2_fill_2 FILLER_54_1846 ();
 sg13g2_fill_1 FILLER_54_1863 ();
 sg13g2_fill_1 FILLER_54_1882 ();
 sg13g2_fill_2 FILLER_54_1888 ();
 sg13g2_fill_1 FILLER_54_1890 ();
 sg13g2_fill_1 FILLER_54_1896 ();
 sg13g2_fill_1 FILLER_54_1924 ();
 sg13g2_decap_8 FILLER_54_1930 ();
 sg13g2_decap_8 FILLER_54_1937 ();
 sg13g2_decap_4 FILLER_54_1944 ();
 sg13g2_fill_1 FILLER_54_1948 ();
 sg13g2_fill_2 FILLER_54_1963 ();
 sg13g2_decap_4 FILLER_54_1968 ();
 sg13g2_fill_1 FILLER_54_1978 ();
 sg13g2_fill_1 FILLER_54_2018 ();
 sg13g2_fill_2 FILLER_54_2026 ();
 sg13g2_fill_2 FILLER_54_2048 ();
 sg13g2_fill_2 FILLER_54_2059 ();
 sg13g2_fill_1 FILLER_54_2061 ();
 sg13g2_fill_2 FILLER_54_2066 ();
 sg13g2_decap_4 FILLER_54_2078 ();
 sg13g2_fill_2 FILLER_54_2082 ();
 sg13g2_decap_8 FILLER_54_2110 ();
 sg13g2_decap_8 FILLER_54_2121 ();
 sg13g2_decap_8 FILLER_54_2128 ();
 sg13g2_fill_2 FILLER_54_2138 ();
 sg13g2_fill_2 FILLER_54_2154 ();
 sg13g2_decap_4 FILLER_54_2192 ();
 sg13g2_fill_1 FILLER_54_2234 ();
 sg13g2_decap_8 FILLER_54_2248 ();
 sg13g2_decap_8 FILLER_54_2255 ();
 sg13g2_fill_1 FILLER_54_2262 ();
 sg13g2_fill_1 FILLER_54_2275 ();
 sg13g2_decap_4 FILLER_54_2300 ();
 sg13g2_decap_4 FILLER_54_2328 ();
 sg13g2_fill_2 FILLER_54_2345 ();
 sg13g2_decap_4 FILLER_54_2356 ();
 sg13g2_fill_2 FILLER_54_2360 ();
 sg13g2_decap_4 FILLER_54_2404 ();
 sg13g2_decap_4 FILLER_54_2434 ();
 sg13g2_fill_2 FILLER_54_2438 ();
 sg13g2_fill_1 FILLER_54_2462 ();
 sg13g2_fill_1 FILLER_54_2527 ();
 sg13g2_decap_4 FILLER_54_2558 ();
 sg13g2_fill_1 FILLER_54_2562 ();
 sg13g2_fill_1 FILLER_54_2586 ();
 sg13g2_decap_4 FILLER_54_2613 ();
 sg13g2_decap_8 FILLER_54_2621 ();
 sg13g2_decap_8 FILLER_54_2628 ();
 sg13g2_decap_8 FILLER_54_2635 ();
 sg13g2_decap_8 FILLER_54_2642 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_decap_8 FILLER_54_2656 ();
 sg13g2_decap_8 FILLER_54_2663 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_28 ();
 sg13g2_fill_1 FILLER_55_32 ();
 sg13g2_fill_1 FILLER_55_37 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_fill_2 FILLER_55_88 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_fill_1 FILLER_55_101 ();
 sg13g2_decap_4 FILLER_55_128 ();
 sg13g2_fill_2 FILLER_55_143 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_fill_1 FILLER_55_176 ();
 sg13g2_decap_4 FILLER_55_210 ();
 sg13g2_fill_2 FILLER_55_219 ();
 sg13g2_fill_1 FILLER_55_259 ();
 sg13g2_fill_2 FILLER_55_268 ();
 sg13g2_fill_1 FILLER_55_274 ();
 sg13g2_fill_1 FILLER_55_331 ();
 sg13g2_fill_1 FILLER_55_341 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_2 FILLER_55_389 ();
 sg13g2_fill_1 FILLER_55_391 ();
 sg13g2_fill_2 FILLER_55_405 ();
 sg13g2_fill_2 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_425 ();
 sg13g2_decap_4 FILLER_55_432 ();
 sg13g2_fill_1 FILLER_55_436 ();
 sg13g2_fill_2 FILLER_55_487 ();
 sg13g2_decap_4 FILLER_55_505 ();
 sg13g2_fill_2 FILLER_55_513 ();
 sg13g2_fill_1 FILLER_55_541 ();
 sg13g2_fill_1 FILLER_55_548 ();
 sg13g2_fill_1 FILLER_55_558 ();
 sg13g2_fill_1 FILLER_55_599 ();
 sg13g2_fill_1 FILLER_55_630 ();
 sg13g2_decap_4 FILLER_55_640 ();
 sg13g2_fill_2 FILLER_55_648 ();
 sg13g2_fill_2 FILLER_55_665 ();
 sg13g2_decap_4 FILLER_55_722 ();
 sg13g2_fill_1 FILLER_55_748 ();
 sg13g2_fill_2 FILLER_55_763 ();
 sg13g2_fill_2 FILLER_55_773 ();
 sg13g2_fill_1 FILLER_55_775 ();
 sg13g2_fill_2 FILLER_55_780 ();
 sg13g2_fill_1 FILLER_55_782 ();
 sg13g2_fill_2 FILLER_55_796 ();
 sg13g2_decap_8 FILLER_55_802 ();
 sg13g2_fill_2 FILLER_55_809 ();
 sg13g2_decap_4 FILLER_55_815 ();
 sg13g2_fill_2 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_887 ();
 sg13g2_fill_1 FILLER_55_894 ();
 sg13g2_decap_8 FILLER_55_917 ();
 sg13g2_fill_2 FILLER_55_924 ();
 sg13g2_decap_4 FILLER_55_962 ();
 sg13g2_fill_1 FILLER_55_966 ();
 sg13g2_decap_8 FILLER_55_1030 ();
 sg13g2_decap_8 FILLER_55_1037 ();
 sg13g2_decap_8 FILLER_55_1044 ();
 sg13g2_decap_8 FILLER_55_1051 ();
 sg13g2_decap_4 FILLER_55_1088 ();
 sg13g2_fill_2 FILLER_55_1118 ();
 sg13g2_fill_1 FILLER_55_1120 ();
 sg13g2_fill_1 FILLER_55_1151 ();
 sg13g2_fill_1 FILLER_55_1166 ();
 sg13g2_decap_4 FILLER_55_1170 ();
 sg13g2_fill_2 FILLER_55_1174 ();
 sg13g2_decap_8 FILLER_55_1182 ();
 sg13g2_fill_2 FILLER_55_1189 ();
 sg13g2_decap_4 FILLER_55_1252 ();
 sg13g2_fill_2 FILLER_55_1270 ();
 sg13g2_fill_1 FILLER_55_1300 ();
 sg13g2_fill_2 FILLER_55_1305 ();
 sg13g2_fill_1 FILLER_55_1312 ();
 sg13g2_decap_8 FILLER_55_1324 ();
 sg13g2_decap_8 FILLER_55_1331 ();
 sg13g2_fill_2 FILLER_55_1348 ();
 sg13g2_fill_1 FILLER_55_1350 ();
 sg13g2_decap_8 FILLER_55_1355 ();
 sg13g2_decap_4 FILLER_55_1362 ();
 sg13g2_fill_2 FILLER_55_1366 ();
 sg13g2_decap_8 FILLER_55_1377 ();
 sg13g2_decap_8 FILLER_55_1384 ();
 sg13g2_fill_1 FILLER_55_1404 ();
 sg13g2_fill_1 FILLER_55_1439 ();
 sg13g2_fill_1 FILLER_55_1445 ();
 sg13g2_fill_2 FILLER_55_1450 ();
 sg13g2_fill_1 FILLER_55_1464 ();
 sg13g2_decap_4 FILLER_55_1477 ();
 sg13g2_fill_1 FILLER_55_1481 ();
 sg13g2_decap_8 FILLER_55_1488 ();
 sg13g2_decap_4 FILLER_55_1495 ();
 sg13g2_fill_2 FILLER_55_1499 ();
 sg13g2_fill_2 FILLER_55_1537 ();
 sg13g2_fill_2 FILLER_55_1566 ();
 sg13g2_fill_1 FILLER_55_1568 ();
 sg13g2_fill_2 FILLER_55_1582 ();
 sg13g2_decap_4 FILLER_55_1601 ();
 sg13g2_fill_2 FILLER_55_1605 ();
 sg13g2_decap_4 FILLER_55_1611 ();
 sg13g2_fill_1 FILLER_55_1615 ();
 sg13g2_decap_8 FILLER_55_1620 ();
 sg13g2_decap_8 FILLER_55_1627 ();
 sg13g2_fill_2 FILLER_55_1634 ();
 sg13g2_fill_1 FILLER_55_1660 ();
 sg13g2_fill_1 FILLER_55_1667 ();
 sg13g2_fill_1 FILLER_55_1681 ();
 sg13g2_fill_1 FILLER_55_1687 ();
 sg13g2_fill_2 FILLER_55_1692 ();
 sg13g2_decap_4 FILLER_55_1724 ();
 sg13g2_decap_4 FILLER_55_1754 ();
 sg13g2_fill_1 FILLER_55_1758 ();
 sg13g2_fill_1 FILLER_55_1802 ();
 sg13g2_decap_8 FILLER_55_1813 ();
 sg13g2_decap_4 FILLER_55_1820 ();
 sg13g2_fill_2 FILLER_55_1828 ();
 sg13g2_fill_1 FILLER_55_1830 ();
 sg13g2_fill_2 FILLER_55_1842 ();
 sg13g2_fill_1 FILLER_55_1853 ();
 sg13g2_fill_1 FILLER_55_1879 ();
 sg13g2_fill_1 FILLER_55_1893 ();
 sg13g2_fill_2 FILLER_55_1925 ();
 sg13g2_fill_1 FILLER_55_1927 ();
 sg13g2_fill_2 FILLER_55_1932 ();
 sg13g2_decap_8 FILLER_55_1939 ();
 sg13g2_decap_4 FILLER_55_1946 ();
 sg13g2_fill_1 FILLER_55_1950 ();
 sg13g2_decap_8 FILLER_55_1955 ();
 sg13g2_decap_8 FILLER_55_1962 ();
 sg13g2_decap_8 FILLER_55_1969 ();
 sg13g2_decap_4 FILLER_55_1976 ();
 sg13g2_fill_1 FILLER_55_2031 ();
 sg13g2_fill_1 FILLER_55_2040 ();
 sg13g2_fill_2 FILLER_55_2056 ();
 sg13g2_fill_1 FILLER_55_2068 ();
 sg13g2_fill_1 FILLER_55_2091 ();
 sg13g2_fill_2 FILLER_55_2125 ();
 sg13g2_fill_2 FILLER_55_2185 ();
 sg13g2_fill_1 FILLER_55_2187 ();
 sg13g2_fill_2 FILLER_55_2204 ();
 sg13g2_fill_1 FILLER_55_2220 ();
 sg13g2_decap_8 FILLER_55_2236 ();
 sg13g2_fill_2 FILLER_55_2243 ();
 sg13g2_fill_2 FILLER_55_2256 ();
 sg13g2_fill_2 FILLER_55_2320 ();
 sg13g2_fill_2 FILLER_55_2338 ();
 sg13g2_decap_8 FILLER_55_2345 ();
 sg13g2_decap_8 FILLER_55_2352 ();
 sg13g2_fill_1 FILLER_55_2359 ();
 sg13g2_fill_1 FILLER_55_2376 ();
 sg13g2_fill_1 FILLER_55_2383 ();
 sg13g2_fill_1 FILLER_55_2389 ();
 sg13g2_fill_1 FILLER_55_2395 ();
 sg13g2_decap_8 FILLER_55_2400 ();
 sg13g2_decap_8 FILLER_55_2421 ();
 sg13g2_decap_8 FILLER_55_2428 ();
 sg13g2_fill_2 FILLER_55_2435 ();
 sg13g2_fill_1 FILLER_55_2437 ();
 sg13g2_fill_1 FILLER_55_2448 ();
 sg13g2_fill_1 FILLER_55_2475 ();
 sg13g2_fill_1 FILLER_55_2486 ();
 sg13g2_fill_1 FILLER_55_2491 ();
 sg13g2_fill_2 FILLER_55_2496 ();
 sg13g2_decap_4 FILLER_55_2503 ();
 sg13g2_fill_2 FILLER_55_2507 ();
 sg13g2_decap_8 FILLER_55_2513 ();
 sg13g2_fill_1 FILLER_55_2526 ();
 sg13g2_fill_2 FILLER_55_2541 ();
 sg13g2_fill_1 FILLER_55_2543 ();
 sg13g2_decap_8 FILLER_55_2640 ();
 sg13g2_decap_8 FILLER_55_2647 ();
 sg13g2_decap_8 FILLER_55_2654 ();
 sg13g2_decap_8 FILLER_55_2661 ();
 sg13g2_fill_2 FILLER_55_2668 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_fill_1 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_decap_4 FILLER_56_146 ();
 sg13g2_fill_2 FILLER_56_150 ();
 sg13g2_fill_2 FILLER_56_223 ();
 sg13g2_fill_1 FILLER_56_225 ();
 sg13g2_fill_2 FILLER_56_235 ();
 sg13g2_fill_2 FILLER_56_247 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_decap_8 FILLER_56_300 ();
 sg13g2_decap_4 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_325 ();
 sg13g2_decap_8 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_1 FILLER_56_359 ();
 sg13g2_decap_4 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_383 ();
 sg13g2_fill_2 FILLER_56_425 ();
 sg13g2_fill_1 FILLER_56_427 ();
 sg13g2_fill_2 FILLER_56_434 ();
 sg13g2_fill_1 FILLER_56_436 ();
 sg13g2_fill_2 FILLER_56_450 ();
 sg13g2_fill_2 FILLER_56_471 ();
 sg13g2_decap_8 FILLER_56_478 ();
 sg13g2_fill_1 FILLER_56_485 ();
 sg13g2_decap_8 FILLER_56_494 ();
 sg13g2_decap_4 FILLER_56_501 ();
 sg13g2_fill_1 FILLER_56_505 ();
 sg13g2_fill_1 FILLER_56_564 ();
 sg13g2_fill_1 FILLER_56_568 ();
 sg13g2_fill_1 FILLER_56_577 ();
 sg13g2_fill_1 FILLER_56_582 ();
 sg13g2_fill_2 FILLER_56_595 ();
 sg13g2_fill_1 FILLER_56_597 ();
 sg13g2_fill_2 FILLER_56_602 ();
 sg13g2_fill_2 FILLER_56_614 ();
 sg13g2_decap_4 FILLER_56_626 ();
 sg13g2_fill_2 FILLER_56_635 ();
 sg13g2_fill_2 FILLER_56_673 ();
 sg13g2_fill_1 FILLER_56_675 ();
 sg13g2_fill_1 FILLER_56_681 ();
 sg13g2_fill_1 FILLER_56_692 ();
 sg13g2_fill_2 FILLER_56_726 ();
 sg13g2_fill_1 FILLER_56_760 ();
 sg13g2_decap_8 FILLER_56_809 ();
 sg13g2_decap_8 FILLER_56_816 ();
 sg13g2_decap_4 FILLER_56_823 ();
 sg13g2_fill_2 FILLER_56_831 ();
 sg13g2_decap_4 FILLER_56_841 ();
 sg13g2_fill_1 FILLER_56_845 ();
 sg13g2_fill_2 FILLER_56_850 ();
 sg13g2_fill_1 FILLER_56_882 ();
 sg13g2_fill_2 FILLER_56_893 ();
 sg13g2_fill_1 FILLER_56_942 ();
 sg13g2_fill_2 FILLER_56_950 ();
 sg13g2_decap_8 FILLER_56_962 ();
 sg13g2_decap_4 FILLER_56_969 ();
 sg13g2_decap_8 FILLER_56_1040 ();
 sg13g2_fill_1 FILLER_56_1051 ();
 sg13g2_fill_2 FILLER_56_1056 ();
 sg13g2_fill_2 FILLER_56_1084 ();
 sg13g2_fill_2 FILLER_56_1096 ();
 sg13g2_fill_1 FILLER_56_1098 ();
 sg13g2_decap_4 FILLER_56_1103 ();
 sg13g2_fill_1 FILLER_56_1167 ();
 sg13g2_fill_1 FILLER_56_1175 ();
 sg13g2_decap_8 FILLER_56_1199 ();
 sg13g2_decap_8 FILLER_56_1206 ();
 sg13g2_decap_8 FILLER_56_1213 ();
 sg13g2_fill_1 FILLER_56_1220 ();
 sg13g2_decap_4 FILLER_56_1227 ();
 sg13g2_decap_8 FILLER_56_1239 ();
 sg13g2_decap_4 FILLER_56_1246 ();
 sg13g2_fill_1 FILLER_56_1250 ();
 sg13g2_fill_1 FILLER_56_1261 ();
 sg13g2_fill_1 FILLER_56_1272 ();
 sg13g2_fill_2 FILLER_56_1293 ();
 sg13g2_fill_1 FILLER_56_1302 ();
 sg13g2_decap_8 FILLER_56_1312 ();
 sg13g2_decap_8 FILLER_56_1319 ();
 sg13g2_decap_8 FILLER_56_1326 ();
 sg13g2_decap_8 FILLER_56_1333 ();
 sg13g2_fill_2 FILLER_56_1340 ();
 sg13g2_decap_4 FILLER_56_1368 ();
 sg13g2_decap_8 FILLER_56_1385 ();
 sg13g2_fill_1 FILLER_56_1392 ();
 sg13g2_fill_2 FILLER_56_1419 ();
 sg13g2_fill_1 FILLER_56_1421 ();
 sg13g2_decap_4 FILLER_56_1451 ();
 sg13g2_fill_2 FILLER_56_1455 ();
 sg13g2_fill_2 FILLER_56_1473 ();
 sg13g2_fill_1 FILLER_56_1475 ();
 sg13g2_fill_2 FILLER_56_1480 ();
 sg13g2_decap_4 FILLER_56_1487 ();
 sg13g2_fill_1 FILLER_56_1491 ();
 sg13g2_fill_2 FILLER_56_1530 ();
 sg13g2_fill_1 FILLER_56_1550 ();
 sg13g2_fill_1 FILLER_56_1556 ();
 sg13g2_fill_1 FILLER_56_1583 ();
 sg13g2_fill_2 FILLER_56_1617 ();
 sg13g2_decap_8 FILLER_56_1623 ();
 sg13g2_fill_2 FILLER_56_1630 ();
 sg13g2_fill_1 FILLER_56_1632 ();
 sg13g2_fill_1 FILLER_56_1643 ();
 sg13g2_fill_1 FILLER_56_1693 ();
 sg13g2_fill_2 FILLER_56_1703 ();
 sg13g2_fill_1 FILLER_56_1705 ();
 sg13g2_fill_1 FILLER_56_1715 ();
 sg13g2_decap_8 FILLER_56_1721 ();
 sg13g2_decap_8 FILLER_56_1728 ();
 sg13g2_decap_4 FILLER_56_1735 ();
 sg13g2_fill_1 FILLER_56_1739 ();
 sg13g2_fill_1 FILLER_56_1766 ();
 sg13g2_decap_4 FILLER_56_1818 ();
 sg13g2_fill_1 FILLER_56_1822 ();
 sg13g2_fill_1 FILLER_56_1828 ();
 sg13g2_fill_1 FILLER_56_1841 ();
 sg13g2_fill_1 FILLER_56_1870 ();
 sg13g2_fill_2 FILLER_56_1882 ();
 sg13g2_decap_4 FILLER_56_1930 ();
 sg13g2_fill_1 FILLER_56_1934 ();
 sg13g2_decap_8 FILLER_56_1940 ();
 sg13g2_fill_2 FILLER_56_1947 ();
 sg13g2_fill_2 FILLER_56_1954 ();
 sg13g2_fill_2 FILLER_56_1961 ();
 sg13g2_fill_1 FILLER_56_1963 ();
 sg13g2_fill_1 FILLER_56_1969 ();
 sg13g2_decap_4 FILLER_56_1975 ();
 sg13g2_fill_2 FILLER_56_1979 ();
 sg13g2_fill_2 FILLER_56_2019 ();
 sg13g2_fill_1 FILLER_56_2021 ();
 sg13g2_fill_1 FILLER_56_2026 ();
 sg13g2_fill_1 FILLER_56_2104 ();
 sg13g2_fill_1 FILLER_56_2142 ();
 sg13g2_fill_1 FILLER_56_2152 ();
 sg13g2_fill_2 FILLER_56_2209 ();
 sg13g2_fill_2 FILLER_56_2215 ();
 sg13g2_fill_1 FILLER_56_2217 ();
 sg13g2_fill_1 FILLER_56_2254 ();
 sg13g2_fill_1 FILLER_56_2263 ();
 sg13g2_fill_2 FILLER_56_2314 ();
 sg13g2_decap_4 FILLER_56_2327 ();
 sg13g2_fill_1 FILLER_56_2331 ();
 sg13g2_fill_2 FILLER_56_2335 ();
 sg13g2_fill_1 FILLER_56_2337 ();
 sg13g2_fill_1 FILLER_56_2343 ();
 sg13g2_fill_1 FILLER_56_2349 ();
 sg13g2_fill_1 FILLER_56_2354 ();
 sg13g2_fill_2 FILLER_56_2365 ();
 sg13g2_decap_8 FILLER_56_2393 ();
 sg13g2_decap_4 FILLER_56_2400 ();
 sg13g2_decap_8 FILLER_56_2484 ();
 sg13g2_decap_8 FILLER_56_2491 ();
 sg13g2_decap_4 FILLER_56_2502 ();
 sg13g2_fill_1 FILLER_56_2506 ();
 sg13g2_decap_4 FILLER_56_2511 ();
 sg13g2_fill_2 FILLER_56_2563 ();
 sg13g2_decap_8 FILLER_56_2642 ();
 sg13g2_decap_8 FILLER_56_2649 ();
 sg13g2_decap_8 FILLER_56_2656 ();
 sg13g2_decap_8 FILLER_56_2663 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_4 ();
 sg13g2_decap_4 FILLER_57_23 ();
 sg13g2_decap_8 FILLER_57_39 ();
 sg13g2_decap_8 FILLER_57_46 ();
 sg13g2_decap_8 FILLER_57_53 ();
 sg13g2_decap_4 FILLER_57_60 ();
 sg13g2_fill_1 FILLER_57_64 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_95 ();
 sg13g2_decap_4 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_132 ();
 sg13g2_decap_4 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_173 ();
 sg13g2_decap_4 FILLER_57_189 ();
 sg13g2_fill_1 FILLER_57_203 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_fill_2 FILLER_57_215 ();
 sg13g2_fill_1 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_276 ();
 sg13g2_fill_1 FILLER_57_289 ();
 sg13g2_fill_2 FILLER_57_294 ();
 sg13g2_fill_1 FILLER_57_296 ();
 sg13g2_fill_1 FILLER_57_370 ();
 sg13g2_fill_1 FILLER_57_376 ();
 sg13g2_fill_2 FILLER_57_400 ();
 sg13g2_decap_4 FILLER_57_432 ();
 sg13g2_fill_2 FILLER_57_436 ();
 sg13g2_decap_4 FILLER_57_447 ();
 sg13g2_fill_1 FILLER_57_451 ();
 sg13g2_fill_1 FILLER_57_457 ();
 sg13g2_fill_1 FILLER_57_463 ();
 sg13g2_fill_1 FILLER_57_469 ();
 sg13g2_fill_1 FILLER_57_474 ();
 sg13g2_fill_2 FILLER_57_479 ();
 sg13g2_decap_4 FILLER_57_485 ();
 sg13g2_fill_2 FILLER_57_503 ();
 sg13g2_decap_8 FILLER_57_509 ();
 sg13g2_decap_4 FILLER_57_516 ();
 sg13g2_fill_1 FILLER_57_520 ();
 sg13g2_fill_1 FILLER_57_555 ();
 sg13g2_decap_4 FILLER_57_595 ();
 sg13g2_fill_2 FILLER_57_599 ();
 sg13g2_decap_8 FILLER_57_619 ();
 sg13g2_decap_8 FILLER_57_626 ();
 sg13g2_fill_1 FILLER_57_633 ();
 sg13g2_decap_8 FILLER_57_664 ();
 sg13g2_decap_8 FILLER_57_671 ();
 sg13g2_fill_1 FILLER_57_678 ();
 sg13g2_decap_4 FILLER_57_739 ();
 sg13g2_fill_2 FILLER_57_743 ();
 sg13g2_fill_2 FILLER_57_750 ();
 sg13g2_fill_1 FILLER_57_802 ();
 sg13g2_decap_8 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_826 ();
 sg13g2_decap_8 FILLER_57_833 ();
 sg13g2_decap_8 FILLER_57_840 ();
 sg13g2_fill_1 FILLER_57_847 ();
 sg13g2_decap_8 FILLER_57_888 ();
 sg13g2_decap_8 FILLER_57_895 ();
 sg13g2_decap_8 FILLER_57_902 ();
 sg13g2_fill_2 FILLER_57_909 ();
 sg13g2_fill_1 FILLER_57_911 ();
 sg13g2_fill_1 FILLER_57_955 ();
 sg13g2_fill_1 FILLER_57_1005 ();
 sg13g2_decap_4 FILLER_57_1010 ();
 sg13g2_fill_1 FILLER_57_1029 ();
 sg13g2_decap_4 FILLER_57_1066 ();
 sg13g2_fill_1 FILLER_57_1070 ();
 sg13g2_fill_2 FILLER_57_1104 ();
 sg13g2_fill_1 FILLER_57_1106 ();
 sg13g2_fill_2 FILLER_57_1115 ();
 sg13g2_decap_4 FILLER_57_1131 ();
 sg13g2_fill_2 FILLER_57_1187 ();
 sg13g2_decap_8 FILLER_57_1199 ();
 sg13g2_decap_8 FILLER_57_1206 ();
 sg13g2_fill_2 FILLER_57_1213 ();
 sg13g2_fill_1 FILLER_57_1215 ();
 sg13g2_decap_8 FILLER_57_1245 ();
 sg13g2_fill_2 FILLER_57_1252 ();
 sg13g2_decap_8 FILLER_57_1259 ();
 sg13g2_fill_2 FILLER_57_1266 ();
 sg13g2_fill_2 FILLER_57_1273 ();
 sg13g2_fill_2 FILLER_57_1278 ();
 sg13g2_fill_1 FILLER_57_1280 ();
 sg13g2_fill_2 FILLER_57_1288 ();
 sg13g2_fill_1 FILLER_57_1290 ();
 sg13g2_fill_2 FILLER_57_1296 ();
 sg13g2_decap_4 FILLER_57_1302 ();
 sg13g2_decap_4 FILLER_57_1334 ();
 sg13g2_decap_4 FILLER_57_1342 ();
 sg13g2_fill_1 FILLER_57_1346 ();
 sg13g2_decap_8 FILLER_57_1351 ();
 sg13g2_fill_2 FILLER_57_1358 ();
 sg13g2_decap_4 FILLER_57_1368 ();
 sg13g2_decap_8 FILLER_57_1387 ();
 sg13g2_decap_4 FILLER_57_1394 ();
 sg13g2_fill_2 FILLER_57_1398 ();
 sg13g2_fill_2 FILLER_57_1410 ();
 sg13g2_fill_2 FILLER_57_1417 ();
 sg13g2_decap_8 FILLER_57_1449 ();
 sg13g2_fill_1 FILLER_57_1482 ();
 sg13g2_fill_1 FILLER_57_1492 ();
 sg13g2_fill_2 FILLER_57_1501 ();
 sg13g2_fill_2 FILLER_57_1520 ();
 sg13g2_fill_1 FILLER_57_1532 ();
 sg13g2_fill_1 FILLER_57_1537 ();
 sg13g2_fill_2 FILLER_57_1584 ();
 sg13g2_fill_1 FILLER_57_1586 ();
 sg13g2_fill_1 FILLER_57_1597 ();
 sg13g2_fill_1 FILLER_57_1615 ();
 sg13g2_fill_1 FILLER_57_1625 ();
 sg13g2_decap_8 FILLER_57_1633 ();
 sg13g2_fill_2 FILLER_57_1640 ();
 sg13g2_fill_1 FILLER_57_1651 ();
 sg13g2_fill_1 FILLER_57_1662 ();
 sg13g2_fill_1 FILLER_57_1668 ();
 sg13g2_fill_1 FILLER_57_1677 ();
 sg13g2_fill_1 FILLER_57_1682 ();
 sg13g2_fill_1 FILLER_57_1698 ();
 sg13g2_decap_8 FILLER_57_1718 ();
 sg13g2_decap_8 FILLER_57_1725 ();
 sg13g2_decap_8 FILLER_57_1732 ();
 sg13g2_fill_2 FILLER_57_1739 ();
 sg13g2_fill_1 FILLER_57_1741 ();
 sg13g2_decap_4 FILLER_57_1746 ();
 sg13g2_fill_1 FILLER_57_1768 ();
 sg13g2_fill_2 FILLER_57_1782 ();
 sg13g2_fill_1 FILLER_57_1796 ();
 sg13g2_decap_8 FILLER_57_1805 ();
 sg13g2_decap_8 FILLER_57_1817 ();
 sg13g2_decap_4 FILLER_57_1828 ();
 sg13g2_fill_1 FILLER_57_1832 ();
 sg13g2_fill_1 FILLER_57_1875 ();
 sg13g2_fill_1 FILLER_57_1884 ();
 sg13g2_fill_2 FILLER_57_1890 ();
 sg13g2_fill_2 FILLER_57_1910 ();
 sg13g2_fill_1 FILLER_57_1917 ();
 sg13g2_decap_8 FILLER_57_1927 ();
 sg13g2_decap_8 FILLER_57_1934 ();
 sg13g2_fill_2 FILLER_57_1941 ();
 sg13g2_fill_1 FILLER_57_1943 ();
 sg13g2_fill_1 FILLER_57_1966 ();
 sg13g2_decap_4 FILLER_57_1972 ();
 sg13g2_fill_1 FILLER_57_1976 ();
 sg13g2_fill_2 FILLER_57_1982 ();
 sg13g2_fill_1 FILLER_57_1984 ();
 sg13g2_fill_1 FILLER_57_1994 ();
 sg13g2_fill_2 FILLER_57_2000 ();
 sg13g2_decap_8 FILLER_57_2011 ();
 sg13g2_fill_1 FILLER_57_2018 ();
 sg13g2_decap_4 FILLER_57_2032 ();
 sg13g2_fill_1 FILLER_57_2036 ();
 sg13g2_decap_4 FILLER_57_2049 ();
 sg13g2_fill_1 FILLER_57_2057 ();
 sg13g2_fill_2 FILLER_57_2067 ();
 sg13g2_fill_2 FILLER_57_2084 ();
 sg13g2_fill_1 FILLER_57_2094 ();
 sg13g2_fill_1 FILLER_57_2099 ();
 sg13g2_decap_8 FILLER_57_2104 ();
 sg13g2_decap_4 FILLER_57_2111 ();
 sg13g2_fill_1 FILLER_57_2115 ();
 sg13g2_decap_8 FILLER_57_2144 ();
 sg13g2_fill_2 FILLER_57_2151 ();
 sg13g2_decap_8 FILLER_57_2163 ();
 sg13g2_fill_2 FILLER_57_2175 ();
 sg13g2_fill_1 FILLER_57_2177 ();
 sg13g2_fill_1 FILLER_57_2196 ();
 sg13g2_fill_1 FILLER_57_2208 ();
 sg13g2_fill_1 FILLER_57_2213 ();
 sg13g2_fill_2 FILLER_57_2218 ();
 sg13g2_fill_1 FILLER_57_2225 ();
 sg13g2_fill_1 FILLER_57_2236 ();
 sg13g2_fill_1 FILLER_57_2273 ();
 sg13g2_fill_2 FILLER_57_2293 ();
 sg13g2_fill_1 FILLER_57_2295 ();
 sg13g2_fill_1 FILLER_57_2328 ();
 sg13g2_fill_1 FILLER_57_2359 ();
 sg13g2_fill_2 FILLER_57_2366 ();
 sg13g2_fill_2 FILLER_57_2372 ();
 sg13g2_fill_2 FILLER_57_2413 ();
 sg13g2_fill_1 FILLER_57_2441 ();
 sg13g2_fill_2 FILLER_57_2452 ();
 sg13g2_fill_1 FILLER_57_2480 ();
 sg13g2_fill_2 FILLER_57_2485 ();
 sg13g2_decap_8 FILLER_57_2548 ();
 sg13g2_fill_1 FILLER_57_2555 ();
 sg13g2_fill_1 FILLER_57_2587 ();
 sg13g2_decap_4 FILLER_57_2616 ();
 sg13g2_fill_1 FILLER_57_2620 ();
 sg13g2_decap_8 FILLER_57_2651 ();
 sg13g2_decap_8 FILLER_57_2658 ();
 sg13g2_decap_4 FILLER_57_2665 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_22 ();
 sg13g2_fill_1 FILLER_58_33 ();
 sg13g2_decap_8 FILLER_58_51 ();
 sg13g2_decap_8 FILLER_58_58 ();
 sg13g2_decap_8 FILLER_58_65 ();
 sg13g2_decap_8 FILLER_58_72 ();
 sg13g2_decap_8 FILLER_58_79 ();
 sg13g2_fill_2 FILLER_58_86 ();
 sg13g2_decap_4 FILLER_58_92 ();
 sg13g2_fill_1 FILLER_58_96 ();
 sg13g2_fill_2 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_149 ();
 sg13g2_fill_2 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_fill_2 FILLER_58_206 ();
 sg13g2_fill_1 FILLER_58_213 ();
 sg13g2_decap_8 FILLER_58_219 ();
 sg13g2_decap_4 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_267 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_fill_2 FILLER_58_308 ();
 sg13g2_fill_1 FILLER_58_310 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_fill_2 FILLER_58_326 ();
 sg13g2_fill_1 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_338 ();
 sg13g2_fill_1 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_381 ();
 sg13g2_fill_1 FILLER_58_414 ();
 sg13g2_fill_2 FILLER_58_421 ();
 sg13g2_decap_8 FILLER_58_427 ();
 sg13g2_fill_2 FILLER_58_434 ();
 sg13g2_fill_2 FILLER_58_467 ();
 sg13g2_fill_1 FILLER_58_469 ();
 sg13g2_fill_2 FILLER_58_506 ();
 sg13g2_fill_1 FILLER_58_508 ();
 sg13g2_decap_8 FILLER_58_514 ();
 sg13g2_fill_1 FILLER_58_524 ();
 sg13g2_fill_2 FILLER_58_530 ();
 sg13g2_fill_1 FILLER_58_548 ();
 sg13g2_fill_2 FILLER_58_604 ();
 sg13g2_fill_1 FILLER_58_606 ();
 sg13g2_fill_1 FILLER_58_619 ();
 sg13g2_fill_1 FILLER_58_630 ();
 sg13g2_fill_1 FILLER_58_647 ();
 sg13g2_fill_1 FILLER_58_660 ();
 sg13g2_decap_4 FILLER_58_675 ();
 sg13g2_fill_2 FILLER_58_679 ();
 sg13g2_fill_1 FILLER_58_704 ();
 sg13g2_fill_1 FILLER_58_724 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_fill_2 FILLER_58_748 ();
 sg13g2_fill_1 FILLER_58_750 ();
 sg13g2_fill_2 FILLER_58_755 ();
 sg13g2_fill_2 FILLER_58_801 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_4 FILLER_58_849 ();
 sg13g2_fill_1 FILLER_58_853 ();
 sg13g2_fill_1 FILLER_58_869 ();
 sg13g2_decap_8 FILLER_58_896 ();
 sg13g2_decap_8 FILLER_58_903 ();
 sg13g2_fill_2 FILLER_58_910 ();
 sg13g2_fill_1 FILLER_58_912 ();
 sg13g2_fill_2 FILLER_58_918 ();
 sg13g2_fill_2 FILLER_58_950 ();
 sg13g2_fill_2 FILLER_58_968 ();
 sg13g2_fill_2 FILLER_58_979 ();
 sg13g2_fill_1 FILLER_58_981 ();
 sg13g2_fill_1 FILLER_58_1015 ();
 sg13g2_fill_1 FILLER_58_1022 ();
 sg13g2_decap_8 FILLER_58_1055 ();
 sg13g2_decap_8 FILLER_58_1062 ();
 sg13g2_decap_8 FILLER_58_1069 ();
 sg13g2_decap_4 FILLER_58_1076 ();
 sg13g2_fill_2 FILLER_58_1080 ();
 sg13g2_fill_2 FILLER_58_1099 ();
 sg13g2_decap_8 FILLER_58_1127 ();
 sg13g2_decap_8 FILLER_58_1134 ();
 sg13g2_fill_1 FILLER_58_1141 ();
 sg13g2_decap_4 FILLER_58_1176 ();
 sg13g2_fill_2 FILLER_58_1180 ();
 sg13g2_decap_4 FILLER_58_1185 ();
 sg13g2_decap_4 FILLER_58_1195 ();
 sg13g2_fill_1 FILLER_58_1199 ();
 sg13g2_decap_4 FILLER_58_1204 ();
 sg13g2_fill_1 FILLER_58_1208 ();
 sg13g2_decap_8 FILLER_58_1239 ();
 sg13g2_decap_4 FILLER_58_1246 ();
 sg13g2_fill_1 FILLER_58_1250 ();
 sg13g2_decap_4 FILLER_58_1255 ();
 sg13g2_fill_2 FILLER_58_1275 ();
 sg13g2_fill_1 FILLER_58_1287 ();
 sg13g2_decap_4 FILLER_58_1294 ();
 sg13g2_fill_2 FILLER_58_1298 ();
 sg13g2_fill_1 FILLER_58_1307 ();
 sg13g2_fill_2 FILLER_58_1317 ();
 sg13g2_fill_1 FILLER_58_1319 ();
 sg13g2_fill_1 FILLER_58_1329 ();
 sg13g2_fill_2 FILLER_58_1345 ();
 sg13g2_fill_1 FILLER_58_1347 ();
 sg13g2_fill_1 FILLER_58_1352 ();
 sg13g2_decap_8 FILLER_58_1366 ();
 sg13g2_decap_4 FILLER_58_1373 ();
 sg13g2_fill_2 FILLER_58_1377 ();
 sg13g2_fill_2 FILLER_58_1384 ();
 sg13g2_fill_1 FILLER_58_1386 ();
 sg13g2_fill_2 FILLER_58_1396 ();
 sg13g2_decap_8 FILLER_58_1411 ();
 sg13g2_fill_2 FILLER_58_1428 ();
 sg13g2_fill_1 FILLER_58_1430 ();
 sg13g2_fill_1 FILLER_58_1439 ();
 sg13g2_decap_8 FILLER_58_1450 ();
 sg13g2_decap_4 FILLER_58_1457 ();
 sg13g2_fill_2 FILLER_58_1465 ();
 sg13g2_fill_2 FILLER_58_1471 ();
 sg13g2_fill_1 FILLER_58_1473 ();
 sg13g2_fill_1 FILLER_58_1505 ();
 sg13g2_fill_1 FILLER_58_1512 ();
 sg13g2_fill_1 FILLER_58_1536 ();
 sg13g2_fill_1 FILLER_58_1542 ();
 sg13g2_fill_1 FILLER_58_1547 ();
 sg13g2_decap_4 FILLER_58_1580 ();
 sg13g2_fill_2 FILLER_58_1594 ();
 sg13g2_fill_1 FILLER_58_1596 ();
 sg13g2_decap_8 FILLER_58_1602 ();
 sg13g2_fill_2 FILLER_58_1609 ();
 sg13g2_decap_4 FILLER_58_1614 ();
 sg13g2_fill_2 FILLER_58_1618 ();
 sg13g2_fill_1 FILLER_58_1625 ();
 sg13g2_decap_8 FILLER_58_1630 ();
 sg13g2_fill_1 FILLER_58_1637 ();
 sg13g2_decap_8 FILLER_58_1642 ();
 sg13g2_fill_2 FILLER_58_1649 ();
 sg13g2_fill_2 FILLER_58_1655 ();
 sg13g2_decap_4 FILLER_58_1666 ();
 sg13g2_fill_1 FILLER_58_1675 ();
 sg13g2_fill_1 FILLER_58_1699 ();
 sg13g2_decap_4 FILLER_58_1705 ();
 sg13g2_decap_8 FILLER_58_1740 ();
 sg13g2_fill_2 FILLER_58_1747 ();
 sg13g2_decap_8 FILLER_58_1757 ();
 sg13g2_decap_4 FILLER_58_1764 ();
 sg13g2_fill_2 FILLER_58_1768 ();
 sg13g2_decap_4 FILLER_58_1803 ();
 sg13g2_decap_8 FILLER_58_1824 ();
 sg13g2_fill_1 FILLER_58_1831 ();
 sg13g2_fill_1 FILLER_58_1836 ();
 sg13g2_fill_1 FILLER_58_1842 ();
 sg13g2_fill_2 FILLER_58_1882 ();
 sg13g2_fill_1 FILLER_58_1901 ();
 sg13g2_fill_1 FILLER_58_1908 ();
 sg13g2_fill_1 FILLER_58_1917 ();
 sg13g2_decap_8 FILLER_58_1922 ();
 sg13g2_decap_8 FILLER_58_1929 ();
 sg13g2_decap_8 FILLER_58_1936 ();
 sg13g2_decap_8 FILLER_58_1943 ();
 sg13g2_fill_1 FILLER_58_1950 ();
 sg13g2_fill_2 FILLER_58_2012 ();
 sg13g2_fill_1 FILLER_58_2046 ();
 sg13g2_decap_4 FILLER_58_2058 ();
 sg13g2_decap_8 FILLER_58_2095 ();
 sg13g2_fill_2 FILLER_58_2140 ();
 sg13g2_fill_1 FILLER_58_2142 ();
 sg13g2_fill_2 FILLER_58_2153 ();
 sg13g2_fill_1 FILLER_58_2155 ();
 sg13g2_fill_2 FILLER_58_2200 ();
 sg13g2_fill_2 FILLER_58_2212 ();
 sg13g2_fill_1 FILLER_58_2214 ();
 sg13g2_fill_1 FILLER_58_2220 ();
 sg13g2_fill_2 FILLER_58_2226 ();
 sg13g2_fill_1 FILLER_58_2254 ();
 sg13g2_fill_1 FILLER_58_2259 ();
 sg13g2_fill_1 FILLER_58_2270 ();
 sg13g2_decap_8 FILLER_58_2281 ();
 sg13g2_fill_1 FILLER_58_2288 ();
 sg13g2_fill_2 FILLER_58_2299 ();
 sg13g2_decap_4 FILLER_58_2357 ();
 sg13g2_fill_2 FILLER_58_2367 ();
 sg13g2_fill_1 FILLER_58_2369 ();
 sg13g2_fill_2 FILLER_58_2541 ();
 sg13g2_decap_4 FILLER_58_2553 ();
 sg13g2_fill_1 FILLER_58_2557 ();
 sg13g2_fill_2 FILLER_58_2593 ();
 sg13g2_fill_1 FILLER_58_2595 ();
 sg13g2_decap_4 FILLER_58_2626 ();
 sg13g2_fill_1 FILLER_58_2630 ();
 sg13g2_decap_8 FILLER_58_2657 ();
 sg13g2_decap_4 FILLER_58_2664 ();
 sg13g2_fill_2 FILLER_58_2668 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_16 ();
 sg13g2_fill_1 FILLER_59_21 ();
 sg13g2_fill_1 FILLER_59_31 ();
 sg13g2_fill_2 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_61 ();
 sg13g2_decap_8 FILLER_59_68 ();
 sg13g2_decap_8 FILLER_59_75 ();
 sg13g2_fill_2 FILLER_59_87 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_decap_4 FILLER_59_238 ();
 sg13g2_fill_2 FILLER_59_249 ();
 sg13g2_fill_1 FILLER_59_251 ();
 sg13g2_fill_2 FILLER_59_272 ();
 sg13g2_fill_1 FILLER_59_274 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_fill_2 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_342 ();
 sg13g2_fill_2 FILLER_59_349 ();
 sg13g2_fill_2 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_376 ();
 sg13g2_decap_8 FILLER_59_383 ();
 sg13g2_fill_2 FILLER_59_390 ();
 sg13g2_decap_8 FILLER_59_396 ();
 sg13g2_fill_1 FILLER_59_403 ();
 sg13g2_decap_4 FILLER_59_414 ();
 sg13g2_fill_1 FILLER_59_418 ();
 sg13g2_fill_2 FILLER_59_454 ();
 sg13g2_fill_1 FILLER_59_456 ();
 sg13g2_fill_2 FILLER_59_500 ();
 sg13g2_fill_2 FILLER_59_539 ();
 sg13g2_fill_2 FILLER_59_595 ();
 sg13g2_fill_2 FILLER_59_623 ();
 sg13g2_fill_2 FILLER_59_630 ();
 sg13g2_decap_4 FILLER_59_642 ();
 sg13g2_fill_2 FILLER_59_646 ();
 sg13g2_decap_8 FILLER_59_653 ();
 sg13g2_decap_4 FILLER_59_660 ();
 sg13g2_fill_2 FILLER_59_664 ();
 sg13g2_fill_1 FILLER_59_691 ();
 sg13g2_fill_2 FILLER_59_708 ();
 sg13g2_fill_1 FILLER_59_710 ();
 sg13g2_decap_4 FILLER_59_715 ();
 sg13g2_fill_1 FILLER_59_742 ();
 sg13g2_fill_2 FILLER_59_749 ();
 sg13g2_fill_1 FILLER_59_780 ();
 sg13g2_fill_2 FILLER_59_785 ();
 sg13g2_decap_4 FILLER_59_800 ();
 sg13g2_decap_4 FILLER_59_809 ();
 sg13g2_decap_4 FILLER_59_817 ();
 sg13g2_fill_2 FILLER_59_821 ();
 sg13g2_decap_4 FILLER_59_827 ();
 sg13g2_fill_2 FILLER_59_831 ();
 sg13g2_fill_2 FILLER_59_928 ();
 sg13g2_fill_2 FILLER_59_934 ();
 sg13g2_fill_1 FILLER_59_936 ();
 sg13g2_fill_1 FILLER_59_966 ();
 sg13g2_fill_1 FILLER_59_1002 ();
 sg13g2_fill_1 FILLER_59_1029 ();
 sg13g2_decap_8 FILLER_59_1069 ();
 sg13g2_decap_4 FILLER_59_1076 ();
 sg13g2_fill_1 FILLER_59_1080 ();
 sg13g2_fill_1 FILLER_59_1107 ();
 sg13g2_fill_1 FILLER_59_1116 ();
 sg13g2_fill_1 FILLER_59_1127 ();
 sg13g2_decap_4 FILLER_59_1132 ();
 sg13g2_fill_2 FILLER_59_1136 ();
 sg13g2_decap_4 FILLER_59_1148 ();
 sg13g2_fill_2 FILLER_59_1152 ();
 sg13g2_decap_4 FILLER_59_1164 ();
 sg13g2_fill_1 FILLER_59_1168 ();
 sg13g2_decap_4 FILLER_59_1173 ();
 sg13g2_fill_1 FILLER_59_1177 ();
 sg13g2_fill_1 FILLER_59_1204 ();
 sg13g2_fill_1 FILLER_59_1215 ();
 sg13g2_fill_1 FILLER_59_1220 ();
 sg13g2_fill_1 FILLER_59_1235 ();
 sg13g2_fill_2 FILLER_59_1241 ();
 sg13g2_fill_1 FILLER_59_1247 ();
 sg13g2_fill_1 FILLER_59_1263 ();
 sg13g2_fill_1 FILLER_59_1290 ();
 sg13g2_fill_2 FILLER_59_1297 ();
 sg13g2_fill_1 FILLER_59_1303 ();
 sg13g2_fill_2 FILLER_59_1310 ();
 sg13g2_fill_1 FILLER_59_1327 ();
 sg13g2_decap_4 FILLER_59_1337 ();
 sg13g2_decap_8 FILLER_59_1351 ();
 sg13g2_fill_1 FILLER_59_1358 ();
 sg13g2_fill_1 FILLER_59_1381 ();
 sg13g2_fill_2 FILLER_59_1386 ();
 sg13g2_fill_2 FILLER_59_1393 ();
 sg13g2_fill_1 FILLER_59_1395 ();
 sg13g2_fill_2 FILLER_59_1409 ();
 sg13g2_fill_1 FILLER_59_1411 ();
 sg13g2_decap_4 FILLER_59_1416 ();
 sg13g2_fill_2 FILLER_59_1420 ();
 sg13g2_decap_4 FILLER_59_1427 ();
 sg13g2_fill_2 FILLER_59_1431 ();
 sg13g2_fill_2 FILLER_59_1438 ();
 sg13g2_decap_4 FILLER_59_1470 ();
 sg13g2_fill_2 FILLER_59_1474 ();
 sg13g2_fill_1 FILLER_59_1498 ();
 sg13g2_decap_4 FILLER_59_1533 ();
 sg13g2_fill_1 FILLER_59_1559 ();
 sg13g2_fill_1 FILLER_59_1569 ();
 sg13g2_fill_2 FILLER_59_1591 ();
 sg13g2_fill_2 FILLER_59_1601 ();
 sg13g2_fill_1 FILLER_59_1607 ();
 sg13g2_decap_8 FILLER_59_1612 ();
 sg13g2_fill_2 FILLER_59_1619 ();
 sg13g2_fill_1 FILLER_59_1641 ();
 sg13g2_fill_2 FILLER_59_1650 ();
 sg13g2_fill_2 FILLER_59_1675 ();
 sg13g2_fill_1 FILLER_59_1715 ();
 sg13g2_fill_1 FILLER_59_1724 ();
 sg13g2_decap_8 FILLER_59_1729 ();
 sg13g2_decap_8 FILLER_59_1736 ();
 sg13g2_decap_4 FILLER_59_1743 ();
 sg13g2_fill_2 FILLER_59_1752 ();
 sg13g2_fill_1 FILLER_59_1754 ();
 sg13g2_decap_8 FILLER_59_1763 ();
 sg13g2_decap_8 FILLER_59_1770 ();
 sg13g2_fill_1 FILLER_59_1777 ();
 sg13g2_fill_1 FILLER_59_1799 ();
 sg13g2_fill_2 FILLER_59_1809 ();
 sg13g2_fill_1 FILLER_59_1811 ();
 sg13g2_decap_8 FILLER_59_1822 ();
 sg13g2_fill_2 FILLER_59_1834 ();
 sg13g2_fill_2 FILLER_59_1897 ();
 sg13g2_decap_8 FILLER_59_1918 ();
 sg13g2_decap_8 FILLER_59_1925 ();
 sg13g2_decap_8 FILLER_59_1932 ();
 sg13g2_decap_8 FILLER_59_1939 ();
 sg13g2_decap_8 FILLER_59_1946 ();
 sg13g2_fill_2 FILLER_59_1953 ();
 sg13g2_fill_1 FILLER_59_1955 ();
 sg13g2_fill_1 FILLER_59_1964 ();
 sg13g2_decap_4 FILLER_59_1970 ();
 sg13g2_fill_2 FILLER_59_1974 ();
 sg13g2_decap_8 FILLER_59_1980 ();
 sg13g2_fill_1 FILLER_59_2021 ();
 sg13g2_fill_1 FILLER_59_2052 ();
 sg13g2_fill_1 FILLER_59_2057 ();
 sg13g2_fill_1 FILLER_59_2068 ();
 sg13g2_fill_1 FILLER_59_2083 ();
 sg13g2_fill_2 FILLER_59_2087 ();
 sg13g2_decap_8 FILLER_59_2093 ();
 sg13g2_decap_8 FILLER_59_2100 ();
 sg13g2_fill_1 FILLER_59_2107 ();
 sg13g2_fill_1 FILLER_59_2118 ();
 sg13g2_fill_2 FILLER_59_2162 ();
 sg13g2_decap_4 FILLER_59_2172 ();
 sg13g2_fill_2 FILLER_59_2176 ();
 sg13g2_fill_1 FILLER_59_2212 ();
 sg13g2_fill_2 FILLER_59_2227 ();
 sg13g2_fill_1 FILLER_59_2239 ();
 sg13g2_fill_1 FILLER_59_2266 ();
 sg13g2_decap_8 FILLER_59_2293 ();
 sg13g2_fill_2 FILLER_59_2314 ();
 sg13g2_fill_1 FILLER_59_2316 ();
 sg13g2_decap_4 FILLER_59_2321 ();
 sg13g2_fill_2 FILLER_59_2348 ();
 sg13g2_decap_4 FILLER_59_2360 ();
 sg13g2_fill_1 FILLER_59_2364 ();
 sg13g2_fill_1 FILLER_59_2371 ();
 sg13g2_decap_8 FILLER_59_2462 ();
 sg13g2_decap_8 FILLER_59_2469 ();
 sg13g2_fill_2 FILLER_59_2476 ();
 sg13g2_decap_4 FILLER_59_2486 ();
 sg13g2_fill_2 FILLER_59_2490 ();
 sg13g2_fill_2 FILLER_59_2496 ();
 sg13g2_decap_8 FILLER_59_2502 ();
 sg13g2_fill_2 FILLER_59_2509 ();
 sg13g2_fill_1 FILLER_59_2515 ();
 sg13g2_fill_2 FILLER_59_2520 ();
 sg13g2_fill_1 FILLER_59_2522 ();
 sg13g2_decap_8 FILLER_59_2555 ();
 sg13g2_fill_2 FILLER_59_2562 ();
 sg13g2_fill_2 FILLER_59_2632 ();
 sg13g2_fill_1 FILLER_59_2634 ();
 sg13g2_decap_8 FILLER_59_2639 ();
 sg13g2_decap_8 FILLER_59_2646 ();
 sg13g2_decap_8 FILLER_59_2653 ();
 sg13g2_decap_8 FILLER_59_2660 ();
 sg13g2_fill_2 FILLER_59_2667 ();
 sg13g2_fill_1 FILLER_59_2669 ();
 sg13g2_fill_1 FILLER_60_19 ();
 sg13g2_fill_2 FILLER_60_37 ();
 sg13g2_fill_1 FILLER_60_62 ();
 sg13g2_fill_1 FILLER_60_94 ();
 sg13g2_decap_4 FILLER_60_129 ();
 sg13g2_fill_1 FILLER_60_133 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_160 ();
 sg13g2_decap_8 FILLER_60_171 ();
 sg13g2_fill_2 FILLER_60_178 ();
 sg13g2_fill_2 FILLER_60_211 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_decap_4 FILLER_60_230 ();
 sg13g2_fill_2 FILLER_60_234 ();
 sg13g2_fill_1 FILLER_60_240 ();
 sg13g2_fill_1 FILLER_60_245 ();
 sg13g2_fill_2 FILLER_60_251 ();
 sg13g2_fill_1 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_263 ();
 sg13g2_decap_4 FILLER_60_304 ();
 sg13g2_decap_8 FILLER_60_344 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_fill_2 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_373 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_4 FILLER_60_398 ();
 sg13g2_fill_1 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_60_419 ();
 sg13g2_decap_8 FILLER_60_426 ();
 sg13g2_fill_1 FILLER_60_433 ();
 sg13g2_fill_1 FILLER_60_468 ();
 sg13g2_fill_1 FILLER_60_510 ();
 sg13g2_fill_2 FILLER_60_515 ();
 sg13g2_fill_2 FILLER_60_570 ();
 sg13g2_fill_1 FILLER_60_609 ();
 sg13g2_fill_1 FILLER_60_614 ();
 sg13g2_fill_2 FILLER_60_627 ();
 sg13g2_decap_8 FILLER_60_659 ();
 sg13g2_decap_8 FILLER_60_666 ();
 sg13g2_fill_1 FILLER_60_673 ();
 sg13g2_decap_8 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_4 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_8 FILLER_60_812 ();
 sg13g2_decap_8 FILLER_60_819 ();
 sg13g2_fill_2 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_fill_1 FILLER_60_851 ();
 sg13g2_fill_2 FILLER_60_891 ();
 sg13g2_fill_1 FILLER_60_908 ();
 sg13g2_decap_4 FILLER_60_917 ();
 sg13g2_fill_2 FILLER_60_921 ();
 sg13g2_fill_1 FILLER_60_928 ();
 sg13g2_fill_1 FILLER_60_938 ();
 sg13g2_fill_1 FILLER_60_961 ();
 sg13g2_fill_2 FILLER_60_984 ();
 sg13g2_fill_2 FILLER_60_1001 ();
 sg13g2_fill_1 FILLER_60_1003 ();
 sg13g2_decap_8 FILLER_60_1008 ();
 sg13g2_fill_2 FILLER_60_1015 ();
 sg13g2_fill_2 FILLER_60_1027 ();
 sg13g2_fill_2 FILLER_60_1059 ();
 sg13g2_fill_2 FILLER_60_1065 ();
 sg13g2_fill_1 FILLER_60_1067 ();
 sg13g2_fill_2 FILLER_60_1116 ();
 sg13g2_fill_2 FILLER_60_1144 ();
 sg13g2_fill_1 FILLER_60_1146 ();
 sg13g2_decap_4 FILLER_60_1199 ();
 sg13g2_fill_2 FILLER_60_1229 ();
 sg13g2_fill_1 FILLER_60_1237 ();
 sg13g2_fill_2 FILLER_60_1242 ();
 sg13g2_fill_1 FILLER_60_1244 ();
 sg13g2_decap_4 FILLER_60_1258 ();
 sg13g2_fill_2 FILLER_60_1273 ();
 sg13g2_fill_1 FILLER_60_1275 ();
 sg13g2_decap_8 FILLER_60_1281 ();
 sg13g2_fill_1 FILLER_60_1288 ();
 sg13g2_decap_4 FILLER_60_1301 ();
 sg13g2_fill_2 FILLER_60_1311 ();
 sg13g2_fill_1 FILLER_60_1313 ();
 sg13g2_decap_8 FILLER_60_1319 ();
 sg13g2_fill_2 FILLER_60_1326 ();
 sg13g2_fill_1 FILLER_60_1328 ();
 sg13g2_fill_2 FILLER_60_1339 ();
 sg13g2_fill_1 FILLER_60_1341 ();
 sg13g2_fill_2 FILLER_60_1370 ();
 sg13g2_fill_1 FILLER_60_1372 ();
 sg13g2_decap_4 FILLER_60_1377 ();
 sg13g2_fill_1 FILLER_60_1395 ();
 sg13g2_fill_2 FILLER_60_1403 ();
 sg13g2_fill_2 FILLER_60_1415 ();
 sg13g2_fill_1 FILLER_60_1417 ();
 sg13g2_decap_4 FILLER_60_1427 ();
 sg13g2_fill_2 FILLER_60_1434 ();
 sg13g2_decap_8 FILLER_60_1463 ();
 sg13g2_decap_8 FILLER_60_1470 ();
 sg13g2_fill_2 FILLER_60_1477 ();
 sg13g2_fill_1 FILLER_60_1479 ();
 sg13g2_fill_1 FILLER_60_1496 ();
 sg13g2_fill_2 FILLER_60_1536 ();
 sg13g2_fill_2 FILLER_60_1550 ();
 sg13g2_decap_8 FILLER_60_1556 ();
 sg13g2_decap_8 FILLER_60_1563 ();
 sg13g2_fill_2 FILLER_60_1570 ();
 sg13g2_fill_2 FILLER_60_1586 ();
 sg13g2_fill_2 FILLER_60_1597 ();
 sg13g2_fill_1 FILLER_60_1599 ();
 sg13g2_fill_2 FILLER_60_1614 ();
 sg13g2_fill_2 FILLER_60_1660 ();
 sg13g2_decap_8 FILLER_60_1720 ();
 sg13g2_decap_8 FILLER_60_1727 ();
 sg13g2_decap_4 FILLER_60_1734 ();
 sg13g2_fill_2 FILLER_60_1738 ();
 sg13g2_decap_4 FILLER_60_1746 ();
 sg13g2_fill_2 FILLER_60_1750 ();
 sg13g2_fill_1 FILLER_60_1757 ();
 sg13g2_fill_1 FILLER_60_1763 ();
 sg13g2_decap_8 FILLER_60_1776 ();
 sg13g2_fill_2 FILLER_60_1783 ();
 sg13g2_fill_1 FILLER_60_1795 ();
 sg13g2_fill_2 FILLER_60_1803 ();
 sg13g2_fill_2 FILLER_60_1810 ();
 sg13g2_decap_8 FILLER_60_1817 ();
 sg13g2_decap_4 FILLER_60_1824 ();
 sg13g2_fill_1 FILLER_60_1828 ();
 sg13g2_fill_1 FILLER_60_1833 ();
 sg13g2_fill_1 FILLER_60_1854 ();
 sg13g2_fill_2 FILLER_60_1864 ();
 sg13g2_fill_1 FILLER_60_1892 ();
 sg13g2_fill_1 FILLER_60_1908 ();
 sg13g2_fill_2 FILLER_60_1918 ();
 sg13g2_fill_1 FILLER_60_1920 ();
 sg13g2_decap_8 FILLER_60_1925 ();
 sg13g2_decap_8 FILLER_60_1932 ();
 sg13g2_decap_8 FILLER_60_1939 ();
 sg13g2_fill_2 FILLER_60_1946 ();
 sg13g2_fill_1 FILLER_60_1970 ();
 sg13g2_decap_8 FILLER_60_1981 ();
 sg13g2_fill_1 FILLER_60_1992 ();
 sg13g2_decap_8 FILLER_60_2007 ();
 sg13g2_decap_4 FILLER_60_2022 ();
 sg13g2_fill_1 FILLER_60_2101 ();
 sg13g2_decap_4 FILLER_60_2128 ();
 sg13g2_fill_1 FILLER_60_2132 ();
 sg13g2_decap_4 FILLER_60_2137 ();
 sg13g2_fill_2 FILLER_60_2141 ();
 sg13g2_decap_8 FILLER_60_2147 ();
 sg13g2_fill_1 FILLER_60_2154 ();
 sg13g2_fill_2 FILLER_60_2167 ();
 sg13g2_fill_2 FILLER_60_2200 ();
 sg13g2_fill_1 FILLER_60_2202 ();
 sg13g2_fill_2 FILLER_60_2212 ();
 sg13g2_fill_1 FILLER_60_2214 ();
 sg13g2_decap_8 FILLER_60_2227 ();
 sg13g2_decap_8 FILLER_60_2234 ();
 sg13g2_decap_4 FILLER_60_2241 ();
 sg13g2_fill_1 FILLER_60_2245 ();
 sg13g2_decap_8 FILLER_60_2250 ();
 sg13g2_decap_8 FILLER_60_2257 ();
 sg13g2_decap_8 FILLER_60_2264 ();
 sg13g2_fill_1 FILLER_60_2271 ();
 sg13g2_decap_8 FILLER_60_2282 ();
 sg13g2_decap_8 FILLER_60_2289 ();
 sg13g2_decap_8 FILLER_60_2296 ();
 sg13g2_decap_4 FILLER_60_2313 ();
 sg13g2_fill_2 FILLER_60_2317 ();
 sg13g2_fill_1 FILLER_60_2324 ();
 sg13g2_decap_4 FILLER_60_2333 ();
 sg13g2_fill_2 FILLER_60_2389 ();
 sg13g2_fill_2 FILLER_60_2439 ();
 sg13g2_decap_8 FILLER_60_2447 ();
 sg13g2_fill_2 FILLER_60_2454 ();
 sg13g2_decap_8 FILLER_60_2499 ();
 sg13g2_decap_4 FILLER_60_2506 ();
 sg13g2_fill_1 FILLER_60_2510 ();
 sg13g2_fill_1 FILLER_60_2516 ();
 sg13g2_fill_1 FILLER_60_2523 ();
 sg13g2_fill_1 FILLER_60_2534 ();
 sg13g2_fill_2 FILLER_60_2539 ();
 sg13g2_fill_2 FILLER_60_2579 ();
 sg13g2_fill_1 FILLER_60_2581 ();
 sg13g2_fill_2 FILLER_60_2588 ();
 sg13g2_fill_2 FILLER_60_2599 ();
 sg13g2_decap_8 FILLER_60_2605 ();
 sg13g2_decap_8 FILLER_60_2612 ();
 sg13g2_decap_8 FILLER_60_2645 ();
 sg13g2_decap_8 FILLER_60_2652 ();
 sg13g2_decap_8 FILLER_60_2659 ();
 sg13g2_decap_4 FILLER_60_2666 ();
 sg13g2_decap_4 FILLER_61_5 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_decap_4 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_120 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_fill_2 FILLER_61_152 ();
 sg13g2_fill_2 FILLER_61_159 ();
 sg13g2_fill_2 FILLER_61_165 ();
 sg13g2_fill_1 FILLER_61_202 ();
 sg13g2_decap_4 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_237 ();
 sg13g2_decap_4 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_261 ();
 sg13g2_fill_2 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_312 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_decap_8 FILLER_61_319 ();
 sg13g2_decap_8 FILLER_61_326 ();
 sg13g2_decap_8 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_349 ();
 sg13g2_fill_1 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_393 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_decap_8 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_61_435 ();
 sg13g2_decap_4 FILLER_61_452 ();
 sg13g2_fill_1 FILLER_61_456 ();
 sg13g2_fill_2 FILLER_61_465 ();
 sg13g2_fill_1 FILLER_61_471 ();
 sg13g2_fill_1 FILLER_61_484 ();
 sg13g2_fill_2 FILLER_61_494 ();
 sg13g2_fill_1 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_558 ();
 sg13g2_fill_1 FILLER_61_603 ();
 sg13g2_fill_2 FILLER_61_633 ();
 sg13g2_decap_4 FILLER_61_639 ();
 sg13g2_fill_1 FILLER_61_643 ();
 sg13g2_decap_4 FILLER_61_653 ();
 sg13g2_fill_1 FILLER_61_728 ();
 sg13g2_fill_1 FILLER_61_739 ();
 sg13g2_decap_8 FILLER_61_814 ();
 sg13g2_fill_2 FILLER_61_821 ();
 sg13g2_fill_1 FILLER_61_823 ();
 sg13g2_fill_2 FILLER_61_864 ();
 sg13g2_fill_1 FILLER_61_890 ();
 sg13g2_decap_4 FILLER_61_907 ();
 sg13g2_fill_1 FILLER_61_969 ();
 sg13g2_fill_1 FILLER_61_983 ();
 sg13g2_decap_4 FILLER_61_1010 ();
 sg13g2_fill_2 FILLER_61_1014 ();
 sg13g2_fill_1 FILLER_61_1036 ();
 sg13g2_fill_2 FILLER_61_1057 ();
 sg13g2_fill_2 FILLER_61_1098 ();
 sg13g2_fill_1 FILLER_61_1150 ();
 sg13g2_fill_1 FILLER_61_1187 ();
 sg13g2_fill_1 FILLER_61_1203 ();
 sg13g2_fill_2 FILLER_61_1238 ();
 sg13g2_fill_1 FILLER_61_1245 ();
 sg13g2_fill_2 FILLER_61_1287 ();
 sg13g2_fill_2 FILLER_61_1293 ();
 sg13g2_decap_4 FILLER_61_1327 ();
 sg13g2_fill_1 FILLER_61_1331 ();
 sg13g2_decap_8 FILLER_61_1341 ();
 sg13g2_decap_4 FILLER_61_1348 ();
 sg13g2_fill_2 FILLER_61_1365 ();
 sg13g2_fill_1 FILLER_61_1377 ();
 sg13g2_decap_8 FILLER_61_1383 ();
 sg13g2_fill_1 FILLER_61_1412 ();
 sg13g2_fill_1 FILLER_61_1442 ();
 sg13g2_fill_2 FILLER_61_1463 ();
 sg13g2_fill_1 FILLER_61_1473 ();
 sg13g2_fill_1 FILLER_61_1498 ();
 sg13g2_fill_1 FILLER_61_1502 ();
 sg13g2_fill_2 FILLER_61_1548 ();
 sg13g2_fill_2 FILLER_61_1575 ();
 sg13g2_fill_1 FILLER_61_1577 ();
 sg13g2_fill_1 FILLER_61_1588 ();
 sg13g2_fill_1 FILLER_61_1594 ();
 sg13g2_decap_4 FILLER_61_1604 ();
 sg13g2_fill_1 FILLER_61_1608 ();
 sg13g2_fill_2 FILLER_61_1618 ();
 sg13g2_fill_2 FILLER_61_1676 ();
 sg13g2_fill_2 FILLER_61_1711 ();
 sg13g2_fill_2 FILLER_61_1717 ();
 sg13g2_decap_4 FILLER_61_1728 ();
 sg13g2_fill_2 FILLER_61_1748 ();
 sg13g2_fill_1 FILLER_61_1771 ();
 sg13g2_fill_2 FILLER_61_1792 ();
 sg13g2_decap_8 FILLER_61_1811 ();
 sg13g2_decap_4 FILLER_61_1818 ();
 sg13g2_fill_1 FILLER_61_1822 ();
 sg13g2_fill_1 FILLER_61_1848 ();
 sg13g2_fill_1 FILLER_61_1854 ();
 sg13g2_fill_1 FILLER_61_1884 ();
 sg13g2_fill_1 FILLER_61_1893 ();
 sg13g2_fill_1 FILLER_61_1915 ();
 sg13g2_decap_8 FILLER_61_1921 ();
 sg13g2_decap_8 FILLER_61_1928 ();
 sg13g2_decap_8 FILLER_61_1935 ();
 sg13g2_decap_4 FILLER_61_1942 ();
 sg13g2_fill_2 FILLER_61_1946 ();
 sg13g2_fill_2 FILLER_61_1982 ();
 sg13g2_fill_1 FILLER_61_1995 ();
 sg13g2_fill_1 FILLER_61_2001 ();
 sg13g2_fill_2 FILLER_61_2012 ();
 sg13g2_fill_1 FILLER_61_2014 ();
 sg13g2_fill_2 FILLER_61_2042 ();
 sg13g2_fill_1 FILLER_61_2049 ();
 sg13g2_fill_2 FILLER_61_2059 ();
 sg13g2_fill_1 FILLER_61_2061 ();
 sg13g2_fill_2 FILLER_61_2066 ();
 sg13g2_fill_1 FILLER_61_2073 ();
 sg13g2_fill_1 FILLER_61_2078 ();
 sg13g2_decap_8 FILLER_61_2098 ();
 sg13g2_decap_4 FILLER_61_2105 ();
 sg13g2_fill_2 FILLER_61_2109 ();
 sg13g2_decap_8 FILLER_61_2115 ();
 sg13g2_decap_8 FILLER_61_2126 ();
 sg13g2_fill_1 FILLER_61_2151 ();
 sg13g2_decap_4 FILLER_61_2171 ();
 sg13g2_fill_2 FILLER_61_2187 ();
 sg13g2_fill_1 FILLER_61_2214 ();
 sg13g2_decap_4 FILLER_61_2225 ();
 sg13g2_fill_2 FILLER_61_2229 ();
 sg13g2_fill_2 FILLER_61_2263 ();
 sg13g2_fill_1 FILLER_61_2265 ();
 sg13g2_fill_2 FILLER_61_2270 ();
 sg13g2_fill_1 FILLER_61_2272 ();
 sg13g2_fill_2 FILLER_61_2299 ();
 sg13g2_fill_1 FILLER_61_2301 ();
 sg13g2_decap_8 FILLER_61_2328 ();
 sg13g2_fill_1 FILLER_61_2381 ();
 sg13g2_fill_2 FILLER_61_2394 ();
 sg13g2_fill_2 FILLER_61_2479 ();
 sg13g2_fill_2 FILLER_61_2504 ();
 sg13g2_decap_4 FILLER_61_2510 ();
 sg13g2_fill_1 FILLER_61_2519 ();
 sg13g2_fill_2 FILLER_61_2533 ();
 sg13g2_fill_1 FILLER_61_2535 ();
 sg13g2_decap_8 FILLER_61_2544 ();
 sg13g2_fill_1 FILLER_61_2551 ();
 sg13g2_fill_2 FILLER_61_2583 ();
 sg13g2_fill_2 FILLER_61_2598 ();
 sg13g2_fill_1 FILLER_61_2625 ();
 sg13g2_decap_8 FILLER_61_2634 ();
 sg13g2_decap_8 FILLER_61_2641 ();
 sg13g2_decap_8 FILLER_61_2648 ();
 sg13g2_decap_8 FILLER_61_2655 ();
 sg13g2_decap_8 FILLER_61_2662 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_17 ();
 sg13g2_fill_2 FILLER_62_24 ();
 sg13g2_fill_1 FILLER_62_41 ();
 sg13g2_decap_4 FILLER_62_46 ();
 sg13g2_fill_2 FILLER_62_55 ();
 sg13g2_decap_8 FILLER_62_61 ();
 sg13g2_decap_8 FILLER_62_68 ();
 sg13g2_fill_2 FILLER_62_75 ();
 sg13g2_fill_1 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_114 ();
 sg13g2_decap_8 FILLER_62_121 ();
 sg13g2_decap_8 FILLER_62_128 ();
 sg13g2_decap_8 FILLER_62_135 ();
 sg13g2_decap_8 FILLER_62_142 ();
 sg13g2_decap_4 FILLER_62_149 ();
 sg13g2_fill_1 FILLER_62_153 ();
 sg13g2_fill_2 FILLER_62_184 ();
 sg13g2_fill_1 FILLER_62_186 ();
 sg13g2_fill_1 FILLER_62_218 ();
 sg13g2_fill_2 FILLER_62_225 ();
 sg13g2_fill_2 FILLER_62_256 ();
 sg13g2_fill_1 FILLER_62_258 ();
 sg13g2_fill_2 FILLER_62_263 ();
 sg13g2_decap_8 FILLER_62_270 ();
 sg13g2_decap_4 FILLER_62_277 ();
 sg13g2_fill_1 FILLER_62_281 ();
 sg13g2_fill_2 FILLER_62_286 ();
 sg13g2_fill_1 FILLER_62_288 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_fill_2 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_328 ();
 sg13g2_fill_1 FILLER_62_355 ();
 sg13g2_fill_1 FILLER_62_361 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_decap_4 FILLER_62_459 ();
 sg13g2_fill_1 FILLER_62_463 ();
 sg13g2_fill_2 FILLER_62_469 ();
 sg13g2_fill_2 FILLER_62_502 ();
 sg13g2_fill_1 FILLER_62_554 ();
 sg13g2_fill_2 FILLER_62_577 ();
 sg13g2_decap_8 FILLER_62_641 ();
 sg13g2_decap_8 FILLER_62_648 ();
 sg13g2_decap_8 FILLER_62_655 ();
 sg13g2_decap_8 FILLER_62_666 ();
 sg13g2_decap_8 FILLER_62_682 ();
 sg13g2_fill_2 FILLER_62_689 ();
 sg13g2_fill_1 FILLER_62_691 ();
 sg13g2_fill_1 FILLER_62_696 ();
 sg13g2_fill_2 FILLER_62_701 ();
 sg13g2_fill_2 FILLER_62_712 ();
 sg13g2_decap_4 FILLER_62_719 ();
 sg13g2_decap_4 FILLER_62_737 ();
 sg13g2_fill_1 FILLER_62_741 ();
 sg13g2_fill_1 FILLER_62_781 ();
 sg13g2_decap_4 FILLER_62_830 ();
 sg13g2_fill_2 FILLER_62_852 ();
 sg13g2_fill_1 FILLER_62_854 ();
 sg13g2_fill_2 FILLER_62_861 ();
 sg13g2_fill_1 FILLER_62_863 ();
 sg13g2_fill_1 FILLER_62_873 ();
 sg13g2_fill_2 FILLER_62_880 ();
 sg13g2_fill_1 FILLER_62_891 ();
 sg13g2_fill_1 FILLER_62_910 ();
 sg13g2_fill_2 FILLER_62_1007 ();
 sg13g2_fill_1 FILLER_62_1029 ();
 sg13g2_decap_4 FILLER_62_1065 ();
 sg13g2_fill_2 FILLER_62_1069 ();
 sg13g2_fill_2 FILLER_62_1081 ();
 sg13g2_fill_1 FILLER_62_1083 ();
 sg13g2_fill_1 FILLER_62_1115 ();
 sg13g2_fill_2 FILLER_62_1160 ();
 sg13g2_fill_1 FILLER_62_1172 ();
 sg13g2_fill_2 FILLER_62_1177 ();
 sg13g2_fill_2 FILLER_62_1186 ();
 sg13g2_fill_1 FILLER_62_1232 ();
 sg13g2_fill_1 FILLER_62_1237 ();
 sg13g2_fill_1 FILLER_62_1245 ();
 sg13g2_fill_2 FILLER_62_1253 ();
 sg13g2_fill_1 FILLER_62_1278 ();
 sg13g2_fill_1 FILLER_62_1290 ();
 sg13g2_fill_1 FILLER_62_1301 ();
 sg13g2_decap_4 FILLER_62_1311 ();
 sg13g2_fill_1 FILLER_62_1315 ();
 sg13g2_decap_4 FILLER_62_1334 ();
 sg13g2_fill_1 FILLER_62_1342 ();
 sg13g2_fill_2 FILLER_62_1352 ();
 sg13g2_fill_2 FILLER_62_1368 ();
 sg13g2_fill_2 FILLER_62_1411 ();
 sg13g2_fill_1 FILLER_62_1419 ();
 sg13g2_fill_1 FILLER_62_1435 ();
 sg13g2_fill_1 FILLER_62_1483 ();
 sg13g2_fill_2 FILLER_62_1494 ();
 sg13g2_fill_1 FILLER_62_1513 ();
 sg13g2_fill_1 FILLER_62_1530 ();
 sg13g2_fill_2 FILLER_62_1578 ();
 sg13g2_fill_1 FILLER_62_1586 ();
 sg13g2_fill_1 FILLER_62_1605 ();
 sg13g2_decap_4 FILLER_62_1614 ();
 sg13g2_fill_2 FILLER_62_1618 ();
 sg13g2_decap_4 FILLER_62_1641 ();
 sg13g2_fill_1 FILLER_62_1645 ();
 sg13g2_fill_1 FILLER_62_1669 ();
 sg13g2_decap_8 FILLER_62_1686 ();
 sg13g2_fill_2 FILLER_62_1693 ();
 sg13g2_fill_1 FILLER_62_1698 ();
 sg13g2_fill_2 FILLER_62_1709 ();
 sg13g2_decap_4 FILLER_62_1716 ();
 sg13g2_fill_2 FILLER_62_1720 ();
 sg13g2_decap_4 FILLER_62_1737 ();
 sg13g2_fill_1 FILLER_62_1773 ();
 sg13g2_fill_2 FILLER_62_1784 ();
 sg13g2_fill_1 FILLER_62_1790 ();
 sg13g2_fill_2 FILLER_62_1798 ();
 sg13g2_decap_4 FILLER_62_1812 ();
 sg13g2_fill_2 FILLER_62_1816 ();
 sg13g2_decap_4 FILLER_62_1823 ();
 sg13g2_fill_1 FILLER_62_1827 ();
 sg13g2_decap_4 FILLER_62_1832 ();
 sg13g2_fill_1 FILLER_62_1847 ();
 sg13g2_fill_1 FILLER_62_1856 ();
 sg13g2_fill_1 FILLER_62_1863 ();
 sg13g2_fill_1 FILLER_62_1868 ();
 sg13g2_fill_1 FILLER_62_1888 ();
 sg13g2_decap_4 FILLER_62_1915 ();
 sg13g2_decap_8 FILLER_62_1924 ();
 sg13g2_decap_8 FILLER_62_1931 ();
 sg13g2_decap_8 FILLER_62_1938 ();
 sg13g2_fill_2 FILLER_62_1945 ();
 sg13g2_fill_2 FILLER_62_1989 ();
 sg13g2_decap_8 FILLER_62_2003 ();
 sg13g2_decap_4 FILLER_62_2010 ();
 sg13g2_fill_1 FILLER_62_2014 ();
 sg13g2_fill_1 FILLER_62_2029 ();
 sg13g2_fill_1 FILLER_62_2046 ();
 sg13g2_fill_1 FILLER_62_2052 ();
 sg13g2_fill_1 FILLER_62_2058 ();
 sg13g2_fill_1 FILLER_62_2105 ();
 sg13g2_decap_8 FILLER_62_2110 ();
 sg13g2_decap_8 FILLER_62_2157 ();
 sg13g2_fill_1 FILLER_62_2164 ();
 sg13g2_decap_8 FILLER_62_2183 ();
 sg13g2_fill_2 FILLER_62_2190 ();
 sg13g2_fill_1 FILLER_62_2196 ();
 sg13g2_decap_4 FILLER_62_2202 ();
 sg13g2_fill_2 FILLER_62_2216 ();
 sg13g2_fill_1 FILLER_62_2218 ();
 sg13g2_fill_2 FILLER_62_2224 ();
 sg13g2_fill_1 FILLER_62_2226 ();
 sg13g2_fill_2 FILLER_62_2316 ();
 sg13g2_decap_8 FILLER_62_2348 ();
 sg13g2_decap_4 FILLER_62_2355 ();
 sg13g2_fill_2 FILLER_62_2359 ();
 sg13g2_fill_1 FILLER_62_2365 ();
 sg13g2_fill_1 FILLER_62_2397 ();
 sg13g2_fill_1 FILLER_62_2424 ();
 sg13g2_fill_2 FILLER_62_2485 ();
 sg13g2_fill_1 FILLER_62_2541 ();
 sg13g2_fill_2 FILLER_62_2551 ();
 sg13g2_fill_1 FILLER_62_2557 ();
 sg13g2_decap_8 FILLER_62_2647 ();
 sg13g2_decap_8 FILLER_62_2654 ();
 sg13g2_decap_8 FILLER_62_2661 ();
 sg13g2_fill_2 FILLER_62_2668 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_50 ();
 sg13g2_fill_2 FILLER_63_57 ();
 sg13g2_fill_2 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_fill_2 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_138 ();
 sg13g2_decap_8 FILLER_63_145 ();
 sg13g2_decap_8 FILLER_63_152 ();
 sg13g2_decap_8 FILLER_63_159 ();
 sg13g2_fill_2 FILLER_63_166 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_1 FILLER_63_186 ();
 sg13g2_fill_1 FILLER_63_200 ();
 sg13g2_fill_1 FILLER_63_239 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_fill_2 FILLER_63_277 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_decap_8 FILLER_63_285 ();
 sg13g2_fill_2 FILLER_63_297 ();
 sg13g2_fill_1 FILLER_63_303 ();
 sg13g2_decap_4 FILLER_63_314 ();
 sg13g2_decap_8 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_365 ();
 sg13g2_fill_1 FILLER_63_374 ();
 sg13g2_fill_1 FILLER_63_380 ();
 sg13g2_fill_2 FILLER_63_386 ();
 sg13g2_fill_2 FILLER_63_392 ();
 sg13g2_fill_1 FILLER_63_407 ();
 sg13g2_fill_1 FILLER_63_422 ();
 sg13g2_fill_2 FILLER_63_436 ();
 sg13g2_fill_1 FILLER_63_438 ();
 sg13g2_fill_2 FILLER_63_470 ();
 sg13g2_decap_8 FILLER_63_477 ();
 sg13g2_fill_1 FILLER_63_484 ();
 sg13g2_fill_1 FILLER_63_497 ();
 sg13g2_fill_1 FILLER_63_503 ();
 sg13g2_fill_2 FILLER_63_519 ();
 sg13g2_fill_2 FILLER_63_526 ();
 sg13g2_fill_1 FILLER_63_543 ();
 sg13g2_fill_2 FILLER_63_579 ();
 sg13g2_fill_1 FILLER_63_634 ();
 sg13g2_decap_8 FILLER_63_650 ();
 sg13g2_decap_8 FILLER_63_657 ();
 sg13g2_decap_8 FILLER_63_664 ();
 sg13g2_decap_4 FILLER_63_676 ();
 sg13g2_fill_1 FILLER_63_680 ();
 sg13g2_decap_4 FILLER_63_691 ();
 sg13g2_fill_2 FILLER_63_695 ();
 sg13g2_decap_4 FILLER_63_701 ();
 sg13g2_decap_4 FILLER_63_709 ();
 sg13g2_fill_1 FILLER_63_713 ();
 sg13g2_fill_2 FILLER_63_724 ();
 sg13g2_fill_2 FILLER_63_774 ();
 sg13g2_decap_8 FILLER_63_820 ();
 sg13g2_fill_2 FILLER_63_827 ();
 sg13g2_fill_1 FILLER_63_829 ();
 sg13g2_fill_2 FILLER_63_840 ();
 sg13g2_fill_1 FILLER_63_842 ();
 sg13g2_fill_2 FILLER_63_853 ();
 sg13g2_fill_1 FILLER_63_891 ();
 sg13g2_fill_2 FILLER_63_956 ();
 sg13g2_fill_2 FILLER_63_986 ();
 sg13g2_fill_1 FILLER_63_996 ();
 sg13g2_fill_2 FILLER_63_1007 ();
 sg13g2_fill_1 FILLER_63_1029 ();
 sg13g2_decap_4 FILLER_63_1055 ();
 sg13g2_fill_2 FILLER_63_1059 ();
 sg13g2_fill_1 FILLER_63_1090 ();
 sg13g2_fill_2 FILLER_63_1101 ();
 sg13g2_decap_4 FILLER_63_1123 ();
 sg13g2_fill_2 FILLER_63_1131 ();
 sg13g2_decap_8 FILLER_63_1141 ();
 sg13g2_decap_4 FILLER_63_1148 ();
 sg13g2_fill_1 FILLER_63_1193 ();
 sg13g2_decap_8 FILLER_63_1220 ();
 sg13g2_decap_8 FILLER_63_1227 ();
 sg13g2_fill_2 FILLER_63_1234 ();
 sg13g2_fill_1 FILLER_63_1239 ();
 sg13g2_fill_1 FILLER_63_1245 ();
 sg13g2_fill_1 FILLER_63_1251 ();
 sg13g2_fill_1 FILLER_63_1265 ();
 sg13g2_fill_1 FILLER_63_1284 ();
 sg13g2_fill_2 FILLER_63_1292 ();
 sg13g2_decap_8 FILLER_63_1303 ();
 sg13g2_decap_8 FILLER_63_1310 ();
 sg13g2_decap_8 FILLER_63_1317 ();
 sg13g2_fill_1 FILLER_63_1329 ();
 sg13g2_decap_4 FILLER_63_1334 ();
 sg13g2_fill_1 FILLER_63_1338 ();
 sg13g2_decap_4 FILLER_63_1352 ();
 sg13g2_fill_1 FILLER_63_1368 ();
 sg13g2_fill_2 FILLER_63_1384 ();
 sg13g2_fill_1 FILLER_63_1386 ();
 sg13g2_decap_8 FILLER_63_1401 ();
 sg13g2_decap_4 FILLER_63_1408 ();
 sg13g2_fill_2 FILLER_63_1427 ();
 sg13g2_fill_2 FILLER_63_1439 ();
 sg13g2_fill_2 FILLER_63_1507 ();
 sg13g2_fill_1 FILLER_63_1543 ();
 sg13g2_fill_1 FILLER_63_1548 ();
 sg13g2_fill_1 FILLER_63_1554 ();
 sg13g2_fill_2 FILLER_63_1561 ();
 sg13g2_fill_2 FILLER_63_1567 ();
 sg13g2_fill_2 FILLER_63_1599 ();
 sg13g2_fill_1 FILLER_63_1601 ();
 sg13g2_fill_2 FILLER_63_1607 ();
 sg13g2_fill_1 FILLER_63_1609 ();
 sg13g2_decap_8 FILLER_63_1615 ();
 sg13g2_decap_8 FILLER_63_1622 ();
 sg13g2_decap_4 FILLER_63_1629 ();
 sg13g2_fill_1 FILLER_63_1633 ();
 sg13g2_fill_1 FILLER_63_1648 ();
 sg13g2_fill_1 FILLER_63_1653 ();
 sg13g2_fill_1 FILLER_63_1663 ();
 sg13g2_fill_1 FILLER_63_1674 ();
 sg13g2_decap_4 FILLER_63_1679 ();
 sg13g2_fill_2 FILLER_63_1683 ();
 sg13g2_fill_2 FILLER_63_1689 ();
 sg13g2_fill_1 FILLER_63_1691 ();
 sg13g2_decap_8 FILLER_63_1704 ();
 sg13g2_decap_8 FILLER_63_1711 ();
 sg13g2_decap_8 FILLER_63_1718 ();
 sg13g2_decap_4 FILLER_63_1725 ();
 sg13g2_fill_1 FILLER_63_1738 ();
 sg13g2_fill_2 FILLER_63_1744 ();
 sg13g2_fill_1 FILLER_63_1746 ();
 sg13g2_fill_1 FILLER_63_1752 ();
 sg13g2_decap_4 FILLER_63_1786 ();
 sg13g2_fill_1 FILLER_63_1790 ();
 sg13g2_decap_8 FILLER_63_1796 ();
 sg13g2_decap_4 FILLER_63_1803 ();
 sg13g2_decap_4 FILLER_63_1811 ();
 sg13g2_decap_4 FILLER_63_1823 ();
 sg13g2_fill_1 FILLER_63_1827 ();
 sg13g2_fill_2 FILLER_63_1833 ();
 sg13g2_fill_1 FILLER_63_1845 ();
 sg13g2_fill_1 FILLER_63_1857 ();
 sg13g2_fill_1 FILLER_63_1864 ();
 sg13g2_decap_4 FILLER_63_1877 ();
 sg13g2_fill_2 FILLER_63_1916 ();
 sg13g2_decap_8 FILLER_63_1928 ();
 sg13g2_decap_8 FILLER_63_1935 ();
 sg13g2_decap_8 FILLER_63_1942 ();
 sg13g2_fill_1 FILLER_63_1996 ();
 sg13g2_decap_8 FILLER_63_2007 ();
 sg13g2_fill_2 FILLER_63_2014 ();
 sg13g2_fill_2 FILLER_63_2031 ();
 sg13g2_fill_1 FILLER_63_2033 ();
 sg13g2_fill_1 FILLER_63_2045 ();
 sg13g2_decap_4 FILLER_63_2050 ();
 sg13g2_fill_1 FILLER_63_2054 ();
 sg13g2_fill_1 FILLER_63_2068 ();
 sg13g2_decap_4 FILLER_63_2073 ();
 sg13g2_decap_4 FILLER_63_2086 ();
 sg13g2_fill_2 FILLER_63_2095 ();
 sg13g2_fill_2 FILLER_63_2101 ();
 sg13g2_fill_1 FILLER_63_2103 ();
 sg13g2_fill_1 FILLER_63_2144 ();
 sg13g2_decap_4 FILLER_63_2159 ();
 sg13g2_fill_1 FILLER_63_2203 ();
 sg13g2_decap_8 FILLER_63_2210 ();
 sg13g2_fill_2 FILLER_63_2217 ();
 sg13g2_fill_1 FILLER_63_2219 ();
 sg13g2_fill_2 FILLER_63_2225 ();
 sg13g2_decap_4 FILLER_63_2245 ();
 sg13g2_fill_2 FILLER_63_2249 ();
 sg13g2_fill_1 FILLER_63_2261 ();
 sg13g2_fill_2 FILLER_63_2329 ();
 sg13g2_fill_2 FILLER_63_2337 ();
 sg13g2_fill_2 FILLER_63_2344 ();
 sg13g2_decap_8 FILLER_63_2350 ();
 sg13g2_decap_8 FILLER_63_2357 ();
 sg13g2_decap_4 FILLER_63_2364 ();
 sg13g2_fill_2 FILLER_63_2440 ();
 sg13g2_fill_1 FILLER_63_2442 ();
 sg13g2_fill_2 FILLER_63_2536 ();
 sg13g2_fill_2 FILLER_63_2544 ();
 sg13g2_fill_1 FILLER_63_2602 ();
 sg13g2_decap_8 FILLER_63_2625 ();
 sg13g2_decap_8 FILLER_63_2632 ();
 sg13g2_decap_8 FILLER_63_2639 ();
 sg13g2_decap_8 FILLER_63_2646 ();
 sg13g2_decap_8 FILLER_63_2653 ();
 sg13g2_decap_8 FILLER_63_2660 ();
 sg13g2_fill_2 FILLER_63_2667 ();
 sg13g2_fill_1 FILLER_63_2669 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_fill_2 FILLER_64_50 ();
 sg13g2_fill_2 FILLER_64_87 ();
 sg13g2_decap_8 FILLER_64_97 ();
 sg13g2_decap_8 FILLER_64_160 ();
 sg13g2_decap_8 FILLER_64_167 ();
 sg13g2_fill_2 FILLER_64_174 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_fill_1 FILLER_64_198 ();
 sg13g2_decap_8 FILLER_64_222 ();
 sg13g2_decap_4 FILLER_64_229 ();
 sg13g2_fill_1 FILLER_64_249 ();
 sg13g2_fill_2 FILLER_64_278 ();
 sg13g2_fill_1 FILLER_64_280 ();
 sg13g2_decap_4 FILLER_64_312 ();
 sg13g2_fill_2 FILLER_64_316 ();
 sg13g2_fill_2 FILLER_64_322 ();
 sg13g2_fill_1 FILLER_64_329 ();
 sg13g2_fill_1 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_339 ();
 sg13g2_fill_2 FILLER_64_365 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_decap_4 FILLER_64_378 ();
 sg13g2_fill_2 FILLER_64_382 ();
 sg13g2_fill_2 FILLER_64_399 ();
 sg13g2_fill_1 FILLER_64_411 ();
 sg13g2_fill_2 FILLER_64_468 ();
 sg13g2_fill_1 FILLER_64_470 ();
 sg13g2_decap_4 FILLER_64_475 ();
 sg13g2_fill_2 FILLER_64_483 ();
 sg13g2_fill_1 FILLER_64_511 ();
 sg13g2_fill_2 FILLER_64_565 ();
 sg13g2_fill_1 FILLER_64_602 ();
 sg13g2_fill_2 FILLER_64_608 ();
 sg13g2_decap_4 FILLER_64_662 ();
 sg13g2_fill_2 FILLER_64_666 ();
 sg13g2_fill_1 FILLER_64_676 ();
 sg13g2_fill_2 FILLER_64_696 ();
 sg13g2_fill_1 FILLER_64_698 ();
 sg13g2_fill_2 FILLER_64_735 ();
 sg13g2_fill_1 FILLER_64_737 ();
 sg13g2_fill_1 FILLER_64_744 ();
 sg13g2_decap_4 FILLER_64_757 ();
 sg13g2_decap_4 FILLER_64_766 ();
 sg13g2_fill_2 FILLER_64_775 ();
 sg13g2_decap_4 FILLER_64_816 ();
 sg13g2_fill_1 FILLER_64_820 ();
 sg13g2_decap_4 FILLER_64_853 ();
 sg13g2_fill_2 FILLER_64_917 ();
 sg13g2_fill_1 FILLER_64_919 ();
 sg13g2_fill_1 FILLER_64_969 ();
 sg13g2_fill_1 FILLER_64_1047 ();
 sg13g2_fill_2 FILLER_64_1061 ();
 sg13g2_fill_1 FILLER_64_1075 ();
 sg13g2_fill_2 FILLER_64_1081 ();
 sg13g2_fill_1 FILLER_64_1083 ();
 sg13g2_fill_1 FILLER_64_1099 ();
 sg13g2_decap_8 FILLER_64_1118 ();
 sg13g2_decap_8 FILLER_64_1135 ();
 sg13g2_decap_8 FILLER_64_1142 ();
 sg13g2_decap_4 FILLER_64_1149 ();
 sg13g2_fill_2 FILLER_64_1153 ();
 sg13g2_fill_2 FILLER_64_1175 ();
 sg13g2_fill_1 FILLER_64_1200 ();
 sg13g2_decap_8 FILLER_64_1211 ();
 sg13g2_fill_1 FILLER_64_1218 ();
 sg13g2_fill_1 FILLER_64_1225 ();
 sg13g2_fill_1 FILLER_64_1231 ();
 sg13g2_fill_1 FILLER_64_1236 ();
 sg13g2_fill_2 FILLER_64_1246 ();
 sg13g2_fill_1 FILLER_64_1280 ();
 sg13g2_decap_8 FILLER_64_1285 ();
 sg13g2_decap_4 FILLER_64_1292 ();
 sg13g2_decap_4 FILLER_64_1304 ();
 sg13g2_fill_2 FILLER_64_1308 ();
 sg13g2_decap_4 FILLER_64_1317 ();
 sg13g2_fill_1 FILLER_64_1321 ();
 sg13g2_decap_8 FILLER_64_1327 ();
 sg13g2_decap_8 FILLER_64_1334 ();
 sg13g2_decap_4 FILLER_64_1341 ();
 sg13g2_decap_4 FILLER_64_1350 ();
 sg13g2_decap_8 FILLER_64_1364 ();
 sg13g2_decap_8 FILLER_64_1371 ();
 sg13g2_decap_8 FILLER_64_1378 ();
 sg13g2_decap_4 FILLER_64_1398 ();
 sg13g2_fill_1 FILLER_64_1402 ();
 sg13g2_fill_2 FILLER_64_1412 ();
 sg13g2_fill_1 FILLER_64_1424 ();
 sg13g2_fill_2 FILLER_64_1429 ();
 sg13g2_decap_8 FILLER_64_1455 ();
 sg13g2_decap_8 FILLER_64_1462 ();
 sg13g2_decap_4 FILLER_64_1469 ();
 sg13g2_fill_1 FILLER_64_1473 ();
 sg13g2_fill_2 FILLER_64_1511 ();
 sg13g2_fill_1 FILLER_64_1522 ();
 sg13g2_decap_8 FILLER_64_1534 ();
 sg13g2_fill_2 FILLER_64_1541 ();
 sg13g2_fill_2 FILLER_64_1553 ();
 sg13g2_decap_8 FILLER_64_1582 ();
 sg13g2_decap_8 FILLER_64_1594 ();
 sg13g2_decap_8 FILLER_64_1601 ();
 sg13g2_decap_8 FILLER_64_1608 ();
 sg13g2_decap_8 FILLER_64_1615 ();
 sg13g2_decap_8 FILLER_64_1627 ();
 sg13g2_decap_8 FILLER_64_1639 ();
 sg13g2_fill_2 FILLER_64_1646 ();
 sg13g2_fill_1 FILLER_64_1658 ();
 sg13g2_decap_8 FILLER_64_1667 ();
 sg13g2_fill_1 FILLER_64_1674 ();
 sg13g2_decap_8 FILLER_64_1679 ();
 sg13g2_fill_2 FILLER_64_1704 ();
 sg13g2_decap_8 FILLER_64_1710 ();
 sg13g2_decap_8 FILLER_64_1717 ();
 sg13g2_decap_4 FILLER_64_1724 ();
 sg13g2_fill_2 FILLER_64_1728 ();
 sg13g2_fill_2 FILLER_64_1743 ();
 sg13g2_fill_1 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1751 ();
 sg13g2_fill_1 FILLER_64_1758 ();
 sg13g2_fill_1 FILLER_64_1766 ();
 sg13g2_fill_1 FILLER_64_1783 ();
 sg13g2_decap_8 FILLER_64_1807 ();
 sg13g2_decap_8 FILLER_64_1814 ();
 sg13g2_decap_8 FILLER_64_1821 ();
 sg13g2_fill_1 FILLER_64_1828 ();
 sg13g2_decap_8 FILLER_64_1838 ();
 sg13g2_fill_1 FILLER_64_1845 ();
 sg13g2_fill_1 FILLER_64_1851 ();
 sg13g2_fill_1 FILLER_64_1862 ();
 sg13g2_fill_1 FILLER_64_1912 ();
 sg13g2_decap_4 FILLER_64_1918 ();
 sg13g2_fill_1 FILLER_64_1922 ();
 sg13g2_decap_8 FILLER_64_1927 ();
 sg13g2_decap_8 FILLER_64_1934 ();
 sg13g2_decap_8 FILLER_64_1941 ();
 sg13g2_decap_4 FILLER_64_1948 ();
 sg13g2_fill_1 FILLER_64_1952 ();
 sg13g2_fill_1 FILLER_64_2008 ();
 sg13g2_decap_4 FILLER_64_2019 ();
 sg13g2_fill_1 FILLER_64_2033 ();
 sg13g2_fill_1 FILLER_64_2039 ();
 sg13g2_fill_1 FILLER_64_2045 ();
 sg13g2_fill_1 FILLER_64_2052 ();
 sg13g2_fill_1 FILLER_64_2064 ();
 sg13g2_fill_1 FILLER_64_2069 ();
 sg13g2_fill_2 FILLER_64_2078 ();
 sg13g2_fill_1 FILLER_64_2080 ();
 sg13g2_fill_2 FILLER_64_2084 ();
 sg13g2_fill_1 FILLER_64_2086 ();
 sg13g2_decap_8 FILLER_64_2097 ();
 sg13g2_decap_4 FILLER_64_2104 ();
 sg13g2_fill_2 FILLER_64_2108 ();
 sg13g2_decap_4 FILLER_64_2118 ();
 sg13g2_fill_2 FILLER_64_2122 ();
 sg13g2_fill_2 FILLER_64_2154 ();
 sg13g2_fill_1 FILLER_64_2156 ();
 sg13g2_decap_8 FILLER_64_2203 ();
 sg13g2_decap_4 FILLER_64_2210 ();
 sg13g2_fill_1 FILLER_64_2214 ();
 sg13g2_fill_2 FILLER_64_2250 ();
 sg13g2_fill_1 FILLER_64_2252 ();
 sg13g2_fill_1 FILLER_64_2279 ();
 sg13g2_decap_4 FILLER_64_2284 ();
 sg13g2_decap_8 FILLER_64_2292 ();
 sg13g2_fill_1 FILLER_64_2299 ();
 sg13g2_fill_1 FILLER_64_2305 ();
 sg13g2_fill_1 FILLER_64_2311 ();
 sg13g2_fill_2 FILLER_64_2318 ();
 sg13g2_fill_1 FILLER_64_2330 ();
 sg13g2_fill_2 FILLER_64_2337 ();
 sg13g2_fill_2 FILLER_64_2365 ();
 sg13g2_fill_2 FILLER_64_2397 ();
 sg13g2_fill_2 FILLER_64_2405 ();
 sg13g2_decap_4 FILLER_64_2411 ();
 sg13g2_fill_2 FILLER_64_2425 ();
 sg13g2_fill_1 FILLER_64_2427 ();
 sg13g2_fill_2 FILLER_64_2438 ();
 sg13g2_fill_2 FILLER_64_2448 ();
 sg13g2_fill_1 FILLER_64_2467 ();
 sg13g2_fill_1 FILLER_64_2499 ();
 sg13g2_fill_1 FILLER_64_2540 ();
 sg13g2_fill_2 FILLER_64_2567 ();
 sg13g2_fill_1 FILLER_64_2588 ();
 sg13g2_fill_2 FILLER_64_2619 ();
 sg13g2_fill_1 FILLER_64_2621 ();
 sg13g2_decap_8 FILLER_64_2648 ();
 sg13g2_decap_8 FILLER_64_2655 ();
 sg13g2_decap_8 FILLER_64_2662 ();
 sg13g2_fill_1 FILLER_64_2669 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_31 ();
 sg13g2_fill_1 FILLER_65_38 ();
 sg13g2_decap_4 FILLER_65_46 ();
 sg13g2_fill_1 FILLER_65_50 ();
 sg13g2_decap_4 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_93 ();
 sg13g2_fill_1 FILLER_65_115 ();
 sg13g2_decap_4 FILLER_65_168 ();
 sg13g2_fill_2 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_179 ();
 sg13g2_decap_8 FILLER_65_195 ();
 sg13g2_fill_2 FILLER_65_202 ();
 sg13g2_decap_8 FILLER_65_214 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_decap_8 FILLER_65_227 ();
 sg13g2_decap_4 FILLER_65_255 ();
 sg13g2_decap_8 FILLER_65_265 ();
 sg13g2_decap_4 FILLER_65_272 ();
 sg13g2_fill_1 FILLER_65_276 ();
 sg13g2_decap_8 FILLER_65_281 ();
 sg13g2_decap_8 FILLER_65_309 ();
 sg13g2_fill_1 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_fill_1 FILLER_65_343 ();
 sg13g2_fill_2 FILLER_65_353 ();
 sg13g2_decap_4 FILLER_65_381 ();
 sg13g2_decap_4 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_397 ();
 sg13g2_fill_2 FILLER_65_404 ();
 sg13g2_fill_1 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_412 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_decap_4 FILLER_65_426 ();
 sg13g2_fill_2 FILLER_65_430 ();
 sg13g2_fill_2 FILLER_65_473 ();
 sg13g2_decap_8 FILLER_65_484 ();
 sg13g2_fill_1 FILLER_65_491 ();
 sg13g2_fill_1 FILLER_65_523 ();
 sg13g2_fill_2 FILLER_65_550 ();
 sg13g2_fill_2 FILLER_65_578 ();
 sg13g2_fill_2 FILLER_65_585 ();
 sg13g2_fill_1 FILLER_65_591 ();
 sg13g2_fill_1 FILLER_65_632 ();
 sg13g2_fill_2 FILLER_65_659 ();
 sg13g2_decap_4 FILLER_65_719 ();
 sg13g2_decap_8 FILLER_65_727 ();
 sg13g2_decap_8 FILLER_65_734 ();
 sg13g2_decap_4 FILLER_65_741 ();
 sg13g2_fill_2 FILLER_65_745 ();
 sg13g2_fill_1 FILLER_65_751 ();
 sg13g2_fill_1 FILLER_65_778 ();
 sg13g2_decap_4 FILLER_65_810 ();
 sg13g2_fill_1 FILLER_65_814 ();
 sg13g2_fill_1 FILLER_65_819 ();
 sg13g2_decap_4 FILLER_65_846 ();
 sg13g2_fill_2 FILLER_65_850 ();
 sg13g2_decap_4 FILLER_65_878 ();
 sg13g2_fill_1 FILLER_65_882 ();
 sg13g2_fill_1 FILLER_65_893 ();
 sg13g2_fill_1 FILLER_65_961 ();
 sg13g2_fill_1 FILLER_65_967 ();
 sg13g2_fill_2 FILLER_65_974 ();
 sg13g2_fill_2 FILLER_65_979 ();
 sg13g2_fill_1 FILLER_65_1039 ();
 sg13g2_decap_8 FILLER_65_1059 ();
 sg13g2_decap_8 FILLER_65_1066 ();
 sg13g2_decap_8 FILLER_65_1073 ();
 sg13g2_decap_4 FILLER_65_1080 ();
 sg13g2_decap_4 FILLER_65_1140 ();
 sg13g2_fill_1 FILLER_65_1174 ();
 sg13g2_decap_8 FILLER_65_1204 ();
 sg13g2_decap_8 FILLER_65_1211 ();
 sg13g2_fill_2 FILLER_65_1218 ();
 sg13g2_fill_1 FILLER_65_1220 ();
 sg13g2_fill_2 FILLER_65_1236 ();
 sg13g2_fill_1 FILLER_65_1248 ();
 sg13g2_decap_4 FILLER_65_1263 ();
 sg13g2_fill_2 FILLER_65_1273 ();
 sg13g2_fill_2 FILLER_65_1280 ();
 sg13g2_fill_1 FILLER_65_1295 ();
 sg13g2_fill_1 FILLER_65_1301 ();
 sg13g2_fill_1 FILLER_65_1306 ();
 sg13g2_fill_1 FILLER_65_1312 ();
 sg13g2_fill_1 FILLER_65_1318 ();
 sg13g2_decap_4 FILLER_65_1324 ();
 sg13g2_fill_1 FILLER_65_1328 ();
 sg13g2_decap_4 FILLER_65_1337 ();
 sg13g2_fill_2 FILLER_65_1341 ();
 sg13g2_fill_1 FILLER_65_1349 ();
 sg13g2_fill_1 FILLER_65_1359 ();
 sg13g2_fill_2 FILLER_65_1365 ();
 sg13g2_fill_1 FILLER_65_1367 ();
 sg13g2_fill_2 FILLER_65_1381 ();
 sg13g2_fill_2 FILLER_65_1387 ();
 sg13g2_fill_1 FILLER_65_1392 ();
 sg13g2_fill_1 FILLER_65_1401 ();
 sg13g2_fill_1 FILLER_65_1407 ();
 sg13g2_fill_2 FILLER_65_1421 ();
 sg13g2_decap_4 FILLER_65_1428 ();
 sg13g2_fill_2 FILLER_65_1438 ();
 sg13g2_decap_8 FILLER_65_1453 ();
 sg13g2_decap_8 FILLER_65_1460 ();
 sg13g2_decap_8 FILLER_65_1467 ();
 sg13g2_fill_2 FILLER_65_1474 ();
 sg13g2_fill_1 FILLER_65_1476 ();
 sg13g2_fill_1 FILLER_65_1511 ();
 sg13g2_fill_1 FILLER_65_1517 ();
 sg13g2_fill_1 FILLER_65_1528 ();
 sg13g2_decap_8 FILLER_65_1542 ();
 sg13g2_decap_8 FILLER_65_1549 ();
 sg13g2_fill_1 FILLER_65_1556 ();
 sg13g2_decap_4 FILLER_65_1570 ();
 sg13g2_fill_1 FILLER_65_1579 ();
 sg13g2_fill_2 FILLER_65_1590 ();
 sg13g2_fill_1 FILLER_65_1592 ();
 sg13g2_fill_2 FILLER_65_1611 ();
 sg13g2_fill_2 FILLER_65_1622 ();
 sg13g2_fill_1 FILLER_65_1632 ();
 sg13g2_fill_2 FILLER_65_1639 ();
 sg13g2_decap_4 FILLER_65_1644 ();
 sg13g2_fill_2 FILLER_65_1652 ();
 sg13g2_decap_8 FILLER_65_1709 ();
 sg13g2_decap_8 FILLER_65_1716 ();
 sg13g2_decap_4 FILLER_65_1723 ();
 sg13g2_fill_1 FILLER_65_1727 ();
 sg13g2_decap_4 FILLER_65_1748 ();
 sg13g2_fill_1 FILLER_65_1760 ();
 sg13g2_fill_1 FILLER_65_1789 ();
 sg13g2_fill_2 FILLER_65_1822 ();
 sg13g2_decap_4 FILLER_65_1829 ();
 sg13g2_fill_1 FILLER_65_1886 ();
 sg13g2_fill_1 FILLER_65_1910 ();
 sg13g2_fill_1 FILLER_65_1916 ();
 sg13g2_fill_2 FILLER_65_1921 ();
 sg13g2_fill_1 FILLER_65_1923 ();
 sg13g2_fill_2 FILLER_65_1929 ();
 sg13g2_fill_1 FILLER_65_1931 ();
 sg13g2_decap_8 FILLER_65_1941 ();
 sg13g2_decap_8 FILLER_65_1948 ();
 sg13g2_decap_8 FILLER_65_1955 ();
 sg13g2_fill_1 FILLER_65_1976 ();
 sg13g2_fill_2 FILLER_65_1981 ();
 sg13g2_fill_1 FILLER_65_1983 ();
 sg13g2_fill_2 FILLER_65_1988 ();
 sg13g2_fill_1 FILLER_65_1998 ();
 sg13g2_fill_1 FILLER_65_2003 ();
 sg13g2_fill_1 FILLER_65_2009 ();
 sg13g2_fill_1 FILLER_65_2019 ();
 sg13g2_fill_1 FILLER_65_2031 ();
 sg13g2_fill_1 FILLER_65_2045 ();
 sg13g2_fill_1 FILLER_65_2052 ();
 sg13g2_fill_1 FILLER_65_2058 ();
 sg13g2_fill_1 FILLER_65_2064 ();
 sg13g2_fill_1 FILLER_65_2074 ();
 sg13g2_fill_1 FILLER_65_2079 ();
 sg13g2_fill_2 FILLER_65_2093 ();
 sg13g2_fill_1 FILLER_65_2107 ();
 sg13g2_fill_2 FILLER_65_2113 ();
 sg13g2_fill_2 FILLER_65_2119 ();
 sg13g2_fill_1 FILLER_65_2131 ();
 sg13g2_decap_4 FILLER_65_2136 ();
 sg13g2_fill_2 FILLER_65_2140 ();
 sg13g2_fill_2 FILLER_65_2180 ();
 sg13g2_decap_8 FILLER_65_2186 ();
 sg13g2_decap_4 FILLER_65_2193 ();
 sg13g2_fill_2 FILLER_65_2206 ();
 sg13g2_fill_1 FILLER_65_2208 ();
 sg13g2_fill_2 FILLER_65_2215 ();
 sg13g2_fill_1 FILLER_65_2217 ();
 sg13g2_fill_1 FILLER_65_2232 ();
 sg13g2_fill_1 FILLER_65_2293 ();
 sg13g2_decap_4 FILLER_65_2298 ();
 sg13g2_fill_2 FILLER_65_2308 ();
 sg13g2_fill_2 FILLER_65_2356 ();
 sg13g2_fill_2 FILLER_65_2362 ();
 sg13g2_fill_1 FILLER_65_2364 ();
 sg13g2_decap_8 FILLER_65_2401 ();
 sg13g2_decap_8 FILLER_65_2408 ();
 sg13g2_decap_8 FILLER_65_2415 ();
 sg13g2_fill_2 FILLER_65_2422 ();
 sg13g2_fill_2 FILLER_65_2434 ();
 sg13g2_fill_1 FILLER_65_2465 ();
 sg13g2_fill_1 FILLER_65_2498 ();
 sg13g2_fill_1 FILLER_65_2509 ();
 sg13g2_fill_1 FILLER_65_2561 ();
 sg13g2_decap_8 FILLER_65_2650 ();
 sg13g2_decap_8 FILLER_65_2657 ();
 sg13g2_decap_4 FILLER_65_2664 ();
 sg13g2_fill_2 FILLER_65_2668 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_12 ();
 sg13g2_decap_8 FILLER_66_46 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_fill_1 FILLER_66_55 ();
 sg13g2_decap_8 FILLER_66_64 ();
 sg13g2_decap_4 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_139 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_fill_2 FILLER_66_146 ();
 sg13g2_fill_1 FILLER_66_148 ();
 sg13g2_fill_2 FILLER_66_153 ();
 sg13g2_fill_1 FILLER_66_155 ();
 sg13g2_decap_8 FILLER_66_180 ();
 sg13g2_fill_1 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_204 ();
 sg13g2_decap_8 FILLER_66_268 ();
 sg13g2_decap_4 FILLER_66_275 ();
 sg13g2_fill_2 FILLER_66_279 ();
 sg13g2_decap_4 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_288 ();
 sg13g2_decap_4 FILLER_66_295 ();
 sg13g2_decap_8 FILLER_66_304 ();
 sg13g2_decap_4 FILLER_66_311 ();
 sg13g2_fill_2 FILLER_66_315 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_fill_2 FILLER_66_370 ();
 sg13g2_fill_1 FILLER_66_372 ();
 sg13g2_fill_1 FILLER_66_391 ();
 sg13g2_fill_2 FILLER_66_427 ();
 sg13g2_fill_2 FILLER_66_473 ();
 sg13g2_fill_2 FILLER_66_484 ();
 sg13g2_fill_1 FILLER_66_486 ();
 sg13g2_fill_1 FILLER_66_502 ();
 sg13g2_fill_1 FILLER_66_508 ();
 sg13g2_fill_1 FILLER_66_530 ();
 sg13g2_fill_2 FILLER_66_585 ();
 sg13g2_fill_1 FILLER_66_617 ();
 sg13g2_fill_2 FILLER_66_656 ();
 sg13g2_fill_2 FILLER_66_699 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_decap_8 FILLER_66_720 ();
 sg13g2_fill_1 FILLER_66_727 ();
 sg13g2_fill_1 FILLER_66_738 ();
 sg13g2_fill_2 FILLER_66_749 ();
 sg13g2_fill_1 FILLER_66_759 ();
 sg13g2_fill_1 FILLER_66_786 ();
 sg13g2_fill_2 FILLER_66_791 ();
 sg13g2_decap_8 FILLER_66_819 ();
 sg13g2_fill_2 FILLER_66_826 ();
 sg13g2_decap_4 FILLER_66_832 ();
 sg13g2_fill_1 FILLER_66_836 ();
 sg13g2_fill_2 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_66_875 ();
 sg13g2_decap_8 FILLER_66_882 ();
 sg13g2_decap_4 FILLER_66_889 ();
 sg13g2_fill_2 FILLER_66_897 ();
 sg13g2_fill_1 FILLER_66_899 ();
 sg13g2_fill_2 FILLER_66_904 ();
 sg13g2_fill_1 FILLER_66_906 ();
 sg13g2_fill_2 FILLER_66_917 ();
 sg13g2_fill_1 FILLER_66_975 ();
 sg13g2_fill_2 FILLER_66_985 ();
 sg13g2_fill_2 FILLER_66_1008 ();
 sg13g2_fill_1 FILLER_66_1028 ();
 sg13g2_decap_4 FILLER_66_1075 ();
 sg13g2_fill_2 FILLER_66_1079 ();
 sg13g2_fill_2 FILLER_66_1104 ();
 sg13g2_fill_1 FILLER_66_1106 ();
 sg13g2_fill_1 FILLER_66_1173 ();
 sg13g2_decap_8 FILLER_66_1200 ();
 sg13g2_decap_8 FILLER_66_1207 ();
 sg13g2_decap_8 FILLER_66_1214 ();
 sg13g2_fill_2 FILLER_66_1221 ();
 sg13g2_fill_2 FILLER_66_1234 ();
 sg13g2_fill_2 FILLER_66_1242 ();
 sg13g2_fill_1 FILLER_66_1244 ();
 sg13g2_fill_1 FILLER_66_1249 ();
 sg13g2_decap_4 FILLER_66_1265 ();
 sg13g2_fill_1 FILLER_66_1322 ();
 sg13g2_decap_4 FILLER_66_1356 ();
 sg13g2_decap_4 FILLER_66_1370 ();
 sg13g2_decap_8 FILLER_66_1378 ();
 sg13g2_fill_2 FILLER_66_1398 ();
 sg13g2_fill_1 FILLER_66_1400 ();
 sg13g2_fill_1 FILLER_66_1409 ();
 sg13g2_decap_4 FILLER_66_1467 ();
 sg13g2_fill_1 FILLER_66_1471 ();
 sg13g2_fill_2 FILLER_66_1497 ();
 sg13g2_fill_1 FILLER_66_1508 ();
 sg13g2_fill_2 FILLER_66_1518 ();
 sg13g2_fill_1 FILLER_66_1520 ();
 sg13g2_fill_1 FILLER_66_1533 ();
 sg13g2_fill_1 FILLER_66_1539 ();
 sg13g2_decap_8 FILLER_66_1561 ();
 sg13g2_fill_2 FILLER_66_1568 ();
 sg13g2_fill_1 FILLER_66_1570 ();
 sg13g2_decap_8 FILLER_66_1575 ();
 sg13g2_decap_8 FILLER_66_1582 ();
 sg13g2_decap_8 FILLER_66_1589 ();
 sg13g2_fill_2 FILLER_66_1613 ();
 sg13g2_fill_1 FILLER_66_1615 ();
 sg13g2_fill_2 FILLER_66_1620 ();
 sg13g2_fill_1 FILLER_66_1622 ();
 sg13g2_fill_1 FILLER_66_1690 ();
 sg13g2_fill_1 FILLER_66_1695 ();
 sg13g2_fill_1 FILLER_66_1736 ();
 sg13g2_decap_8 FILLER_66_1746 ();
 sg13g2_fill_2 FILLER_66_1753 ();
 sg13g2_decap_4 FILLER_66_1760 ();
 sg13g2_fill_1 FILLER_66_1764 ();
 sg13g2_fill_1 FILLER_66_1770 ();
 sg13g2_fill_1 FILLER_66_1775 ();
 sg13g2_decap_8 FILLER_66_1801 ();
 sg13g2_decap_4 FILLER_66_1808 ();
 sg13g2_fill_1 FILLER_66_1830 ();
 sg13g2_fill_2 FILLER_66_1845 ();
 sg13g2_fill_1 FILLER_66_1847 ();
 sg13g2_fill_2 FILLER_66_1863 ();
 sg13g2_fill_2 FILLER_66_1884 ();
 sg13g2_fill_1 FILLER_66_1892 ();
 sg13g2_fill_2 FILLER_66_1904 ();
 sg13g2_fill_1 FILLER_66_1906 ();
 sg13g2_fill_1 FILLER_66_1912 ();
 sg13g2_fill_2 FILLER_66_1918 ();
 sg13g2_fill_2 FILLER_66_1925 ();
 sg13g2_decap_8 FILLER_66_1937 ();
 sg13g2_fill_2 FILLER_66_1944 ();
 sg13g2_decap_8 FILLER_66_1950 ();
 sg13g2_fill_1 FILLER_66_1975 ();
 sg13g2_decap_4 FILLER_66_1981 ();
 sg13g2_fill_2 FILLER_66_1991 ();
 sg13g2_fill_1 FILLER_66_1993 ();
 sg13g2_fill_1 FILLER_66_2027 ();
 sg13g2_fill_1 FILLER_66_2042 ();
 sg13g2_fill_2 FILLER_66_2047 ();
 sg13g2_fill_1 FILLER_66_2066 ();
 sg13g2_fill_1 FILLER_66_2072 ();
 sg13g2_fill_2 FILLER_66_2099 ();
 sg13g2_fill_1 FILLER_66_2114 ();
 sg13g2_fill_1 FILLER_66_2118 ();
 sg13g2_decap_8 FILLER_66_2127 ();
 sg13g2_fill_2 FILLER_66_2134 ();
 sg13g2_decap_4 FILLER_66_2141 ();
 sg13g2_fill_1 FILLER_66_2157 ();
 sg13g2_fill_2 FILLER_66_2177 ();
 sg13g2_decap_8 FILLER_66_2185 ();
 sg13g2_decap_8 FILLER_66_2192 ();
 sg13g2_decap_8 FILLER_66_2229 ();
 sg13g2_decap_8 FILLER_66_2236 ();
 sg13g2_decap_8 FILLER_66_2243 ();
 sg13g2_decap_4 FILLER_66_2250 ();
 sg13g2_fill_1 FILLER_66_2254 ();
 sg13g2_fill_2 FILLER_66_2263 ();
 sg13g2_fill_1 FILLER_66_2285 ();
 sg13g2_fill_1 FILLER_66_2312 ();
 sg13g2_fill_1 FILLER_66_2317 ();
 sg13g2_fill_2 FILLER_66_2324 ();
 sg13g2_fill_2 FILLER_66_2362 ();
 sg13g2_fill_1 FILLER_66_2367 ();
 sg13g2_decap_4 FILLER_66_2373 ();
 sg13g2_fill_2 FILLER_66_2377 ();
 sg13g2_decap_8 FILLER_66_2402 ();
 sg13g2_decap_8 FILLER_66_2409 ();
 sg13g2_fill_1 FILLER_66_2416 ();
 sg13g2_decap_4 FILLER_66_2420 ();
 sg13g2_decap_8 FILLER_66_2427 ();
 sg13g2_fill_2 FILLER_66_2548 ();
 sg13g2_decap_8 FILLER_66_2619 ();
 sg13g2_decap_4 FILLER_66_2626 ();
 sg13g2_fill_1 FILLER_66_2630 ();
 sg13g2_decap_8 FILLER_66_2635 ();
 sg13g2_decap_8 FILLER_66_2642 ();
 sg13g2_decap_8 FILLER_66_2649 ();
 sg13g2_decap_8 FILLER_66_2656 ();
 sg13g2_decap_8 FILLER_66_2663 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_27 ();
 sg13g2_decap_8 FILLER_67_34 ();
 sg13g2_decap_8 FILLER_67_41 ();
 sg13g2_decap_8 FILLER_67_48 ();
 sg13g2_decap_8 FILLER_67_55 ();
 sg13g2_decap_8 FILLER_67_66 ();
 sg13g2_fill_1 FILLER_67_73 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_fill_2 FILLER_67_131 ();
 sg13g2_decap_4 FILLER_67_143 ();
 sg13g2_fill_2 FILLER_67_178 ();
 sg13g2_decap_8 FILLER_67_215 ();
 sg13g2_decap_8 FILLER_67_222 ();
 sg13g2_fill_2 FILLER_67_229 ();
 sg13g2_fill_1 FILLER_67_231 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_285 ();
 sg13g2_decap_4 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_328 ();
 sg13g2_fill_1 FILLER_67_330 ();
 sg13g2_fill_2 FILLER_67_340 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_decap_4 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_375 ();
 sg13g2_fill_2 FILLER_67_394 ();
 sg13g2_fill_2 FILLER_67_436 ();
 sg13g2_decap_4 FILLER_67_442 ();
 sg13g2_fill_1 FILLER_67_462 ();
 sg13g2_fill_1 FILLER_67_512 ();
 sg13g2_fill_1 FILLER_67_526 ();
 sg13g2_fill_2 FILLER_67_540 ();
 sg13g2_fill_1 FILLER_67_563 ();
 sg13g2_fill_2 FILLER_67_579 ();
 sg13g2_fill_1 FILLER_67_585 ();
 sg13g2_decap_4 FILLER_67_590 ();
 sg13g2_fill_2 FILLER_67_594 ();
 sg13g2_decap_4 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_646 ();
 sg13g2_decap_8 FILLER_67_655 ();
 sg13g2_decap_8 FILLER_67_666 ();
 sg13g2_fill_1 FILLER_67_673 ();
 sg13g2_fill_2 FILLER_67_698 ();
 sg13g2_fill_1 FILLER_67_700 ();
 sg13g2_fill_2 FILLER_67_706 ();
 sg13g2_fill_2 FILLER_67_719 ();
 sg13g2_fill_1 FILLER_67_721 ();
 sg13g2_fill_2 FILLER_67_731 ();
 sg13g2_fill_2 FILLER_67_767 ();
 sg13g2_fill_1 FILLER_67_774 ();
 sg13g2_fill_2 FILLER_67_801 ();
 sg13g2_decap_8 FILLER_67_807 ();
 sg13g2_decap_4 FILLER_67_814 ();
 sg13g2_fill_2 FILLER_67_818 ();
 sg13g2_fill_2 FILLER_67_856 ();
 sg13g2_decap_4 FILLER_67_868 ();
 sg13g2_fill_2 FILLER_67_878 ();
 sg13g2_fill_1 FILLER_67_880 ();
 sg13g2_fill_2 FILLER_67_885 ();
 sg13g2_fill_1 FILLER_67_887 ();
 sg13g2_decap_4 FILLER_67_906 ();
 sg13g2_fill_1 FILLER_67_910 ();
 sg13g2_decap_8 FILLER_67_917 ();
 sg13g2_fill_2 FILLER_67_924 ();
 sg13g2_fill_1 FILLER_67_926 ();
 sg13g2_decap_8 FILLER_67_930 ();
 sg13g2_decap_8 FILLER_67_937 ();
 sg13g2_fill_2 FILLER_67_1024 ();
 sg13g2_fill_1 FILLER_67_1026 ();
 sg13g2_fill_1 FILLER_67_1030 ();
 sg13g2_fill_2 FILLER_67_1038 ();
 sg13g2_fill_1 FILLER_67_1040 ();
 sg13g2_decap_8 FILLER_67_1070 ();
 sg13g2_decap_4 FILLER_67_1077 ();
 sg13g2_fill_2 FILLER_67_1117 ();
 sg13g2_fill_1 FILLER_67_1119 ();
 sg13g2_fill_2 FILLER_67_1184 ();
 sg13g2_decap_8 FILLER_67_1195 ();
 sg13g2_decap_8 FILLER_67_1202 ();
 sg13g2_fill_1 FILLER_67_1209 ();
 sg13g2_fill_1 FILLER_67_1225 ();
 sg13g2_decap_4 FILLER_67_1234 ();
 sg13g2_fill_2 FILLER_67_1243 ();
 sg13g2_fill_1 FILLER_67_1245 ();
 sg13g2_fill_1 FILLER_67_1256 ();
 sg13g2_decap_4 FILLER_67_1263 ();
 sg13g2_fill_1 FILLER_67_1267 ();
 sg13g2_decap_8 FILLER_67_1273 ();
 sg13g2_decap_8 FILLER_67_1280 ();
 sg13g2_decap_8 FILLER_67_1287 ();
 sg13g2_fill_1 FILLER_67_1294 ();
 sg13g2_decap_4 FILLER_67_1317 ();
 sg13g2_decap_8 FILLER_67_1325 ();
 sg13g2_decap_8 FILLER_67_1332 ();
 sg13g2_fill_2 FILLER_67_1339 ();
 sg13g2_fill_1 FILLER_67_1347 ();
 sg13g2_decap_8 FILLER_67_1364 ();
 sg13g2_fill_1 FILLER_67_1386 ();
 sg13g2_fill_2 FILLER_67_1396 ();
 sg13g2_fill_1 FILLER_67_1398 ();
 sg13g2_fill_2 FILLER_67_1420 ();
 sg13g2_fill_2 FILLER_67_1452 ();
 sg13g2_fill_1 FILLER_67_1459 ();
 sg13g2_fill_1 FILLER_67_1490 ();
 sg13g2_fill_2 FILLER_67_1494 ();
 sg13g2_fill_1 FILLER_67_1500 ();
 sg13g2_fill_1 FILLER_67_1506 ();
 sg13g2_fill_2 FILLER_67_1511 ();
 sg13g2_fill_1 FILLER_67_1513 ();
 sg13g2_fill_2 FILLER_67_1518 ();
 sg13g2_fill_1 FILLER_67_1520 ();
 sg13g2_fill_2 FILLER_67_1540 ();
 sg13g2_fill_1 FILLER_67_1542 ();
 sg13g2_decap_8 FILLER_67_1573 ();
 sg13g2_decap_8 FILLER_67_1580 ();
 sg13g2_decap_8 FILLER_67_1587 ();
 sg13g2_decap_4 FILLER_67_1594 ();
 sg13g2_decap_8 FILLER_67_1615 ();
 sg13g2_decap_8 FILLER_67_1622 ();
 sg13g2_fill_1 FILLER_67_1629 ();
 sg13g2_fill_1 FILLER_67_1689 ();
 sg13g2_fill_2 FILLER_67_1702 ();
 sg13g2_fill_1 FILLER_67_1704 ();
 sg13g2_fill_2 FILLER_67_1740 ();
 sg13g2_fill_1 FILLER_67_1742 ();
 sg13g2_decap_8 FILLER_67_1747 ();
 sg13g2_fill_2 FILLER_67_1754 ();
 sg13g2_fill_1 FILLER_67_1756 ();
 sg13g2_decap_4 FILLER_67_1766 ();
 sg13g2_fill_2 FILLER_67_1774 ();
 sg13g2_fill_2 FILLER_67_1786 ();
 sg13g2_fill_1 FILLER_67_1788 ();
 sg13g2_decap_4 FILLER_67_1808 ();
 sg13g2_fill_1 FILLER_67_1812 ();
 sg13g2_fill_1 FILLER_67_1819 ();
 sg13g2_fill_2 FILLER_67_1829 ();
 sg13g2_fill_1 FILLER_67_1851 ();
 sg13g2_fill_1 FILLER_67_1858 ();
 sg13g2_fill_1 FILLER_67_1887 ();
 sg13g2_fill_1 FILLER_67_1898 ();
 sg13g2_fill_2 FILLER_67_1905 ();
 sg13g2_fill_2 FILLER_67_1925 ();
 sg13g2_fill_1 FILLER_67_1927 ();
 sg13g2_fill_2 FILLER_67_1954 ();
 sg13g2_fill_1 FILLER_67_1956 ();
 sg13g2_decap_4 FILLER_67_1961 ();
 sg13g2_fill_2 FILLER_67_1965 ();
 sg13g2_decap_4 FILLER_67_1973 ();
 sg13g2_fill_1 FILLER_67_1982 ();
 sg13g2_fill_2 FILLER_67_1987 ();
 sg13g2_fill_2 FILLER_67_2012 ();
 sg13g2_fill_1 FILLER_67_2014 ();
 sg13g2_fill_2 FILLER_67_2032 ();
 sg13g2_fill_2 FILLER_67_2041 ();
 sg13g2_fill_2 FILLER_67_2068 ();
 sg13g2_fill_2 FILLER_67_2087 ();
 sg13g2_fill_1 FILLER_67_2094 ();
 sg13g2_fill_2 FILLER_67_2099 ();
 sg13g2_fill_2 FILLER_67_2106 ();
 sg13g2_fill_1 FILLER_67_2121 ();
 sg13g2_decap_4 FILLER_67_2130 ();
 sg13g2_decap_8 FILLER_67_2138 ();
 sg13g2_fill_2 FILLER_67_2145 ();
 sg13g2_fill_1 FILLER_67_2152 ();
 sg13g2_fill_1 FILLER_67_2167 ();
 sg13g2_fill_1 FILLER_67_2173 ();
 sg13g2_decap_8 FILLER_67_2178 ();
 sg13g2_decap_4 FILLER_67_2241 ();
 sg13g2_decap_8 FILLER_67_2263 ();
 sg13g2_fill_1 FILLER_67_2270 ();
 sg13g2_fill_2 FILLER_67_2284 ();
 sg13g2_fill_2 FILLER_67_2325 ();
 sg13g2_fill_1 FILLER_67_2353 ();
 sg13g2_decap_4 FILLER_67_2370 ();
 sg13g2_fill_1 FILLER_67_2374 ();
 sg13g2_decap_4 FILLER_67_2411 ();
 sg13g2_fill_2 FILLER_67_2415 ();
 sg13g2_fill_1 FILLER_67_2423 ();
 sg13g2_fill_2 FILLER_67_2468 ();
 sg13g2_fill_1 FILLER_67_2477 ();
 sg13g2_fill_1 FILLER_67_2540 ();
 sg13g2_fill_2 FILLER_67_2580 ();
 sg13g2_fill_2 FILLER_67_2595 ();
 sg13g2_decap_8 FILLER_67_2624 ();
 sg13g2_decap_8 FILLER_67_2631 ();
 sg13g2_decap_8 FILLER_67_2638 ();
 sg13g2_decap_8 FILLER_67_2645 ();
 sg13g2_decap_8 FILLER_67_2652 ();
 sg13g2_decap_8 FILLER_67_2659 ();
 sg13g2_decap_4 FILLER_67_2666 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_4 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_53 ();
 sg13g2_fill_2 FILLER_68_127 ();
 sg13g2_decap_8 FILLER_68_142 ();
 sg13g2_fill_1 FILLER_68_149 ();
 sg13g2_decap_4 FILLER_68_224 ();
 sg13g2_fill_2 FILLER_68_228 ();
 sg13g2_fill_1 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_decap_8 FILLER_68_313 ();
 sg13g2_fill_2 FILLER_68_320 ();
 sg13g2_fill_1 FILLER_68_419 ();
 sg13g2_decap_8 FILLER_68_429 ();
 sg13g2_fill_2 FILLER_68_436 ();
 sg13g2_fill_1 FILLER_68_438 ();
 sg13g2_fill_2 FILLER_68_462 ();
 sg13g2_fill_1 FILLER_68_469 ();
 sg13g2_fill_1 FILLER_68_509 ();
 sg13g2_fill_2 FILLER_68_515 ();
 sg13g2_fill_2 FILLER_68_540 ();
 sg13g2_fill_1 FILLER_68_546 ();
 sg13g2_fill_1 FILLER_68_575 ();
 sg13g2_fill_2 FILLER_68_581 ();
 sg13g2_fill_1 FILLER_68_588 ();
 sg13g2_fill_2 FILLER_68_597 ();
 sg13g2_fill_1 FILLER_68_599 ();
 sg13g2_fill_2 FILLER_68_623 ();
 sg13g2_decap_4 FILLER_68_651 ();
 sg13g2_decap_4 FILLER_68_663 ();
 sg13g2_fill_2 FILLER_68_672 ();
 sg13g2_decap_4 FILLER_68_700 ();
 sg13g2_fill_1 FILLER_68_734 ();
 sg13g2_fill_1 FILLER_68_745 ();
 sg13g2_fill_1 FILLER_68_759 ();
 sg13g2_fill_2 FILLER_68_771 ();
 sg13g2_fill_2 FILLER_68_816 ();
 sg13g2_fill_1 FILLER_68_818 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_fill_2 FILLER_68_845 ();
 sg13g2_fill_1 FILLER_68_847 ();
 sg13g2_fill_1 FILLER_68_883 ();
 sg13g2_fill_2 FILLER_68_889 ();
 sg13g2_decap_8 FILLER_68_947 ();
 sg13g2_fill_1 FILLER_68_957 ();
 sg13g2_fill_2 FILLER_68_962 ();
 sg13g2_fill_1 FILLER_68_1010 ();
 sg13g2_fill_2 FILLER_68_1065 ();
 sg13g2_fill_2 FILLER_68_1072 ();
 sg13g2_decap_4 FILLER_68_1078 ();
 sg13g2_fill_1 FILLER_68_1082 ();
 sg13g2_fill_1 FILLER_68_1126 ();
 sg13g2_fill_1 FILLER_68_1139 ();
 sg13g2_fill_1 FILLER_68_1158 ();
 sg13g2_decap_4 FILLER_68_1163 ();
 sg13g2_fill_1 FILLER_68_1167 ();
 sg13g2_fill_1 FILLER_68_1199 ();
 sg13g2_fill_1 FILLER_68_1238 ();
 sg13g2_fill_1 FILLER_68_1244 ();
 sg13g2_fill_1 FILLER_68_1249 ();
 sg13g2_fill_1 FILLER_68_1255 ();
 sg13g2_decap_8 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1269 ();
 sg13g2_decap_4 FILLER_68_1276 ();
 sg13g2_fill_1 FILLER_68_1280 ();
 sg13g2_fill_1 FILLER_68_1319 ();
 sg13g2_fill_2 FILLER_68_1334 ();
 sg13g2_fill_1 FILLER_68_1336 ();
 sg13g2_fill_1 FILLER_68_1342 ();
 sg13g2_fill_1 FILLER_68_1347 ();
 sg13g2_fill_1 FILLER_68_1353 ();
 sg13g2_fill_1 FILLER_68_1359 ();
 sg13g2_fill_2 FILLER_68_1365 ();
 sg13g2_decap_8 FILLER_68_1372 ();
 sg13g2_fill_1 FILLER_68_1379 ();
 sg13g2_decap_4 FILLER_68_1390 ();
 sg13g2_fill_1 FILLER_68_1394 ();
 sg13g2_fill_1 FILLER_68_1404 ();
 sg13g2_fill_2 FILLER_68_1418 ();
 sg13g2_decap_8 FILLER_68_1464 ();
 sg13g2_fill_2 FILLER_68_1471 ();
 sg13g2_decap_4 FILLER_68_1479 ();
 sg13g2_fill_1 FILLER_68_1483 ();
 sg13g2_decap_4 FILLER_68_1487 ();
 sg13g2_fill_2 FILLER_68_1503 ();
 sg13g2_fill_1 FILLER_68_1505 ();
 sg13g2_fill_2 FILLER_68_1520 ();
 sg13g2_fill_1 FILLER_68_1522 ();
 sg13g2_decap_4 FILLER_68_1528 ();
 sg13g2_fill_1 FILLER_68_1540 ();
 sg13g2_decap_4 FILLER_68_1559 ();
 sg13g2_fill_1 FILLER_68_1569 ();
 sg13g2_decap_8 FILLER_68_1583 ();
 sg13g2_decap_4 FILLER_68_1590 ();
 sg13g2_fill_1 FILLER_68_1594 ();
 sg13g2_decap_8 FILLER_68_1617 ();
 sg13g2_decap_8 FILLER_68_1624 ();
 sg13g2_decap_8 FILLER_68_1653 ();
 sg13g2_decap_8 FILLER_68_1660 ();
 sg13g2_fill_2 FILLER_68_1667 ();
 sg13g2_fill_1 FILLER_68_1669 ();
 sg13g2_fill_1 FILLER_68_1675 ();
 sg13g2_fill_1 FILLER_68_1680 ();
 sg13g2_decap_4 FILLER_68_1690 ();
 sg13g2_fill_1 FILLER_68_1694 ();
 sg13g2_decap_4 FILLER_68_1703 ();
 sg13g2_fill_2 FILLER_68_1707 ();
 sg13g2_fill_1 FILLER_68_1713 ();
 sg13g2_fill_1 FILLER_68_1724 ();
 sg13g2_fill_2 FILLER_68_1755 ();
 sg13g2_fill_2 FILLER_68_1768 ();
 sg13g2_fill_1 FILLER_68_1770 ();
 sg13g2_fill_1 FILLER_68_1781 ();
 sg13g2_fill_1 FILLER_68_1787 ();
 sg13g2_decap_4 FILLER_68_1793 ();
 sg13g2_decap_4 FILLER_68_1802 ();
 sg13g2_decap_8 FILLER_68_1814 ();
 sg13g2_fill_2 FILLER_68_1826 ();
 sg13g2_fill_2 FILLER_68_1834 ();
 sg13g2_fill_1 FILLER_68_1836 ();
 sg13g2_fill_2 FILLER_68_1842 ();
 sg13g2_fill_1 FILLER_68_1844 ();
 sg13g2_decap_4 FILLER_68_1850 ();
 sg13g2_fill_2 FILLER_68_1854 ();
 sg13g2_fill_2 FILLER_68_1866 ();
 sg13g2_fill_2 FILLER_68_1872 ();
 sg13g2_fill_1 FILLER_68_1874 ();
 sg13g2_fill_2 FILLER_68_1879 ();
 sg13g2_fill_1 FILLER_68_1881 ();
 sg13g2_fill_2 FILLER_68_1891 ();
 sg13g2_decap_8 FILLER_68_1922 ();
 sg13g2_decap_4 FILLER_68_1929 ();
 sg13g2_fill_2 FILLER_68_1933 ();
 sg13g2_decap_8 FILLER_68_1939 ();
 sg13g2_decap_8 FILLER_68_1946 ();
 sg13g2_decap_8 FILLER_68_1953 ();
 sg13g2_decap_8 FILLER_68_1960 ();
 sg13g2_fill_1 FILLER_68_1995 ();
 sg13g2_fill_2 FILLER_68_2012 ();
 sg13g2_fill_1 FILLER_68_2014 ();
 sg13g2_fill_1 FILLER_68_2041 ();
 sg13g2_fill_1 FILLER_68_2046 ();
 sg13g2_fill_2 FILLER_68_2051 ();
 sg13g2_fill_1 FILLER_68_2058 ();
 sg13g2_fill_1 FILLER_68_2070 ();
 sg13g2_fill_2 FILLER_68_2095 ();
 sg13g2_decap_4 FILLER_68_2169 ();
 sg13g2_fill_1 FILLER_68_2173 ();
 sg13g2_decap_8 FILLER_68_2184 ();
 sg13g2_fill_2 FILLER_68_2191 ();
 sg13g2_fill_1 FILLER_68_2193 ();
 sg13g2_fill_2 FILLER_68_2198 ();
 sg13g2_decap_4 FILLER_68_2229 ();
 sg13g2_fill_2 FILLER_68_2243 ();
 sg13g2_fill_1 FILLER_68_2245 ();
 sg13g2_fill_1 FILLER_68_2276 ();
 sg13g2_fill_1 FILLER_68_2347 ();
 sg13g2_decap_4 FILLER_68_2418 ();
 sg13g2_fill_2 FILLER_68_2430 ();
 sg13g2_fill_2 FILLER_68_2442 ();
 sg13g2_fill_2 FILLER_68_2448 ();
 sg13g2_fill_1 FILLER_68_2450 ();
 sg13g2_fill_2 FILLER_68_2461 ();
 sg13g2_fill_1 FILLER_68_2463 ();
 sg13g2_fill_2 FILLER_68_2534 ();
 sg13g2_fill_2 FILLER_68_2556 ();
 sg13g2_fill_2 FILLER_68_2562 ();
 sg13g2_fill_2 FILLER_68_2590 ();
 sg13g2_decap_8 FILLER_68_2618 ();
 sg13g2_decap_8 FILLER_68_2625 ();
 sg13g2_decap_8 FILLER_68_2632 ();
 sg13g2_decap_8 FILLER_68_2639 ();
 sg13g2_decap_8 FILLER_68_2646 ();
 sg13g2_decap_8 FILLER_68_2653 ();
 sg13g2_decap_8 FILLER_68_2660 ();
 sg13g2_fill_2 FILLER_68_2667 ();
 sg13g2_fill_1 FILLER_68_2669 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_72 ();
 sg13g2_fill_1 FILLER_69_83 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_decap_4 FILLER_69_111 ();
 sg13g2_fill_2 FILLER_69_120 ();
 sg13g2_decap_4 FILLER_69_127 ();
 sg13g2_decap_4 FILLER_69_157 ();
 sg13g2_decap_4 FILLER_69_165 ();
 sg13g2_fill_1 FILLER_69_169 ();
 sg13g2_fill_1 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_fill_1 FILLER_69_199 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_4 FILLER_69_217 ();
 sg13g2_fill_2 FILLER_69_230 ();
 sg13g2_fill_1 FILLER_69_235 ();
 sg13g2_fill_2 FILLER_69_260 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_fill_1 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_342 ();
 sg13g2_fill_2 FILLER_69_349 ();
 sg13g2_decap_4 FILLER_69_355 ();
 sg13g2_fill_2 FILLER_69_359 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_4 FILLER_69_420 ();
 sg13g2_fill_1 FILLER_69_424 ();
 sg13g2_decap_8 FILLER_69_474 ();
 sg13g2_fill_1 FILLER_69_485 ();
 sg13g2_fill_1 FILLER_69_496 ();
 sg13g2_fill_1 FILLER_69_545 ();
 sg13g2_decap_8 FILLER_69_577 ();
 sg13g2_fill_2 FILLER_69_584 ();
 sg13g2_fill_1 FILLER_69_596 ();
 sg13g2_fill_1 FILLER_69_607 ();
 sg13g2_fill_2 FILLER_69_617 ();
 sg13g2_fill_1 FILLER_69_623 ();
 sg13g2_fill_1 FILLER_69_629 ();
 sg13g2_decap_8 FILLER_69_656 ();
 sg13g2_decap_4 FILLER_69_663 ();
 sg13g2_fill_2 FILLER_69_703 ();
 sg13g2_fill_2 FILLER_69_727 ();
 sg13g2_decap_4 FILLER_69_739 ();
 sg13g2_fill_2 FILLER_69_743 ();
 sg13g2_fill_2 FILLER_69_767 ();
 sg13g2_fill_1 FILLER_69_794 ();
 sg13g2_fill_1 FILLER_69_821 ();
 sg13g2_fill_2 FILLER_69_848 ();
 sg13g2_fill_1 FILLER_69_891 ();
 sg13g2_decap_4 FILLER_69_918 ();
 sg13g2_fill_1 FILLER_69_922 ();
 sg13g2_fill_2 FILLER_69_958 ();
 sg13g2_fill_2 FILLER_69_979 ();
 sg13g2_fill_1 FILLER_69_981 ();
 sg13g2_fill_1 FILLER_69_995 ();
 sg13g2_fill_1 FILLER_69_1002 ();
 sg13g2_fill_1 FILLER_69_1029 ();
 sg13g2_fill_2 FILLER_69_1036 ();
 sg13g2_fill_1 FILLER_69_1038 ();
 sg13g2_decap_8 FILLER_69_1044 ();
 sg13g2_decap_4 FILLER_69_1051 ();
 sg13g2_fill_2 FILLER_69_1059 ();
 sg13g2_fill_1 FILLER_69_1061 ();
 sg13g2_fill_2 FILLER_69_1069 ();
 sg13g2_fill_1 FILLER_69_1087 ();
 sg13g2_fill_2 FILLER_69_1096 ();
 sg13g2_fill_1 FILLER_69_1098 ();
 sg13g2_decap_8 FILLER_69_1135 ();
 sg13g2_decap_8 FILLER_69_1168 ();
 sg13g2_decap_4 FILLER_69_1175 ();
 sg13g2_fill_2 FILLER_69_1179 ();
 sg13g2_decap_8 FILLER_69_1184 ();
 sg13g2_decap_8 FILLER_69_1191 ();
 sg13g2_fill_1 FILLER_69_1198 ();
 sg13g2_fill_1 FILLER_69_1237 ();
 sg13g2_fill_1 FILLER_69_1244 ();
 sg13g2_fill_1 FILLER_69_1250 ();
 sg13g2_fill_1 FILLER_69_1256 ();
 sg13g2_fill_1 FILLER_69_1263 ();
 sg13g2_decap_8 FILLER_69_1272 ();
 sg13g2_fill_2 FILLER_69_1279 ();
 sg13g2_fill_1 FILLER_69_1281 ();
 sg13g2_fill_1 FILLER_69_1312 ();
 sg13g2_decap_4 FILLER_69_1328 ();
 sg13g2_fill_1 FILLER_69_1348 ();
 sg13g2_fill_1 FILLER_69_1354 ();
 sg13g2_fill_2 FILLER_69_1385 ();
 sg13g2_decap_4 FILLER_69_1391 ();
 sg13g2_fill_1 FILLER_69_1395 ();
 sg13g2_fill_1 FILLER_69_1431 ();
 sg13g2_fill_2 FILLER_69_1443 ();
 sg13g2_decap_4 FILLER_69_1455 ();
 sg13g2_decap_4 FILLER_69_1463 ();
 sg13g2_fill_1 FILLER_69_1467 ();
 sg13g2_fill_1 FILLER_69_1472 ();
 sg13g2_fill_2 FILLER_69_1476 ();
 sg13g2_decap_4 FILLER_69_1487 ();
 sg13g2_fill_2 FILLER_69_1499 ();
 sg13g2_fill_1 FILLER_69_1501 ();
 sg13g2_fill_1 FILLER_69_1522 ();
 sg13g2_fill_1 FILLER_69_1526 ();
 sg13g2_decap_8 FILLER_69_1531 ();
 sg13g2_fill_2 FILLER_69_1538 ();
 sg13g2_fill_1 FILLER_69_1591 ();
 sg13g2_decap_8 FILLER_69_1621 ();
 sg13g2_decap_8 FILLER_69_1628 ();
 sg13g2_decap_8 FILLER_69_1635 ();
 sg13g2_fill_1 FILLER_69_1642 ();
 sg13g2_decap_8 FILLER_69_1646 ();
 sg13g2_fill_2 FILLER_69_1653 ();
 sg13g2_fill_1 FILLER_69_1655 ();
 sg13g2_decap_8 FILLER_69_1660 ();
 sg13g2_decap_8 FILLER_69_1667 ();
 sg13g2_decap_4 FILLER_69_1674 ();
 sg13g2_fill_2 FILLER_69_1687 ();
 sg13g2_decap_4 FILLER_69_1728 ();
 sg13g2_fill_1 FILLER_69_1732 ();
 sg13g2_decap_4 FILLER_69_1752 ();
 sg13g2_fill_2 FILLER_69_1756 ();
 sg13g2_decap_4 FILLER_69_1770 ();
 sg13g2_fill_2 FILLER_69_1778 ();
 sg13g2_decap_8 FILLER_69_1823 ();
 sg13g2_decap_8 FILLER_69_1830 ();
 sg13g2_decap_8 FILLER_69_1837 ();
 sg13g2_decap_4 FILLER_69_1848 ();
 sg13g2_fill_2 FILLER_69_1852 ();
 sg13g2_fill_1 FILLER_69_1859 ();
 sg13g2_fill_1 FILLER_69_1864 ();
 sg13g2_decap_4 FILLER_69_1881 ();
 sg13g2_decap_8 FILLER_69_1890 ();
 sg13g2_fill_1 FILLER_69_1897 ();
 sg13g2_fill_2 FILLER_69_1903 ();
 sg13g2_decap_4 FILLER_69_1930 ();
 sg13g2_decap_8 FILLER_69_1945 ();
 sg13g2_decap_4 FILLER_69_1952 ();
 sg13g2_fill_1 FILLER_69_1961 ();
 sg13g2_fill_2 FILLER_69_1968 ();
 sg13g2_fill_1 FILLER_69_2023 ();
 sg13g2_fill_2 FILLER_69_2056 ();
 sg13g2_fill_2 FILLER_69_2071 ();
 sg13g2_fill_2 FILLER_69_2091 ();
 sg13g2_decap_4 FILLER_69_2153 ();
 sg13g2_fill_1 FILLER_69_2165 ();
 sg13g2_fill_1 FILLER_69_2199 ();
 sg13g2_decap_4 FILLER_69_2226 ();
 sg13g2_decap_8 FILLER_69_2235 ();
 sg13g2_decap_4 FILLER_69_2260 ();
 sg13g2_fill_2 FILLER_69_2264 ();
 sg13g2_fill_2 FILLER_69_2321 ();
 sg13g2_decap_8 FILLER_69_2379 ();
 sg13g2_decap_8 FILLER_69_2386 ();
 sg13g2_decap_8 FILLER_69_2393 ();
 sg13g2_decap_4 FILLER_69_2400 ();
 sg13g2_fill_1 FILLER_69_2408 ();
 sg13g2_fill_1 FILLER_69_2431 ();
 sg13g2_decap_8 FILLER_69_2458 ();
 sg13g2_decap_4 FILLER_69_2465 ();
 sg13g2_fill_1 FILLER_69_2469 ();
 sg13g2_fill_2 FILLER_69_2524 ();
 sg13g2_fill_1 FILLER_69_2584 ();
 sg13g2_fill_1 FILLER_69_2596 ();
 sg13g2_fill_2 FILLER_69_2630 ();
 sg13g2_decap_8 FILLER_69_2636 ();
 sg13g2_decap_8 FILLER_69_2643 ();
 sg13g2_decap_8 FILLER_69_2650 ();
 sg13g2_decap_8 FILLER_69_2657 ();
 sg13g2_decap_4 FILLER_69_2664 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_4 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_46 ();
 sg13g2_decap_4 FILLER_70_78 ();
 sg13g2_fill_1 FILLER_70_102 ();
 sg13g2_fill_2 FILLER_70_129 ();
 sg13g2_decap_4 FILLER_70_136 ();
 sg13g2_fill_2 FILLER_70_150 ();
 sg13g2_decap_4 FILLER_70_178 ();
 sg13g2_fill_2 FILLER_70_188 ();
 sg13g2_fill_1 FILLER_70_190 ();
 sg13g2_fill_2 FILLER_70_199 ();
 sg13g2_decap_8 FILLER_70_207 ();
 sg13g2_decap_4 FILLER_70_214 ();
 sg13g2_fill_1 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_2 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_256 ();
 sg13g2_decap_8 FILLER_70_274 ();
 sg13g2_fill_2 FILLER_70_281 ();
 sg13g2_decap_8 FILLER_70_293 ();
 sg13g2_decap_8 FILLER_70_305 ();
 sg13g2_decap_8 FILLER_70_352 ();
 sg13g2_decap_4 FILLER_70_359 ();
 sg13g2_fill_1 FILLER_70_363 ();
 sg13g2_fill_1 FILLER_70_390 ();
 sg13g2_fill_1 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_446 ();
 sg13g2_fill_2 FILLER_70_451 ();
 sg13g2_fill_1 FILLER_70_453 ();
 sg13g2_fill_1 FILLER_70_459 ();
 sg13g2_decap_8 FILLER_70_464 ();
 sg13g2_decap_8 FILLER_70_471 ();
 sg13g2_decap_8 FILLER_70_478 ();
 sg13g2_decap_4 FILLER_70_485 ();
 sg13g2_decap_4 FILLER_70_494 ();
 sg13g2_fill_1 FILLER_70_498 ();
 sg13g2_fill_2 FILLER_70_503 ();
 sg13g2_fill_1 FILLER_70_548 ();
 sg13g2_fill_2 FILLER_70_553 ();
 sg13g2_fill_1 FILLER_70_559 ();
 sg13g2_fill_1 FILLER_70_586 ();
 sg13g2_fill_1 FILLER_70_635 ();
 sg13g2_decap_8 FILLER_70_649 ();
 sg13g2_decap_4 FILLER_70_656 ();
 sg13g2_fill_1 FILLER_70_665 ();
 sg13g2_fill_2 FILLER_70_727 ();
 sg13g2_fill_1 FILLER_70_801 ();
 sg13g2_decap_8 FILLER_70_810 ();
 sg13g2_fill_2 FILLER_70_817 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_decap_4 FILLER_70_882 ();
 sg13g2_fill_2 FILLER_70_886 ();
 sg13g2_fill_1 FILLER_70_897 ();
 sg13g2_decap_4 FILLER_70_924 ();
 sg13g2_fill_2 FILLER_70_938 ();
 sg13g2_fill_2 FILLER_70_944 ();
 sg13g2_fill_1 FILLER_70_956 ();
 sg13g2_fill_1 FILLER_70_997 ();
 sg13g2_fill_1 FILLER_70_1008 ();
 sg13g2_fill_1 FILLER_70_1039 ();
 sg13g2_fill_2 FILLER_70_1056 ();
 sg13g2_decap_8 FILLER_70_1084 ();
 sg13g2_decap_8 FILLER_70_1091 ();
 sg13g2_fill_2 FILLER_70_1098 ();
 sg13g2_fill_1 FILLER_70_1100 ();
 sg13g2_fill_2 FILLER_70_1122 ();
 sg13g2_fill_2 FILLER_70_1158 ();
 sg13g2_fill_1 FILLER_70_1160 ();
 sg13g2_decap_4 FILLER_70_1169 ();
 sg13g2_fill_2 FILLER_70_1202 ();
 sg13g2_fill_1 FILLER_70_1221 ();
 sg13g2_fill_1 FILLER_70_1240 ();
 sg13g2_fill_1 FILLER_70_1246 ();
 sg13g2_fill_2 FILLER_70_1274 ();
 sg13g2_fill_2 FILLER_70_1295 ();
 sg13g2_fill_1 FILLER_70_1302 ();
 sg13g2_fill_1 FILLER_70_1323 ();
 sg13g2_fill_2 FILLER_70_1329 ();
 sg13g2_fill_1 FILLER_70_1331 ();
 sg13g2_fill_1 FILLER_70_1369 ();
 sg13g2_fill_1 FILLER_70_1376 ();
 sg13g2_decap_8 FILLER_70_1398 ();
 sg13g2_fill_1 FILLER_70_1405 ();
 sg13g2_decap_4 FILLER_70_1409 ();
 sg13g2_fill_1 FILLER_70_1418 ();
 sg13g2_fill_1 FILLER_70_1423 ();
 sg13g2_decap_8 FILLER_70_1434 ();
 sg13g2_decap_8 FILLER_70_1441 ();
 sg13g2_decap_4 FILLER_70_1448 ();
 sg13g2_decap_4 FILLER_70_1503 ();
 sg13g2_decap_8 FILLER_70_1530 ();
 sg13g2_decap_8 FILLER_70_1537 ();
 sg13g2_decap_4 FILLER_70_1544 ();
 sg13g2_fill_2 FILLER_70_1548 ();
 sg13g2_decap_4 FILLER_70_1570 ();
 sg13g2_decap_4 FILLER_70_1587 ();
 sg13g2_fill_2 FILLER_70_1591 ();
 sg13g2_decap_8 FILLER_70_1622 ();
 sg13g2_decap_8 FILLER_70_1629 ();
 sg13g2_decap_8 FILLER_70_1636 ();
 sg13g2_fill_1 FILLER_70_1643 ();
 sg13g2_decap_8 FILLER_70_1648 ();
 sg13g2_decap_8 FILLER_70_1655 ();
 sg13g2_fill_1 FILLER_70_1666 ();
 sg13g2_fill_2 FILLER_70_1672 ();
 sg13g2_fill_1 FILLER_70_1691 ();
 sg13g2_fill_2 FILLER_70_1699 ();
 sg13g2_fill_2 FILLER_70_1723 ();
 sg13g2_fill_1 FILLER_70_1725 ();
 sg13g2_decap_4 FILLER_70_1735 ();
 sg13g2_decap_4 FILLER_70_1743 ();
 sg13g2_fill_1 FILLER_70_1747 ();
 sg13g2_decap_8 FILLER_70_1753 ();
 sg13g2_decap_4 FILLER_70_1760 ();
 sg13g2_fill_1 FILLER_70_1772 ();
 sg13g2_fill_2 FILLER_70_1802 ();
 sg13g2_decap_4 FILLER_70_1809 ();
 sg13g2_fill_1 FILLER_70_1813 ();
 sg13g2_fill_1 FILLER_70_1818 ();
 sg13g2_decap_8 FILLER_70_1830 ();
 sg13g2_decap_8 FILLER_70_1837 ();
 sg13g2_decap_8 FILLER_70_1844 ();
 sg13g2_decap_8 FILLER_70_1851 ();
 sg13g2_decap_4 FILLER_70_1858 ();
 sg13g2_decap_4 FILLER_70_1866 ();
 sg13g2_fill_2 FILLER_70_1870 ();
 sg13g2_fill_1 FILLER_70_1897 ();
 sg13g2_decap_8 FILLER_70_1916 ();
 sg13g2_decap_4 FILLER_70_1923 ();
 sg13g2_fill_1 FILLER_70_1927 ();
 sg13g2_decap_4 FILLER_70_1932 ();
 sg13g2_fill_1 FILLER_70_1962 ();
 sg13g2_fill_1 FILLER_70_1968 ();
 sg13g2_fill_2 FILLER_70_2003 ();
 sg13g2_fill_2 FILLER_70_2025 ();
 sg13g2_fill_1 FILLER_70_2034 ();
 sg13g2_fill_2 FILLER_70_2075 ();
 sg13g2_fill_1 FILLER_70_2109 ();
 sg13g2_fill_2 FILLER_70_2114 ();
 sg13g2_fill_2 FILLER_70_2138 ();
 sg13g2_fill_2 FILLER_70_2145 ();
 sg13g2_fill_2 FILLER_70_2152 ();
 sg13g2_decap_8 FILLER_70_2180 ();
 sg13g2_decap_4 FILLER_70_2187 ();
 sg13g2_fill_1 FILLER_70_2191 ();
 sg13g2_fill_1 FILLER_70_2203 ();
 sg13g2_decap_8 FILLER_70_2210 ();
 sg13g2_fill_1 FILLER_70_2217 ();
 sg13g2_fill_1 FILLER_70_2227 ();
 sg13g2_decap_4 FILLER_70_2238 ();
 sg13g2_fill_2 FILLER_70_2247 ();
 sg13g2_fill_2 FILLER_70_2255 ();
 sg13g2_fill_1 FILLER_70_2263 ();
 sg13g2_fill_2 FILLER_70_2268 ();
 sg13g2_fill_1 FILLER_70_2270 ();
 sg13g2_fill_2 FILLER_70_2278 ();
 sg13g2_fill_1 FILLER_70_2286 ();
 sg13g2_fill_1 FILLER_70_2293 ();
 sg13g2_fill_2 FILLER_70_2351 ();
 sg13g2_fill_2 FILLER_70_2358 ();
 sg13g2_fill_1 FILLER_70_2373 ();
 sg13g2_fill_1 FILLER_70_2386 ();
 sg13g2_fill_2 FILLER_70_2423 ();
 sg13g2_fill_1 FILLER_70_2425 ();
 sg13g2_decap_4 FILLER_70_2445 ();
 sg13g2_fill_2 FILLER_70_2449 ();
 sg13g2_decap_4 FILLER_70_2455 ();
 sg13g2_fill_2 FILLER_70_2459 ();
 sg13g2_fill_2 FILLER_70_2467 ();
 sg13g2_decap_8 FILLER_70_2511 ();
 sg13g2_fill_2 FILLER_70_2518 ();
 sg13g2_decap_8 FILLER_70_2525 ();
 sg13g2_decap_4 FILLER_70_2532 ();
 sg13g2_decap_4 FILLER_70_2570 ();
 sg13g2_decap_4 FILLER_70_2577 ();
 sg13g2_decap_8 FILLER_70_2584 ();
 sg13g2_decap_4 FILLER_70_2591 ();
 sg13g2_decap_8 FILLER_70_2631 ();
 sg13g2_decap_8 FILLER_70_2638 ();
 sg13g2_decap_8 FILLER_70_2645 ();
 sg13g2_decap_8 FILLER_70_2652 ();
 sg13g2_decap_8 FILLER_70_2659 ();
 sg13g2_decap_4 FILLER_70_2666 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_decap_4 FILLER_71_150 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_1 FILLER_71_173 ();
 sg13g2_decap_4 FILLER_71_186 ();
 sg13g2_decap_8 FILLER_71_194 ();
 sg13g2_fill_2 FILLER_71_201 ();
 sg13g2_decap_4 FILLER_71_213 ();
 sg13g2_decap_4 FILLER_71_221 ();
 sg13g2_decap_8 FILLER_71_236 ();
 sg13g2_decap_8 FILLER_71_243 ();
 sg13g2_decap_8 FILLER_71_250 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_274 ();
 sg13g2_fill_2 FILLER_71_286 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_4 FILLER_71_315 ();
 sg13g2_fill_2 FILLER_71_345 ();
 sg13g2_fill_1 FILLER_71_347 ();
 sg13g2_fill_1 FILLER_71_353 ();
 sg13g2_decap_8 FILLER_71_359 ();
 sg13g2_decap_4 FILLER_71_366 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_375 ();
 sg13g2_fill_2 FILLER_71_380 ();
 sg13g2_fill_1 FILLER_71_382 ();
 sg13g2_fill_2 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_438 ();
 sg13g2_fill_2 FILLER_71_442 ();
 sg13g2_decap_8 FILLER_71_464 ();
 sg13g2_decap_8 FILLER_71_471 ();
 sg13g2_fill_2 FILLER_71_478 ();
 sg13g2_fill_1 FILLER_71_480 ();
 sg13g2_decap_4 FILLER_71_489 ();
 sg13g2_fill_2 FILLER_71_493 ();
 sg13g2_fill_1 FILLER_71_553 ();
 sg13g2_fill_1 FILLER_71_559 ();
 sg13g2_fill_2 FILLER_71_570 ();
 sg13g2_fill_1 FILLER_71_577 ();
 sg13g2_fill_1 FILLER_71_582 ();
 sg13g2_fill_1 FILLER_71_588 ();
 sg13g2_fill_1 FILLER_71_593 ();
 sg13g2_fill_2 FILLER_71_598 ();
 sg13g2_fill_2 FILLER_71_610 ();
 sg13g2_fill_1 FILLER_71_612 ();
 sg13g2_fill_1 FILLER_71_628 ();
 sg13g2_decap_8 FILLER_71_639 ();
 sg13g2_fill_2 FILLER_71_646 ();
 sg13g2_fill_1 FILLER_71_648 ();
 sg13g2_decap_4 FILLER_71_659 ();
 sg13g2_fill_2 FILLER_71_663 ();
 sg13g2_fill_2 FILLER_71_695 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_fill_1 FILLER_71_718 ();
 sg13g2_decap_4 FILLER_71_725 ();
 sg13g2_fill_2 FILLER_71_772 ();
 sg13g2_fill_1 FILLER_71_784 ();
 sg13g2_fill_1 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_818 ();
 sg13g2_fill_2 FILLER_71_825 ();
 sg13g2_fill_1 FILLER_71_827 ();
 sg13g2_fill_2 FILLER_71_848 ();
 sg13g2_fill_1 FILLER_71_850 ();
 sg13g2_decap_4 FILLER_71_859 ();
 sg13g2_fill_2 FILLER_71_863 ();
 sg13g2_fill_2 FILLER_71_874 ();
 sg13g2_decap_4 FILLER_71_881 ();
 sg13g2_decap_4 FILLER_71_895 ();
 sg13g2_fill_2 FILLER_71_899 ();
 sg13g2_fill_2 FILLER_71_938 ();
 sg13g2_fill_1 FILLER_71_961 ();
 sg13g2_fill_1 FILLER_71_988 ();
 sg13g2_fill_2 FILLER_71_994 ();
 sg13g2_fill_2 FILLER_71_1009 ();
 sg13g2_fill_1 FILLER_71_1011 ();
 sg13g2_decap_8 FILLER_71_1053 ();
 sg13g2_decap_8 FILLER_71_1060 ();
 sg13g2_decap_8 FILLER_71_1067 ();
 sg13g2_decap_8 FILLER_71_1074 ();
 sg13g2_decap_8 FILLER_71_1081 ();
 sg13g2_decap_4 FILLER_71_1088 ();
 sg13g2_fill_2 FILLER_71_1092 ();
 sg13g2_decap_4 FILLER_71_1124 ();
 sg13g2_fill_1 FILLER_71_1128 ();
 sg13g2_fill_1 FILLER_71_1195 ();
 sg13g2_fill_1 FILLER_71_1235 ();
 sg13g2_fill_2 FILLER_71_1246 ();
 sg13g2_fill_2 FILLER_71_1282 ();
 sg13g2_fill_1 FILLER_71_1284 ();
 sg13g2_fill_1 FILLER_71_1289 ();
 sg13g2_fill_1 FILLER_71_1300 ();
 sg13g2_fill_1 FILLER_71_1316 ();
 sg13g2_fill_1 FILLER_71_1360 ();
 sg13g2_fill_2 FILLER_71_1369 ();
 sg13g2_decap_4 FILLER_71_1376 ();
 sg13g2_fill_1 FILLER_71_1380 ();
 sg13g2_decap_8 FILLER_71_1399 ();
 sg13g2_decap_8 FILLER_71_1414 ();
 sg13g2_fill_1 FILLER_71_1421 ();
 sg13g2_decap_4 FILLER_71_1426 ();
 sg13g2_decap_8 FILLER_71_1443 ();
 sg13g2_decap_8 FILLER_71_1450 ();
 sg13g2_decap_8 FILLER_71_1457 ();
 sg13g2_decap_8 FILLER_71_1464 ();
 sg13g2_fill_2 FILLER_71_1471 ();
 sg13g2_fill_1 FILLER_71_1473 ();
 sg13g2_decap_4 FILLER_71_1509 ();
 sg13g2_fill_2 FILLER_71_1513 ();
 sg13g2_fill_2 FILLER_71_1526 ();
 sg13g2_fill_1 FILLER_71_1528 ();
 sg13g2_fill_1 FILLER_71_1535 ();
 sg13g2_fill_1 FILLER_71_1541 ();
 sg13g2_fill_2 FILLER_71_1568 ();
 sg13g2_fill_1 FILLER_71_1570 ();
 sg13g2_fill_2 FILLER_71_1576 ();
 sg13g2_fill_1 FILLER_71_1610 ();
 sg13g2_decap_8 FILLER_71_1625 ();
 sg13g2_decap_8 FILLER_71_1632 ();
 sg13g2_fill_1 FILLER_71_1639 ();
 sg13g2_fill_2 FILLER_71_1653 ();
 sg13g2_fill_1 FILLER_71_1655 ();
 sg13g2_fill_2 FILLER_71_1693 ();
 sg13g2_decap_4 FILLER_71_1725 ();
 sg13g2_fill_1 FILLER_71_1729 ();
 sg13g2_fill_2 FILLER_71_1733 ();
 sg13g2_fill_1 FILLER_71_1735 ();
 sg13g2_fill_2 FILLER_71_1741 ();
 sg13g2_fill_1 FILLER_71_1743 ();
 sg13g2_decap_8 FILLER_71_1749 ();
 sg13g2_decap_8 FILLER_71_1756 ();
 sg13g2_decap_8 FILLER_71_1763 ();
 sg13g2_decap_8 FILLER_71_1770 ();
 sg13g2_decap_8 FILLER_71_1777 ();
 sg13g2_decap_4 FILLER_71_1784 ();
 sg13g2_decap_4 FILLER_71_1814 ();
 sg13g2_fill_2 FILLER_71_1822 ();
 sg13g2_fill_1 FILLER_71_1824 ();
 sg13g2_fill_1 FILLER_71_1830 ();
 sg13g2_decap_8 FILLER_71_1835 ();
 sg13g2_decap_8 FILLER_71_1842 ();
 sg13g2_fill_2 FILLER_71_1849 ();
 sg13g2_fill_1 FILLER_71_1851 ();
 sg13g2_decap_4 FILLER_71_1856 ();
 sg13g2_decap_4 FILLER_71_1870 ();
 sg13g2_fill_1 FILLER_71_1898 ();
 sg13g2_fill_2 FILLER_71_1908 ();
 sg13g2_fill_1 FILLER_71_1910 ();
 sg13g2_fill_2 FILLER_71_1955 ();
 sg13g2_fill_1 FILLER_71_1962 ();
 sg13g2_fill_2 FILLER_71_1967 ();
 sg13g2_fill_1 FILLER_71_1969 ();
 sg13g2_decap_4 FILLER_71_1974 ();
 sg13g2_fill_2 FILLER_71_1989 ();
 sg13g2_fill_1 FILLER_71_2019 ();
 sg13g2_fill_1 FILLER_71_2029 ();
 sg13g2_fill_2 FILLER_71_2052 ();
 sg13g2_fill_2 FILLER_71_2070 ();
 sg13g2_fill_2 FILLER_71_2116 ();
 sg13g2_fill_2 FILLER_71_2161 ();
 sg13g2_decap_8 FILLER_71_2173 ();
 sg13g2_fill_1 FILLER_71_2180 ();
 sg13g2_decap_8 FILLER_71_2190 ();
 sg13g2_decap_4 FILLER_71_2197 ();
 sg13g2_decap_4 FILLER_71_2206 ();
 sg13g2_fill_1 FILLER_71_2210 ();
 sg13g2_fill_1 FILLER_71_2247 ();
 sg13g2_fill_1 FILLER_71_2258 ();
 sg13g2_fill_1 FILLER_71_2263 ();
 sg13g2_fill_2 FILLER_71_2274 ();
 sg13g2_fill_1 FILLER_71_2289 ();
 sg13g2_fill_1 FILLER_71_2316 ();
 sg13g2_fill_1 FILLER_71_2350 ();
 sg13g2_fill_2 FILLER_71_2359 ();
 sg13g2_fill_2 FILLER_71_2371 ();
 sg13g2_decap_8 FILLER_71_2400 ();
 sg13g2_decap_8 FILLER_71_2407 ();
 sg13g2_decap_8 FILLER_71_2414 ();
 sg13g2_decap_4 FILLER_71_2421 ();
 sg13g2_fill_2 FILLER_71_2425 ();
 sg13g2_decap_8 FILLER_71_2431 ();
 sg13g2_decap_4 FILLER_71_2438 ();
 sg13g2_fill_1 FILLER_71_2442 ();
 sg13g2_decap_8 FILLER_71_2503 ();
 sg13g2_decap_8 FILLER_71_2536 ();
 sg13g2_decap_4 FILLER_71_2543 ();
 sg13g2_fill_2 FILLER_71_2550 ();
 sg13g2_fill_1 FILLER_71_2552 ();
 sg13g2_fill_2 FILLER_71_2563 ();
 sg13g2_fill_1 FILLER_71_2601 ();
 sg13g2_fill_2 FILLER_71_2616 ();
 sg13g2_decap_8 FILLER_71_2622 ();
 sg13g2_decap_8 FILLER_71_2629 ();
 sg13g2_decap_8 FILLER_71_2636 ();
 sg13g2_decap_8 FILLER_71_2643 ();
 sg13g2_decap_8 FILLER_71_2650 ();
 sg13g2_decap_8 FILLER_71_2657 ();
 sg13g2_decap_4 FILLER_71_2664 ();
 sg13g2_fill_2 FILLER_71_2668 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_60 ();
 sg13g2_decap_8 FILLER_72_67 ();
 sg13g2_decap_8 FILLER_72_74 ();
 sg13g2_decap_8 FILLER_72_81 ();
 sg13g2_fill_1 FILLER_72_88 ();
 sg13g2_decap_4 FILLER_72_110 ();
 sg13g2_fill_1 FILLER_72_114 ();
 sg13g2_decap_8 FILLER_72_129 ();
 sg13g2_decap_4 FILLER_72_136 ();
 sg13g2_fill_2 FILLER_72_140 ();
 sg13g2_fill_1 FILLER_72_155 ();
 sg13g2_fill_2 FILLER_72_187 ();
 sg13g2_decap_4 FILLER_72_236 ();
 sg13g2_fill_2 FILLER_72_240 ();
 sg13g2_fill_2 FILLER_72_257 ();
 sg13g2_fill_1 FILLER_72_259 ();
 sg13g2_decap_4 FILLER_72_264 ();
 sg13g2_fill_2 FILLER_72_268 ();
 sg13g2_fill_2 FILLER_72_277 ();
 sg13g2_decap_8 FILLER_72_309 ();
 sg13g2_decap_8 FILLER_72_316 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_decap_4 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_368 ();
 sg13g2_fill_1 FILLER_72_374 ();
 sg13g2_fill_1 FILLER_72_380 ();
 sg13g2_fill_1 FILLER_72_390 ();
 sg13g2_fill_2 FILLER_72_400 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_fill_1 FILLER_72_413 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_decap_8 FILLER_72_465 ();
 sg13g2_fill_1 FILLER_72_480 ();
 sg13g2_fill_1 FILLER_72_537 ();
 sg13g2_fill_1 FILLER_72_556 ();
 sg13g2_decap_4 FILLER_72_585 ();
 sg13g2_fill_1 FILLER_72_589 ();
 sg13g2_fill_2 FILLER_72_595 ();
 sg13g2_fill_1 FILLER_72_597 ();
 sg13g2_fill_2 FILLER_72_607 ();
 sg13g2_decap_8 FILLER_72_645 ();
 sg13g2_fill_1 FILLER_72_722 ();
 sg13g2_fill_1 FILLER_72_741 ();
 sg13g2_fill_1 FILLER_72_746 ();
 sg13g2_fill_1 FILLER_72_751 ();
 sg13g2_fill_2 FILLER_72_756 ();
 sg13g2_fill_1 FILLER_72_794 ();
 sg13g2_decap_8 FILLER_72_803 ();
 sg13g2_decap_8 FILLER_72_810 ();
 sg13g2_decap_4 FILLER_72_817 ();
 sg13g2_fill_1 FILLER_72_821 ();
 sg13g2_fill_2 FILLER_72_904 ();
 sg13g2_fill_1 FILLER_72_916 ();
 sg13g2_fill_1 FILLER_72_953 ();
 sg13g2_fill_1 FILLER_72_959 ();
 sg13g2_fill_1 FILLER_72_970 ();
 sg13g2_fill_1 FILLER_72_975 ();
 sg13g2_fill_2 FILLER_72_984 ();
 sg13g2_decap_4 FILLER_72_991 ();
 sg13g2_fill_2 FILLER_72_995 ();
 sg13g2_fill_2 FILLER_72_1005 ();
 sg13g2_fill_2 FILLER_72_1012 ();
 sg13g2_fill_2 FILLER_72_1018 ();
 sg13g2_fill_1 FILLER_72_1020 ();
 sg13g2_fill_1 FILLER_72_1031 ();
 sg13g2_fill_2 FILLER_72_1058 ();
 sg13g2_fill_1 FILLER_72_1060 ();
 sg13g2_decap_8 FILLER_72_1087 ();
 sg13g2_decap_4 FILLER_72_1094 ();
 sg13g2_fill_2 FILLER_72_1098 ();
 sg13g2_fill_2 FILLER_72_1152 ();
 sg13g2_fill_1 FILLER_72_1154 ();
 sg13g2_decap_4 FILLER_72_1165 ();
 sg13g2_fill_1 FILLER_72_1195 ();
 sg13g2_fill_2 FILLER_72_1202 ();
 sg13g2_fill_2 FILLER_72_1214 ();
 sg13g2_fill_1 FILLER_72_1216 ();
 sg13g2_fill_1 FILLER_72_1220 ();
 sg13g2_decap_4 FILLER_72_1227 ();
 sg13g2_fill_1 FILLER_72_1257 ();
 sg13g2_fill_1 FILLER_72_1267 ();
 sg13g2_decap_8 FILLER_72_1273 ();
 sg13g2_fill_1 FILLER_72_1280 ();
 sg13g2_fill_1 FILLER_72_1296 ();
 sg13g2_fill_1 FILLER_72_1302 ();
 sg13g2_fill_2 FILLER_72_1308 ();
 sg13g2_fill_2 FILLER_72_1314 ();
 sg13g2_fill_2 FILLER_72_1321 ();
 sg13g2_fill_1 FILLER_72_1331 ();
 sg13g2_fill_2 FILLER_72_1337 ();
 sg13g2_fill_1 FILLER_72_1343 ();
 sg13g2_fill_1 FILLER_72_1349 ();
 sg13g2_fill_1 FILLER_72_1354 ();
 sg13g2_fill_1 FILLER_72_1368 ();
 sg13g2_fill_2 FILLER_72_1379 ();
 sg13g2_decap_8 FILLER_72_1391 ();
 sg13g2_fill_2 FILLER_72_1398 ();
 sg13g2_fill_1 FILLER_72_1400 ();
 sg13g2_fill_1 FILLER_72_1405 ();
 sg13g2_decap_8 FILLER_72_1442 ();
 sg13g2_decap_4 FILLER_72_1449 ();
 sg13g2_fill_1 FILLER_72_1453 ();
 sg13g2_fill_1 FILLER_72_1506 ();
 sg13g2_fill_1 FILLER_72_1519 ();
 sg13g2_decap_4 FILLER_72_1525 ();
 sg13g2_fill_2 FILLER_72_1529 ();
 sg13g2_fill_1 FILLER_72_1538 ();
 sg13g2_decap_8 FILLER_72_1544 ();
 sg13g2_decap_4 FILLER_72_1551 ();
 sg13g2_fill_1 FILLER_72_1570 ();
 sg13g2_fill_1 FILLER_72_1589 ();
 sg13g2_fill_2 FILLER_72_1603 ();
 sg13g2_fill_1 FILLER_72_1605 ();
 sg13g2_fill_1 FILLER_72_1624 ();
 sg13g2_decap_4 FILLER_72_1651 ();
 sg13g2_fill_2 FILLER_72_1689 ();
 sg13g2_decap_8 FILLER_72_1695 ();
 sg13g2_fill_2 FILLER_72_1702 ();
 sg13g2_fill_1 FILLER_72_1704 ();
 sg13g2_fill_2 FILLER_72_1719 ();
 sg13g2_fill_2 FILLER_72_1725 ();
 sg13g2_decap_4 FILLER_72_1731 ();
 sg13g2_fill_2 FILLER_72_1735 ();
 sg13g2_fill_1 FILLER_72_1743 ();
 sg13g2_fill_2 FILLER_72_1758 ();
 sg13g2_fill_1 FILLER_72_1760 ();
 sg13g2_decap_8 FILLER_72_1765 ();
 sg13g2_decap_8 FILLER_72_1772 ();
 sg13g2_fill_1 FILLER_72_1779 ();
 sg13g2_decap_8 FILLER_72_1830 ();
 sg13g2_fill_2 FILLER_72_1837 ();
 sg13g2_fill_1 FILLER_72_1839 ();
 sg13g2_fill_1 FILLER_72_1844 ();
 sg13g2_fill_1 FILLER_72_1863 ();
 sg13g2_fill_1 FILLER_72_1869 ();
 sg13g2_fill_1 FILLER_72_1875 ();
 sg13g2_decap_4 FILLER_72_1887 ();
 sg13g2_fill_2 FILLER_72_1896 ();
 sg13g2_fill_1 FILLER_72_1907 ();
 sg13g2_decap_8 FILLER_72_1925 ();
 sg13g2_decap_8 FILLER_72_1932 ();
 sg13g2_decap_8 FILLER_72_1939 ();
 sg13g2_decap_8 FILLER_72_1950 ();
 sg13g2_fill_1 FILLER_72_1957 ();
 sg13g2_decap_8 FILLER_72_1962 ();
 sg13g2_fill_2 FILLER_72_1969 ();
 sg13g2_decap_8 FILLER_72_1976 ();
 sg13g2_decap_4 FILLER_72_1983 ();
 sg13g2_fill_2 FILLER_72_1987 ();
 sg13g2_fill_1 FILLER_72_2012 ();
 sg13g2_fill_2 FILLER_72_2016 ();
 sg13g2_fill_2 FILLER_72_2027 ();
 sg13g2_fill_2 FILLER_72_2043 ();
 sg13g2_fill_1 FILLER_72_2066 ();
 sg13g2_fill_2 FILLER_72_2105 ();
 sg13g2_fill_1 FILLER_72_2118 ();
 sg13g2_fill_1 FILLER_72_2129 ();
 sg13g2_fill_1 FILLER_72_2140 ();
 sg13g2_decap_8 FILLER_72_2177 ();
 sg13g2_decap_8 FILLER_72_2184 ();
 sg13g2_fill_2 FILLER_72_2191 ();
 sg13g2_fill_1 FILLER_72_2193 ();
 sg13g2_fill_2 FILLER_72_2226 ();
 sg13g2_fill_1 FILLER_72_2348 ();
 sg13g2_fill_2 FILLER_72_2383 ();
 sg13g2_decap_8 FILLER_72_2425 ();
 sg13g2_decap_4 FILLER_72_2432 ();
 sg13g2_fill_1 FILLER_72_2440 ();
 sg13g2_decap_4 FILLER_72_2494 ();
 sg13g2_fill_2 FILLER_72_2528 ();
 sg13g2_fill_1 FILLER_72_2591 ();
 sg13g2_decap_8 FILLER_72_2632 ();
 sg13g2_decap_8 FILLER_72_2639 ();
 sg13g2_decap_8 FILLER_72_2646 ();
 sg13g2_decap_8 FILLER_72_2653 ();
 sg13g2_decap_8 FILLER_72_2660 ();
 sg13g2_fill_2 FILLER_72_2667 ();
 sg13g2_fill_1 FILLER_72_2669 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_54 ();
 sg13g2_decap_8 FILLER_73_61 ();
 sg13g2_decap_8 FILLER_73_68 ();
 sg13g2_decap_8 FILLER_73_75 ();
 sg13g2_decap_4 FILLER_73_82 ();
 sg13g2_fill_1 FILLER_73_86 ();
 sg13g2_decap_8 FILLER_73_97 ();
 sg13g2_decap_8 FILLER_73_104 ();
 sg13g2_decap_8 FILLER_73_111 ();
 sg13g2_fill_2 FILLER_73_118 ();
 sg13g2_decap_4 FILLER_73_151 ();
 sg13g2_fill_1 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_177 ();
 sg13g2_fill_1 FILLER_73_182 ();
 sg13g2_fill_1 FILLER_73_214 ();
 sg13g2_decap_8 FILLER_73_227 ();
 sg13g2_fill_1 FILLER_73_234 ();
 sg13g2_decap_8 FILLER_73_323 ();
 sg13g2_decap_8 FILLER_73_330 ();
 sg13g2_fill_1 FILLER_73_341 ();
 sg13g2_fill_1 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_418 ();
 sg13g2_fill_2 FILLER_73_422 ();
 sg13g2_decap_8 FILLER_73_428 ();
 sg13g2_decap_4 FILLER_73_439 ();
 sg13g2_fill_1 FILLER_73_451 ();
 sg13g2_fill_2 FILLER_73_500 ();
 sg13g2_fill_2 FILLER_73_507 ();
 sg13g2_fill_1 FILLER_73_521 ();
 sg13g2_fill_1 FILLER_73_557 ();
 sg13g2_fill_1 FILLER_73_573 ();
 sg13g2_fill_1 FILLER_73_585 ();
 sg13g2_decap_8 FILLER_73_590 ();
 sg13g2_fill_2 FILLER_73_597 ();
 sg13g2_fill_2 FILLER_73_603 ();
 sg13g2_fill_1 FILLER_73_605 ();
 sg13g2_fill_2 FILLER_73_622 ();
 sg13g2_fill_1 FILLER_73_624 ();
 sg13g2_decap_8 FILLER_73_629 ();
 sg13g2_decap_8 FILLER_73_636 ();
 sg13g2_fill_2 FILLER_73_643 ();
 sg13g2_fill_1 FILLER_73_645 ();
 sg13g2_decap_8 FILLER_73_652 ();
 sg13g2_fill_2 FILLER_73_659 ();
 sg13g2_fill_1 FILLER_73_661 ();
 sg13g2_decap_4 FILLER_73_672 ();
 sg13g2_fill_2 FILLER_73_716 ();
 sg13g2_fill_2 FILLER_73_724 ();
 sg13g2_fill_2 FILLER_73_739 ();
 sg13g2_fill_1 FILLER_73_741 ();
 sg13g2_fill_1 FILLER_73_746 ();
 sg13g2_fill_1 FILLER_73_752 ();
 sg13g2_fill_2 FILLER_73_758 ();
 sg13g2_fill_2 FILLER_73_775 ();
 sg13g2_fill_1 FILLER_73_781 ();
 sg13g2_fill_2 FILLER_73_788 ();
 sg13g2_fill_1 FILLER_73_829 ();
 sg13g2_fill_1 FILLER_73_836 ();
 sg13g2_fill_1 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_874 ();
 sg13g2_decap_8 FILLER_73_881 ();
 sg13g2_fill_2 FILLER_73_893 ();
 sg13g2_fill_1 FILLER_73_895 ();
 sg13g2_fill_1 FILLER_73_910 ();
 sg13g2_fill_2 FILLER_73_941 ();
 sg13g2_fill_2 FILLER_73_948 ();
 sg13g2_decap_8 FILLER_73_980 ();
 sg13g2_decap_8 FILLER_73_987 ();
 sg13g2_decap_4 FILLER_73_994 ();
 sg13g2_fill_1 FILLER_73_998 ();
 sg13g2_decap_8 FILLER_73_1015 ();
 sg13g2_decap_8 FILLER_73_1022 ();
 sg13g2_decap_8 FILLER_73_1029 ();
 sg13g2_fill_2 FILLER_73_1036 ();
 sg13g2_fill_2 FILLER_73_1062 ();
 sg13g2_fill_1 FILLER_73_1064 ();
 sg13g2_fill_2 FILLER_73_1115 ();
 sg13g2_fill_1 FILLER_73_1117 ();
 sg13g2_fill_2 FILLER_73_1158 ();
 sg13g2_fill_1 FILLER_73_1160 ();
 sg13g2_decap_4 FILLER_73_1187 ();
 sg13g2_fill_1 FILLER_73_1191 ();
 sg13g2_fill_2 FILLER_73_1205 ();
 sg13g2_fill_2 FILLER_73_1233 ();
 sg13g2_fill_1 FILLER_73_1235 ();
 sg13g2_decap_4 FILLER_73_1257 ();
 sg13g2_fill_2 FILLER_73_1261 ();
 sg13g2_decap_4 FILLER_73_1273 ();
 sg13g2_fill_2 FILLER_73_1277 ();
 sg13g2_decap_8 FILLER_73_1317 ();
 sg13g2_decap_4 FILLER_73_1324 ();
 sg13g2_fill_2 FILLER_73_1328 ();
 sg13g2_fill_2 FILLER_73_1340 ();
 sg13g2_fill_1 FILLER_73_1342 ();
 sg13g2_decap_8 FILLER_73_1379 ();
 sg13g2_fill_1 FILLER_73_1386 ();
 sg13g2_decap_8 FILLER_73_1423 ();
 sg13g2_decap_8 FILLER_73_1430 ();
 sg13g2_fill_2 FILLER_73_1437 ();
 sg13g2_decap_8 FILLER_73_1443 ();
 sg13g2_fill_2 FILLER_73_1450 ();
 sg13g2_fill_1 FILLER_73_1452 ();
 sg13g2_fill_1 FILLER_73_1499 ();
 sg13g2_fill_1 FILLER_73_1505 ();
 sg13g2_fill_1 FILLER_73_1511 ();
 sg13g2_fill_1 FILLER_73_1520 ();
 sg13g2_fill_1 FILLER_73_1525 ();
 sg13g2_decap_8 FILLER_73_1530 ();
 sg13g2_decap_8 FILLER_73_1537 ();
 sg13g2_decap_8 FILLER_73_1544 ();
 sg13g2_fill_2 FILLER_73_1551 ();
 sg13g2_fill_1 FILLER_73_1561 ();
 sg13g2_decap_4 FILLER_73_1604 ();
 sg13g2_fill_1 FILLER_73_1608 ();
 sg13g2_fill_2 FILLER_73_1614 ();
 sg13g2_decap_8 FILLER_73_1625 ();
 sg13g2_fill_1 FILLER_73_1632 ();
 sg13g2_fill_1 FILLER_73_1637 ();
 sg13g2_fill_2 FILLER_73_1648 ();
 sg13g2_fill_1 FILLER_73_1655 ();
 sg13g2_fill_2 FILLER_73_1660 ();
 sg13g2_fill_1 FILLER_73_1685 ();
 sg13g2_fill_2 FILLER_73_1691 ();
 sg13g2_fill_1 FILLER_73_1693 ();
 sg13g2_fill_1 FILLER_73_1712 ();
 sg13g2_fill_1 FILLER_73_1717 ();
 sg13g2_fill_1 FILLER_73_1727 ();
 sg13g2_fill_2 FILLER_73_1736 ();
 sg13g2_fill_1 FILLER_73_1738 ();
 sg13g2_decap_4 FILLER_73_1757 ();
 sg13g2_fill_2 FILLER_73_1761 ();
 sg13g2_decap_8 FILLER_73_1767 ();
 sg13g2_decap_8 FILLER_73_1774 ();
 sg13g2_fill_1 FILLER_73_1795 ();
 sg13g2_fill_1 FILLER_73_1824 ();
 sg13g2_decap_4 FILLER_73_1830 ();
 sg13g2_fill_2 FILLER_73_1834 ();
 sg13g2_fill_2 FILLER_73_1840 ();
 sg13g2_fill_2 FILLER_73_1846 ();
 sg13g2_fill_1 FILLER_73_1894 ();
 sg13g2_fill_1 FILLER_73_1908 ();
 sg13g2_fill_1 FILLER_73_1917 ();
 sg13g2_fill_2 FILLER_73_1927 ();
 sg13g2_fill_1 FILLER_73_1929 ();
 sg13g2_fill_1 FILLER_73_1938 ();
 sg13g2_decap_8 FILLER_73_1944 ();
 sg13g2_fill_1 FILLER_73_1951 ();
 sg13g2_fill_1 FILLER_73_1960 ();
 sg13g2_decap_4 FILLER_73_1966 ();
 sg13g2_fill_2 FILLER_73_1970 ();
 sg13g2_fill_1 FILLER_73_1977 ();
 sg13g2_fill_1 FILLER_73_1982 ();
 sg13g2_fill_1 FILLER_73_1988 ();
 sg13g2_fill_2 FILLER_73_1998 ();
 sg13g2_fill_1 FILLER_73_2000 ();
 sg13g2_decap_4 FILLER_73_2006 ();
 sg13g2_fill_1 FILLER_73_2010 ();
 sg13g2_decap_4 FILLER_73_2020 ();
 sg13g2_decap_4 FILLER_73_2028 ();
 sg13g2_fill_2 FILLER_73_2032 ();
 sg13g2_fill_1 FILLER_73_2060 ();
 sg13g2_fill_1 FILLER_73_2087 ();
 sg13g2_fill_1 FILLER_73_2098 ();
 sg13g2_fill_1 FILLER_73_2105 ();
 sg13g2_fill_2 FILLER_73_2142 ();
 sg13g2_fill_2 FILLER_73_2185 ();
 sg13g2_fill_1 FILLER_73_2234 ();
 sg13g2_fill_2 FILLER_73_2245 ();
 sg13g2_fill_1 FILLER_73_2315 ();
 sg13g2_fill_1 FILLER_73_2334 ();
 sg13g2_fill_2 FILLER_73_2354 ();
 sg13g2_fill_1 FILLER_73_2360 ();
 sg13g2_fill_1 FILLER_73_2365 ();
 sg13g2_decap_4 FILLER_73_2411 ();
 sg13g2_fill_2 FILLER_73_2451 ();
 sg13g2_decap_4 FILLER_73_2457 ();
 sg13g2_fill_2 FILLER_73_2503 ();
 sg13g2_fill_1 FILLER_73_2571 ();
 sg13g2_fill_1 FILLER_73_2581 ();
 sg13g2_fill_2 FILLER_73_2595 ();
 sg13g2_decap_8 FILLER_73_2603 ();
 sg13g2_decap_8 FILLER_73_2610 ();
 sg13g2_decap_8 FILLER_73_2617 ();
 sg13g2_decap_8 FILLER_73_2624 ();
 sg13g2_decap_8 FILLER_73_2631 ();
 sg13g2_decap_8 FILLER_73_2638 ();
 sg13g2_decap_8 FILLER_73_2645 ();
 sg13g2_decap_8 FILLER_73_2652 ();
 sg13g2_decap_8 FILLER_73_2659 ();
 sg13g2_decap_4 FILLER_73_2666 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_fill_1 FILLER_74_42 ();
 sg13g2_decap_4 FILLER_74_83 ();
 sg13g2_fill_1 FILLER_74_87 ();
 sg13g2_decap_8 FILLER_74_93 ();
 sg13g2_decap_4 FILLER_74_100 ();
 sg13g2_fill_2 FILLER_74_104 ();
 sg13g2_decap_4 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_155 ();
 sg13g2_fill_2 FILLER_74_178 ();
 sg13g2_fill_1 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_206 ();
 sg13g2_fill_1 FILLER_74_217 ();
 sg13g2_fill_1 FILLER_74_244 ();
 sg13g2_fill_1 FILLER_74_249 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_decap_4 FILLER_74_316 ();
 sg13g2_fill_2 FILLER_74_320 ();
 sg13g2_decap_8 FILLER_74_327 ();
 sg13g2_decap_8 FILLER_74_334 ();
 sg13g2_decap_4 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_345 ();
 sg13g2_decap_8 FILLER_74_424 ();
 sg13g2_decap_4 FILLER_74_436 ();
 sg13g2_fill_2 FILLER_74_471 ();
 sg13g2_fill_1 FILLER_74_477 ();
 sg13g2_fill_2 FILLER_74_488 ();
 sg13g2_fill_1 FILLER_74_516 ();
 sg13g2_fill_2 FILLER_74_556 ();
 sg13g2_decap_4 FILLER_74_593 ();
 sg13g2_fill_2 FILLER_74_602 ();
 sg13g2_fill_1 FILLER_74_634 ();
 sg13g2_fill_2 FILLER_74_674 ();
 sg13g2_decap_4 FILLER_74_685 ();
 sg13g2_decap_8 FILLER_74_707 ();
 sg13g2_decap_4 FILLER_74_714 ();
 sg13g2_fill_1 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_fill_2 FILLER_74_800 ();
 sg13g2_fill_1 FILLER_74_802 ();
 sg13g2_fill_2 FILLER_74_839 ();
 sg13g2_fill_1 FILLER_74_841 ();
 sg13g2_fill_2 FILLER_74_846 ();
 sg13g2_decap_4 FILLER_74_872 ();
 sg13g2_fill_2 FILLER_74_884 ();
 sg13g2_fill_1 FILLER_74_886 ();
 sg13g2_fill_2 FILLER_74_949 ();
 sg13g2_decap_4 FILLER_74_957 ();
 sg13g2_decap_4 FILLER_74_971 ();
 sg13g2_fill_2 FILLER_74_985 ();
 sg13g2_fill_1 FILLER_74_987 ();
 sg13g2_decap_4 FILLER_74_994 ();
 sg13g2_decap_8 FILLER_74_1034 ();
 sg13g2_decap_8 FILLER_74_1041 ();
 sg13g2_decap_8 FILLER_74_1048 ();
 sg13g2_fill_1 FILLER_74_1055 ();
 sg13g2_decap_8 FILLER_74_1083 ();
 sg13g2_fill_2 FILLER_74_1090 ();
 sg13g2_fill_2 FILLER_74_1118 ();
 sg13g2_fill_1 FILLER_74_1120 ();
 sg13g2_fill_2 FILLER_74_1131 ();
 sg13g2_fill_1 FILLER_74_1133 ();
 sg13g2_decap_8 FILLER_74_1220 ();
 sg13g2_decap_8 FILLER_74_1227 ();
 sg13g2_fill_1 FILLER_74_1234 ();
 sg13g2_decap_8 FILLER_74_1255 ();
 sg13g2_fill_2 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1326 ();
 sg13g2_decap_4 FILLER_74_1333 ();
 sg13g2_fill_1 FILLER_74_1337 ();
 sg13g2_fill_2 FILLER_74_1364 ();
 sg13g2_decap_4 FILLER_74_1392 ();
 sg13g2_fill_1 FILLER_74_1396 ();
 sg13g2_decap_4 FILLER_74_1459 ();
 sg13g2_fill_1 FILLER_74_1463 ();
 sg13g2_decap_8 FILLER_74_1468 ();
 sg13g2_fill_1 FILLER_74_1475 ();
 sg13g2_decap_4 FILLER_74_1481 ();
 sg13g2_fill_1 FILLER_74_1485 ();
 sg13g2_decap_4 FILLER_74_1490 ();
 sg13g2_fill_1 FILLER_74_1518 ();
 sg13g2_fill_2 FILLER_74_1528 ();
 sg13g2_fill_1 FILLER_74_1534 ();
 sg13g2_decap_8 FILLER_74_1553 ();
 sg13g2_decap_8 FILLER_74_1560 ();
 sg13g2_fill_2 FILLER_74_1567 ();
 sg13g2_fill_1 FILLER_74_1569 ();
 sg13g2_fill_2 FILLER_74_1579 ();
 sg13g2_fill_1 FILLER_74_1581 ();
 sg13g2_fill_2 FILLER_74_1592 ();
 sg13g2_decap_4 FILLER_74_1598 ();
 sg13g2_fill_1 FILLER_74_1602 ();
 sg13g2_fill_1 FILLER_74_1608 ();
 sg13g2_decap_8 FILLER_74_1614 ();
 sg13g2_decap_8 FILLER_74_1621 ();
 sg13g2_decap_8 FILLER_74_1628 ();
 sg13g2_decap_8 FILLER_74_1635 ();
 sg13g2_decap_8 FILLER_74_1642 ();
 sg13g2_fill_2 FILLER_74_1649 ();
 sg13g2_fill_1 FILLER_74_1651 ();
 sg13g2_fill_2 FILLER_74_1662 ();
 sg13g2_fill_1 FILLER_74_1664 ();
 sg13g2_fill_2 FILLER_74_1669 ();
 sg13g2_fill_1 FILLER_74_1671 ();
 sg13g2_fill_1 FILLER_74_1677 ();
 sg13g2_fill_1 FILLER_74_1684 ();
 sg13g2_fill_1 FILLER_74_1690 ();
 sg13g2_decap_8 FILLER_74_1695 ();
 sg13g2_fill_1 FILLER_74_1702 ();
 sg13g2_decap_8 FILLER_74_1708 ();
 sg13g2_fill_1 FILLER_74_1715 ();
 sg13g2_fill_1 FILLER_74_1720 ();
 sg13g2_fill_1 FILLER_74_1726 ();
 sg13g2_fill_1 FILLER_74_1731 ();
 sg13g2_fill_1 FILLER_74_1751 ();
 sg13g2_decap_8 FILLER_74_1762 ();
 sg13g2_decap_8 FILLER_74_1769 ();
 sg13g2_decap_8 FILLER_74_1776 ();
 sg13g2_decap_8 FILLER_74_1783 ();
 sg13g2_fill_1 FILLER_74_1790 ();
 sg13g2_fill_1 FILLER_74_1816 ();
 sg13g2_fill_1 FILLER_74_1822 ();
 sg13g2_fill_2 FILLER_74_1854 ();
 sg13g2_fill_1 FILLER_74_1875 ();
 sg13g2_fill_1 FILLER_74_1905 ();
 sg13g2_fill_2 FILLER_74_1921 ();
 sg13g2_fill_1 FILLER_74_1923 ();
 sg13g2_decap_8 FILLER_74_1947 ();
 sg13g2_fill_1 FILLER_74_1954 ();
 sg13g2_fill_2 FILLER_74_1960 ();
 sg13g2_decap_8 FILLER_74_1988 ();
 sg13g2_decap_8 FILLER_74_1995 ();
 sg13g2_decap_8 FILLER_74_2002 ();
 sg13g2_decap_4 FILLER_74_2009 ();
 sg13g2_fill_2 FILLER_74_2039 ();
 sg13g2_decap_8 FILLER_74_2045 ();
 sg13g2_decap_4 FILLER_74_2152 ();
 sg13g2_fill_2 FILLER_74_2156 ();
 sg13g2_fill_1 FILLER_74_2166 ();
 sg13g2_fill_1 FILLER_74_2181 ();
 sg13g2_fill_2 FILLER_74_2186 ();
 sg13g2_fill_2 FILLER_74_2221 ();
 sg13g2_fill_1 FILLER_74_2303 ();
 sg13g2_fill_1 FILLER_74_2327 ();
 sg13g2_fill_1 FILLER_74_2373 ();
 sg13g2_fill_1 FILLER_74_2403 ();
 sg13g2_fill_2 FILLER_74_2438 ();
 sg13g2_decap_4 FILLER_74_2492 ();
 sg13g2_fill_1 FILLER_74_2496 ();
 sg13g2_decap_8 FILLER_74_2507 ();
 sg13g2_fill_2 FILLER_74_2514 ();
 sg13g2_fill_1 FILLER_74_2516 ();
 sg13g2_decap_4 FILLER_74_2536 ();
 sg13g2_fill_2 FILLER_74_2540 ();
 sg13g2_fill_2 FILLER_74_2568 ();
 sg13g2_fill_1 FILLER_74_2570 ();
 sg13g2_fill_2 FILLER_74_2575 ();
 sg13g2_decap_8 FILLER_74_2617 ();
 sg13g2_decap_8 FILLER_74_2624 ();
 sg13g2_decap_8 FILLER_74_2631 ();
 sg13g2_decap_8 FILLER_74_2638 ();
 sg13g2_decap_8 FILLER_74_2645 ();
 sg13g2_decap_8 FILLER_74_2652 ();
 sg13g2_decap_8 FILLER_74_2659 ();
 sg13g2_decap_4 FILLER_74_2666 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_fill_1 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_87 ();
 sg13g2_decap_8 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_100 ();
 sg13g2_fill_1 FILLER_75_137 ();
 sg13g2_decap_8 FILLER_75_143 ();
 sg13g2_decap_8 FILLER_75_150 ();
 sg13g2_fill_1 FILLER_75_157 ();
 sg13g2_decap_8 FILLER_75_179 ();
 sg13g2_decap_8 FILLER_75_186 ();
 sg13g2_decap_8 FILLER_75_193 ();
 sg13g2_decap_4 FILLER_75_200 ();
 sg13g2_fill_1 FILLER_75_207 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_decap_4 FILLER_75_220 ();
 sg13g2_fill_2 FILLER_75_224 ();
 sg13g2_decap_4 FILLER_75_230 ();
 sg13g2_fill_2 FILLER_75_234 ();
 sg13g2_decap_4 FILLER_75_244 ();
 sg13g2_fill_2 FILLER_75_248 ();
 sg13g2_fill_2 FILLER_75_254 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_fill_1 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_330 ();
 sg13g2_fill_2 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_fill_2 FILLER_75_350 ();
 sg13g2_decap_4 FILLER_75_357 ();
 sg13g2_fill_2 FILLER_75_361 ();
 sg13g2_decap_4 FILLER_75_371 ();
 sg13g2_fill_1 FILLER_75_375 ();
 sg13g2_decap_8 FILLER_75_380 ();
 sg13g2_decap_4 FILLER_75_387 ();
 sg13g2_fill_1 FILLER_75_391 ();
 sg13g2_fill_2 FILLER_75_410 ();
 sg13g2_fill_1 FILLER_75_412 ();
 sg13g2_decap_8 FILLER_75_421 ();
 sg13g2_decap_4 FILLER_75_428 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_465 ();
 sg13g2_fill_1 FILLER_75_485 ();
 sg13g2_fill_1 FILLER_75_515 ();
 sg13g2_decap_8 FILLER_75_582 ();
 sg13g2_fill_1 FILLER_75_589 ();
 sg13g2_decap_8 FILLER_75_594 ();
 sg13g2_fill_1 FILLER_75_601 ();
 sg13g2_fill_2 FILLER_75_612 ();
 sg13g2_fill_1 FILLER_75_614 ();
 sg13g2_decap_4 FILLER_75_628 ();
 sg13g2_fill_1 FILLER_75_632 ();
 sg13g2_fill_2 FILLER_75_644 ();
 sg13g2_fill_1 FILLER_75_646 ();
 sg13g2_decap_4 FILLER_75_657 ();
 sg13g2_fill_2 FILLER_75_661 ();
 sg13g2_fill_2 FILLER_75_671 ();
 sg13g2_decap_4 FILLER_75_712 ();
 sg13g2_fill_1 FILLER_75_746 ();
 sg13g2_fill_1 FILLER_75_761 ();
 sg13g2_fill_2 FILLER_75_776 ();
 sg13g2_decap_8 FILLER_75_788 ();
 sg13g2_fill_2 FILLER_75_795 ();
 sg13g2_fill_1 FILLER_75_797 ();
 sg13g2_decap_4 FILLER_75_804 ();
 sg13g2_fill_1 FILLER_75_808 ();
 sg13g2_fill_2 FILLER_75_813 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_fill_1 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_856 ();
 sg13g2_decap_8 FILLER_75_863 ();
 sg13g2_fill_1 FILLER_75_870 ();
 sg13g2_fill_2 FILLER_75_877 ();
 sg13g2_fill_1 FILLER_75_879 ();
 sg13g2_decap_8 FILLER_75_893 ();
 sg13g2_fill_1 FILLER_75_900 ();
 sg13g2_fill_2 FILLER_75_911 ();
 sg13g2_fill_1 FILLER_75_913 ();
 sg13g2_fill_1 FILLER_75_920 ();
 sg13g2_fill_2 FILLER_75_925 ();
 sg13g2_decap_4 FILLER_75_931 ();
 sg13g2_fill_1 FILLER_75_948 ();
 sg13g2_fill_2 FILLER_75_980 ();
 sg13g2_decap_8 FILLER_75_1040 ();
 sg13g2_decap_8 FILLER_75_1047 ();
 sg13g2_fill_1 FILLER_75_1054 ();
 sg13g2_decap_8 FILLER_75_1059 ();
 sg13g2_fill_1 FILLER_75_1066 ();
 sg13g2_decap_8 FILLER_75_1071 ();
 sg13g2_decap_4 FILLER_75_1078 ();
 sg13g2_fill_2 FILLER_75_1082 ();
 sg13g2_decap_4 FILLER_75_1114 ();
 sg13g2_fill_1 FILLER_75_1118 ();
 sg13g2_decap_8 FILLER_75_1162 ();
 sg13g2_decap_8 FILLER_75_1169 ();
 sg13g2_decap_8 FILLER_75_1180 ();
 sg13g2_fill_1 FILLER_75_1197 ();
 sg13g2_fill_2 FILLER_75_1225 ();
 sg13g2_decap_8 FILLER_75_1253 ();
 sg13g2_decap_8 FILLER_75_1260 ();
 sg13g2_decap_8 FILLER_75_1271 ();
 sg13g2_fill_2 FILLER_75_1278 ();
 sg13g2_fill_1 FILLER_75_1280 ();
 sg13g2_fill_2 FILLER_75_1294 ();
 sg13g2_decap_8 FILLER_75_1326 ();
 sg13g2_decap_8 FILLER_75_1333 ();
 sg13g2_fill_2 FILLER_75_1340 ();
 sg13g2_fill_1 FILLER_75_1342 ();
 sg13g2_fill_2 FILLER_75_1347 ();
 sg13g2_fill_1 FILLER_75_1349 ();
 sg13g2_decap_8 FILLER_75_1353 ();
 sg13g2_decap_4 FILLER_75_1364 ();
 sg13g2_fill_1 FILLER_75_1368 ();
 sg13g2_decap_8 FILLER_75_1383 ();
 sg13g2_decap_8 FILLER_75_1390 ();
 sg13g2_decap_4 FILLER_75_1397 ();
 sg13g2_fill_1 FILLER_75_1411 ();
 sg13g2_fill_1 FILLER_75_1438 ();
 sg13g2_fill_2 FILLER_75_1465 ();
 sg13g2_fill_2 FILLER_75_1470 ();
 sg13g2_fill_1 FILLER_75_1472 ();
 sg13g2_decap_8 FILLER_75_1477 ();
 sg13g2_fill_2 FILLER_75_1528 ();
 sg13g2_decap_8 FILLER_75_1535 ();
 sg13g2_decap_8 FILLER_75_1545 ();
 sg13g2_decap_8 FILLER_75_1552 ();
 sg13g2_fill_1 FILLER_75_1570 ();
 sg13g2_fill_2 FILLER_75_1580 ();
 sg13g2_fill_1 FILLER_75_1591 ();
 sg13g2_decap_8 FILLER_75_1596 ();
 sg13g2_fill_1 FILLER_75_1607 ();
 sg13g2_decap_8 FILLER_75_1623 ();
 sg13g2_fill_2 FILLER_75_1630 ();
 sg13g2_fill_1 FILLER_75_1636 ();
 sg13g2_fill_2 FILLER_75_1641 ();
 sg13g2_fill_2 FILLER_75_1711 ();
 sg13g2_decap_4 FILLER_75_1729 ();
 sg13g2_fill_1 FILLER_75_1733 ();
 sg13g2_fill_2 FILLER_75_1751 ();
 sg13g2_decap_8 FILLER_75_1779 ();
 sg13g2_decap_8 FILLER_75_1786 ();
 sg13g2_decap_8 FILLER_75_1793 ();
 sg13g2_fill_1 FILLER_75_1800 ();
 sg13g2_fill_1 FILLER_75_1806 ();
 sg13g2_fill_1 FILLER_75_1831 ();
 sg13g2_fill_2 FILLER_75_1853 ();
 sg13g2_fill_1 FILLER_75_1911 ();
 sg13g2_fill_1 FILLER_75_1916 ();
 sg13g2_decap_8 FILLER_75_1922 ();
 sg13g2_fill_2 FILLER_75_2022 ();
 sg13g2_fill_1 FILLER_75_2024 ();
 sg13g2_decap_4 FILLER_75_2055 ();
 sg13g2_fill_1 FILLER_75_2066 ();
 sg13g2_decap_8 FILLER_75_2077 ();
 sg13g2_decap_4 FILLER_75_2084 ();
 sg13g2_fill_2 FILLER_75_2088 ();
 sg13g2_fill_1 FILLER_75_2133 ();
 sg13g2_decap_4 FILLER_75_2157 ();
 sg13g2_fill_2 FILLER_75_2161 ();
 sg13g2_decap_4 FILLER_75_2171 ();
 sg13g2_fill_1 FILLER_75_2179 ();
 sg13g2_fill_1 FILLER_75_2186 ();
 sg13g2_decap_8 FILLER_75_2205 ();
 sg13g2_fill_1 FILLER_75_2212 ();
 sg13g2_fill_1 FILLER_75_2334 ();
 sg13g2_fill_1 FILLER_75_2339 ();
 sg13g2_fill_2 FILLER_75_2350 ();
 sg13g2_fill_2 FILLER_75_2378 ();
 sg13g2_decap_8 FILLER_75_2414 ();
 sg13g2_decap_4 FILLER_75_2421 ();
 sg13g2_fill_1 FILLER_75_2425 ();
 sg13g2_decap_4 FILLER_75_2462 ();
 sg13g2_decap_4 FILLER_75_2472 ();
 sg13g2_fill_2 FILLER_75_2476 ();
 sg13g2_decap_8 FILLER_75_2488 ();
 sg13g2_decap_8 FILLER_75_2495 ();
 sg13g2_decap_8 FILLER_75_2502 ();
 sg13g2_decap_8 FILLER_75_2509 ();
 sg13g2_decap_8 FILLER_75_2516 ();
 sg13g2_decap_4 FILLER_75_2523 ();
 sg13g2_fill_2 FILLER_75_2527 ();
 sg13g2_fill_2 FILLER_75_2533 ();
 sg13g2_fill_1 FILLER_75_2535 ();
 sg13g2_fill_2 FILLER_75_2540 ();
 sg13g2_decap_8 FILLER_75_2556 ();
 sg13g2_decap_8 FILLER_75_2563 ();
 sg13g2_decap_4 FILLER_75_2585 ();
 sg13g2_fill_1 FILLER_75_2589 ();
 sg13g2_decap_8 FILLER_75_2616 ();
 sg13g2_decap_8 FILLER_75_2623 ();
 sg13g2_decap_8 FILLER_75_2630 ();
 sg13g2_decap_8 FILLER_75_2637 ();
 sg13g2_decap_8 FILLER_75_2644 ();
 sg13g2_decap_8 FILLER_75_2651 ();
 sg13g2_decap_8 FILLER_75_2658 ();
 sg13g2_decap_4 FILLER_75_2665 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_102 ();
 sg13g2_fill_1 FILLER_76_129 ();
 sg13g2_fill_1 FILLER_76_135 ();
 sg13g2_decap_4 FILLER_76_156 ();
 sg13g2_fill_2 FILLER_76_160 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_183 ();
 sg13g2_fill_1 FILLER_76_185 ();
 sg13g2_fill_2 FILLER_76_191 ();
 sg13g2_fill_1 FILLER_76_193 ();
 sg13g2_decap_4 FILLER_76_204 ();
 sg13g2_fill_1 FILLER_76_208 ();
 sg13g2_decap_8 FILLER_76_212 ();
 sg13g2_decap_8 FILLER_76_219 ();
 sg13g2_fill_2 FILLER_76_226 ();
 sg13g2_fill_1 FILLER_76_231 ();
 sg13g2_decap_4 FILLER_76_258 ();
 sg13g2_fill_1 FILLER_76_271 ();
 sg13g2_decap_8 FILLER_76_275 ();
 sg13g2_decap_4 FILLER_76_282 ();
 sg13g2_decap_4 FILLER_76_291 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_decap_4 FILLER_76_306 ();
 sg13g2_fill_1 FILLER_76_310 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_fill_2 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_328 ();
 sg13g2_fill_1 FILLER_76_335 ();
 sg13g2_decap_4 FILLER_76_345 ();
 sg13g2_decap_4 FILLER_76_354 ();
 sg13g2_fill_1 FILLER_76_358 ();
 sg13g2_fill_2 FILLER_76_363 ();
 sg13g2_fill_1 FILLER_76_365 ();
 sg13g2_decap_4 FILLER_76_376 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_1 FILLER_76_391 ();
 sg13g2_fill_2 FILLER_76_397 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_409 ();
 sg13g2_fill_2 FILLER_76_468 ();
 sg13g2_fill_2 FILLER_76_473 ();
 sg13g2_decap_4 FILLER_76_506 ();
 sg13g2_fill_2 FILLER_76_510 ();
 sg13g2_fill_2 FILLER_76_565 ();
 sg13g2_fill_2 FILLER_76_633 ();
 sg13g2_fill_2 FILLER_76_659 ();
 sg13g2_decap_4 FILLER_76_671 ();
 sg13g2_fill_2 FILLER_76_675 ();
 sg13g2_fill_1 FILLER_76_692 ();
 sg13g2_fill_2 FILLER_76_697 ();
 sg13g2_fill_1 FILLER_76_699 ();
 sg13g2_fill_2 FILLER_76_709 ();
 sg13g2_fill_2 FILLER_76_796 ();
 sg13g2_decap_4 FILLER_76_852 ();
 sg13g2_decap_8 FILLER_76_882 ();
 sg13g2_decap_8 FILLER_76_889 ();
 sg13g2_decap_4 FILLER_76_896 ();
 sg13g2_decap_8 FILLER_76_926 ();
 sg13g2_decap_8 FILLER_76_943 ();
 sg13g2_fill_1 FILLER_76_950 ();
 sg13g2_fill_2 FILLER_76_957 ();
 sg13g2_fill_1 FILLER_76_959 ();
 sg13g2_fill_1 FILLER_76_974 ();
 sg13g2_fill_1 FILLER_76_987 ();
 sg13g2_fill_1 FILLER_76_993 ();
 sg13g2_fill_1 FILLER_76_998 ();
 sg13g2_fill_1 FILLER_76_1009 ();
 sg13g2_fill_1 FILLER_76_1020 ();
 sg13g2_fill_1 FILLER_76_1026 ();
 sg13g2_fill_1 FILLER_76_1031 ();
 sg13g2_decap_8 FILLER_76_1074 ();
 sg13g2_decap_8 FILLER_76_1081 ();
 sg13g2_decap_8 FILLER_76_1088 ();
 sg13g2_decap_8 FILLER_76_1095 ();
 sg13g2_decap_8 FILLER_76_1102 ();
 sg13g2_decap_8 FILLER_76_1109 ();
 sg13g2_decap_8 FILLER_76_1116 ();
 sg13g2_fill_2 FILLER_76_1137 ();
 sg13g2_fill_1 FILLER_76_1139 ();
 sg13g2_decap_8 FILLER_76_1166 ();
 sg13g2_decap_8 FILLER_76_1173 ();
 sg13g2_fill_2 FILLER_76_1180 ();
 sg13g2_fill_1 FILLER_76_1186 ();
 sg13g2_decap_8 FILLER_76_1190 ();
 sg13g2_fill_1 FILLER_76_1197 ();
 sg13g2_decap_8 FILLER_76_1227 ();
 sg13g2_fill_1 FILLER_76_1234 ();
 sg13g2_fill_2 FILLER_76_1242 ();
 sg13g2_fill_2 FILLER_76_1303 ();
 sg13g2_decap_4 FILLER_76_1329 ();
 sg13g2_fill_1 FILLER_76_1343 ();
 sg13g2_fill_2 FILLER_76_1358 ();
 sg13g2_decap_8 FILLER_76_1370 ();
 sg13g2_decap_8 FILLER_76_1377 ();
 sg13g2_decap_8 FILLER_76_1384 ();
 sg13g2_decap_8 FILLER_76_1391 ();
 sg13g2_fill_2 FILLER_76_1398 ();
 sg13g2_fill_2 FILLER_76_1410 ();
 sg13g2_fill_1 FILLER_76_1416 ();
 sg13g2_fill_1 FILLER_76_1444 ();
 sg13g2_decap_8 FILLER_76_1449 ();
 sg13g2_decap_8 FILLER_76_1456 ();
 sg13g2_decap_8 FILLER_76_1463 ();
 sg13g2_fill_2 FILLER_76_1470 ();
 sg13g2_fill_1 FILLER_76_1472 ();
 sg13g2_decap_4 FILLER_76_1479 ();
 sg13g2_fill_2 FILLER_76_1483 ();
 sg13g2_fill_1 FILLER_76_1489 ();
 sg13g2_fill_2 FILLER_76_1521 ();
 sg13g2_fill_2 FILLER_76_1528 ();
 sg13g2_fill_1 FILLER_76_1535 ();
 sg13g2_fill_1 FILLER_76_1541 ();
 sg13g2_fill_1 FILLER_76_1546 ();
 sg13g2_fill_1 FILLER_76_1552 ();
 sg13g2_fill_1 FILLER_76_1571 ();
 sg13g2_decap_8 FILLER_76_1624 ();
 sg13g2_fill_1 FILLER_76_1631 ();
 sg13g2_fill_1 FILLER_76_1637 ();
 sg13g2_fill_1 FILLER_76_1675 ();
 sg13g2_fill_1 FILLER_76_1684 ();
 sg13g2_fill_1 FILLER_76_1692 ();
 sg13g2_fill_1 FILLER_76_1715 ();
 sg13g2_fill_1 FILLER_76_1750 ();
 sg13g2_fill_2 FILLER_76_1755 ();
 sg13g2_decap_8 FILLER_76_1771 ();
 sg13g2_decap_8 FILLER_76_1778 ();
 sg13g2_decap_4 FILLER_76_1785 ();
 sg13g2_fill_1 FILLER_76_1789 ();
 sg13g2_decap_4 FILLER_76_1793 ();
 sg13g2_fill_1 FILLER_76_1797 ();
 sg13g2_fill_2 FILLER_76_1813 ();
 sg13g2_fill_2 FILLER_76_1829 ();
 sg13g2_fill_1 FILLER_76_1865 ();
 sg13g2_fill_2 FILLER_76_1879 ();
 sg13g2_fill_2 FILLER_76_1915 ();
 sg13g2_fill_1 FILLER_76_1917 ();
 sg13g2_fill_2 FILLER_76_1927 ();
 sg13g2_fill_1 FILLER_76_1933 ();
 sg13g2_fill_1 FILLER_76_1960 ();
 sg13g2_fill_1 FILLER_76_1965 ();
 sg13g2_fill_1 FILLER_76_1975 ();
 sg13g2_decap_8 FILLER_76_1988 ();
 sg13g2_fill_2 FILLER_76_1995 ();
 sg13g2_fill_2 FILLER_76_2005 ();
 sg13g2_fill_1 FILLER_76_2007 ();
 sg13g2_fill_2 FILLER_76_2018 ();
 sg13g2_decap_8 FILLER_76_2024 ();
 sg13g2_decap_8 FILLER_76_2035 ();
 sg13g2_decap_8 FILLER_76_2042 ();
 sg13g2_decap_8 FILLER_76_2049 ();
 sg13g2_decap_8 FILLER_76_2056 ();
 sg13g2_decap_8 FILLER_76_2063 ();
 sg13g2_decap_8 FILLER_76_2070 ();
 sg13g2_decap_8 FILLER_76_2077 ();
 sg13g2_decap_4 FILLER_76_2084 ();
 sg13g2_fill_2 FILLER_76_2088 ();
 sg13g2_decap_8 FILLER_76_2100 ();
 sg13g2_fill_2 FILLER_76_2107 ();
 sg13g2_fill_2 FILLER_76_2113 ();
 sg13g2_decap_4 FILLER_76_2125 ();
 sg13g2_fill_2 FILLER_76_2129 ();
 sg13g2_fill_1 FILLER_76_2144 ();
 sg13g2_decap_8 FILLER_76_2154 ();
 sg13g2_fill_1 FILLER_76_2187 ();
 sg13g2_fill_2 FILLER_76_2192 ();
 sg13g2_fill_2 FILLER_76_2204 ();
 sg13g2_fill_1 FILLER_76_2206 ();
 sg13g2_fill_1 FILLER_76_2232 ();
 sg13g2_fill_2 FILLER_76_2246 ();
 sg13g2_fill_2 FILLER_76_2264 ();
 sg13g2_fill_1 FILLER_76_2271 ();
 sg13g2_fill_2 FILLER_76_2357 ();
 sg13g2_fill_2 FILLER_76_2376 ();
 sg13g2_decap_8 FILLER_76_2414 ();
 sg13g2_decap_8 FILLER_76_2421 ();
 sg13g2_fill_1 FILLER_76_2460 ();
 sg13g2_fill_1 FILLER_76_2471 ();
 sg13g2_decap_4 FILLER_76_2478 ();
 sg13g2_fill_2 FILLER_76_2482 ();
 sg13g2_fill_1 FILLER_76_2494 ();
 sg13g2_fill_1 FILLER_76_2545 ();
 sg13g2_fill_1 FILLER_76_2556 ();
 sg13g2_fill_2 FILLER_76_2605 ();
 sg13g2_decap_8 FILLER_76_2612 ();
 sg13g2_decap_8 FILLER_76_2619 ();
 sg13g2_decap_8 FILLER_76_2626 ();
 sg13g2_decap_8 FILLER_76_2633 ();
 sg13g2_decap_8 FILLER_76_2640 ();
 sg13g2_decap_8 FILLER_76_2647 ();
 sg13g2_decap_8 FILLER_76_2654 ();
 sg13g2_decap_8 FILLER_76_2661 ();
 sg13g2_fill_2 FILLER_76_2668 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_4 FILLER_77_63 ();
 sg13g2_fill_2 FILLER_77_67 ();
 sg13g2_decap_8 FILLER_77_73 ();
 sg13g2_fill_2 FILLER_77_100 ();
 sg13g2_fill_1 FILLER_77_127 ();
 sg13g2_fill_2 FILLER_77_138 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_2 FILLER_77_200 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_decap_8 FILLER_77_303 ();
 sg13g2_decap_8 FILLER_77_310 ();
 sg13g2_decap_8 FILLER_77_317 ();
 sg13g2_fill_2 FILLER_77_324 ();
 sg13g2_fill_1 FILLER_77_326 ();
 sg13g2_fill_1 FILLER_77_367 ();
 sg13g2_fill_1 FILLER_77_394 ();
 sg13g2_fill_2 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_417 ();
 sg13g2_fill_1 FILLER_77_423 ();
 sg13g2_fill_1 FILLER_77_428 ();
 sg13g2_fill_1 FILLER_77_434 ();
 sg13g2_fill_1 FILLER_77_439 ();
 sg13g2_fill_2 FILLER_77_446 ();
 sg13g2_fill_2 FILLER_77_480 ();
 sg13g2_fill_2 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_496 ();
 sg13g2_decap_8 FILLER_77_503 ();
 sg13g2_fill_2 FILLER_77_510 ();
 sg13g2_fill_1 FILLER_77_526 ();
 sg13g2_fill_1 FILLER_77_599 ();
 sg13g2_fill_1 FILLER_77_610 ();
 sg13g2_fill_2 FILLER_77_689 ();
 sg13g2_fill_2 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_fill_1 FILLER_77_797 ();
 sg13g2_decap_4 FILLER_77_810 ();
 sg13g2_fill_1 FILLER_77_814 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_fill_2 FILLER_77_825 ();
 sg13g2_fill_2 FILLER_77_863 ();
 sg13g2_fill_1 FILLER_77_865 ();
 sg13g2_decap_8 FILLER_77_892 ();
 sg13g2_decap_4 FILLER_77_899 ();
 sg13g2_fill_2 FILLER_77_903 ();
 sg13g2_decap_8 FILLER_77_909 ();
 sg13g2_fill_2 FILLER_77_916 ();
 sg13g2_fill_1 FILLER_77_918 ();
 sg13g2_decap_8 FILLER_77_1005 ();
 sg13g2_fill_2 FILLER_77_1012 ();
 sg13g2_fill_1 FILLER_77_1040 ();
 sg13g2_fill_1 FILLER_77_1087 ();
 sg13g2_fill_2 FILLER_77_1124 ();
 sg13g2_decap_4 FILLER_77_1201 ();
 sg13g2_decap_4 FILLER_77_1209 ();
 sg13g2_fill_1 FILLER_77_1213 ();
 sg13g2_decap_8 FILLER_77_1240 ();
 sg13g2_decap_8 FILLER_77_1247 ();
 sg13g2_decap_8 FILLER_77_1254 ();
 sg13g2_fill_2 FILLER_77_1261 ();
 sg13g2_fill_2 FILLER_77_1267 ();
 sg13g2_fill_1 FILLER_77_1269 ();
 sg13g2_decap_4 FILLER_77_1296 ();
 sg13g2_fill_1 FILLER_77_1300 ();
 sg13g2_fill_1 FILLER_77_1327 ();
 sg13g2_decap_8 FILLER_77_1332 ();
 sg13g2_fill_2 FILLER_77_1339 ();
 sg13g2_fill_1 FILLER_77_1341 ();
 sg13g2_fill_2 FILLER_77_1382 ();
 sg13g2_fill_1 FILLER_77_1384 ();
 sg13g2_fill_1 FILLER_77_1399 ();
 sg13g2_decap_8 FILLER_77_1452 ();
 sg13g2_fill_1 FILLER_77_1459 ();
 sg13g2_fill_1 FILLER_77_1486 ();
 sg13g2_fill_2 FILLER_77_1492 ();
 sg13g2_fill_1 FILLER_77_1520 ();
 sg13g2_fill_2 FILLER_77_1552 ();
 sg13g2_fill_1 FILLER_77_1581 ();
 sg13g2_fill_2 FILLER_77_1589 ();
 sg13g2_fill_1 FILLER_77_1614 ();
 sg13g2_fill_2 FILLER_77_1677 ();
 sg13g2_fill_1 FILLER_77_1679 ();
 sg13g2_fill_2 FILLER_77_1708 ();
 sg13g2_decap_8 FILLER_77_1762 ();
 sg13g2_decap_8 FILLER_77_1769 ();
 sg13g2_decap_4 FILLER_77_1776 ();
 sg13g2_decap_8 FILLER_77_1783 ();
 sg13g2_fill_1 FILLER_77_1790 ();
 sg13g2_decap_4 FILLER_77_1796 ();
 sg13g2_fill_1 FILLER_77_1800 ();
 sg13g2_fill_2 FILLER_77_1809 ();
 sg13g2_fill_1 FILLER_77_1814 ();
 sg13g2_fill_2 FILLER_77_1827 ();
 sg13g2_fill_1 FILLER_77_1838 ();
 sg13g2_fill_1 FILLER_77_1856 ();
 sg13g2_fill_2 FILLER_77_1881 ();
 sg13g2_fill_1 FILLER_77_1883 ();
 sg13g2_fill_1 FILLER_77_1899 ();
 sg13g2_fill_2 FILLER_77_1930 ();
 sg13g2_fill_2 FILLER_77_1936 ();
 sg13g2_fill_2 FILLER_77_1964 ();
 sg13g2_fill_1 FILLER_77_1966 ();
 sg13g2_fill_2 FILLER_77_1980 ();
 sg13g2_fill_1 FILLER_77_1982 ();
 sg13g2_decap_8 FILLER_77_2009 ();
 sg13g2_decap_8 FILLER_77_2016 ();
 sg13g2_decap_8 FILLER_77_2023 ();
 sg13g2_decap_8 FILLER_77_2030 ();
 sg13g2_decap_8 FILLER_77_2037 ();
 sg13g2_decap_8 FILLER_77_2044 ();
 sg13g2_decap_8 FILLER_77_2051 ();
 sg13g2_decap_8 FILLER_77_2058 ();
 sg13g2_decap_8 FILLER_77_2065 ();
 sg13g2_decap_8 FILLER_77_2072 ();
 sg13g2_decap_4 FILLER_77_2079 ();
 sg13g2_fill_2 FILLER_77_2083 ();
 sg13g2_decap_8 FILLER_77_2111 ();
 sg13g2_fill_2 FILLER_77_2118 ();
 sg13g2_decap_8 FILLER_77_2130 ();
 sg13g2_fill_1 FILLER_77_2169 ();
 sg13g2_fill_1 FILLER_77_2180 ();
 sg13g2_fill_1 FILLER_77_2187 ();
 sg13g2_fill_1 FILLER_77_2198 ();
 sg13g2_fill_1 FILLER_77_2231 ();
 sg13g2_fill_1 FILLER_77_2242 ();
 sg13g2_fill_1 FILLER_77_2287 ();
 sg13g2_fill_2 FILLER_77_2349 ();
 sg13g2_fill_2 FILLER_77_2435 ();
 sg13g2_decap_8 FILLER_77_2441 ();
 sg13g2_fill_2 FILLER_77_2484 ();
 sg13g2_decap_8 FILLER_77_2520 ();
 sg13g2_fill_1 FILLER_77_2527 ();
 sg13g2_fill_2 FILLER_77_2541 ();
 sg13g2_decap_8 FILLER_77_2603 ();
 sg13g2_decap_8 FILLER_77_2610 ();
 sg13g2_decap_8 FILLER_77_2617 ();
 sg13g2_decap_8 FILLER_77_2624 ();
 sg13g2_decap_8 FILLER_77_2631 ();
 sg13g2_decap_8 FILLER_77_2638 ();
 sg13g2_decap_8 FILLER_77_2645 ();
 sg13g2_decap_8 FILLER_77_2652 ();
 sg13g2_decap_8 FILLER_77_2659 ();
 sg13g2_decap_4 FILLER_77_2666 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_81 ();
 sg13g2_fill_1 FILLER_78_108 ();
 sg13g2_fill_1 FILLER_78_114 ();
 sg13g2_fill_1 FILLER_78_155 ();
 sg13g2_fill_1 FILLER_78_272 ();
 sg13g2_fill_1 FILLER_78_278 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_fill_2 FILLER_78_322 ();
 sg13g2_decap_4 FILLER_78_355 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_fill_1 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_428 ();
 sg13g2_fill_1 FILLER_78_434 ();
 sg13g2_fill_1 FILLER_78_440 ();
 sg13g2_fill_2 FILLER_78_467 ();
 sg13g2_fill_1 FILLER_78_479 ();
 sg13g2_fill_2 FILLER_78_510 ();
 sg13g2_fill_1 FILLER_78_512 ();
 sg13g2_fill_1 FILLER_78_586 ();
 sg13g2_fill_1 FILLER_78_592 ();
 sg13g2_fill_1 FILLER_78_597 ();
 sg13g2_fill_1 FILLER_78_629 ();
 sg13g2_fill_1 FILLER_78_635 ();
 sg13g2_fill_2 FILLER_78_665 ();
 sg13g2_fill_2 FILLER_78_673 ();
 sg13g2_decap_4 FILLER_78_684 ();
 sg13g2_fill_2 FILLER_78_688 ();
 sg13g2_fill_2 FILLER_78_751 ();
 sg13g2_decap_8 FILLER_78_800 ();
 sg13g2_decap_4 FILLER_78_807 ();
 sg13g2_fill_1 FILLER_78_811 ();
 sg13g2_fill_2 FILLER_78_872 ();
 sg13g2_fill_1 FILLER_78_874 ();
 sg13g2_decap_8 FILLER_78_884 ();
 sg13g2_decap_8 FILLER_78_891 ();
 sg13g2_decap_8 FILLER_78_898 ();
 sg13g2_decap_4 FILLER_78_905 ();
 sg13g2_fill_1 FILLER_78_961 ();
 sg13g2_fill_1 FILLER_78_1028 ();
 sg13g2_fill_2 FILLER_78_1055 ();
 sg13g2_fill_2 FILLER_78_1088 ();
 sg13g2_fill_1 FILLER_78_1090 ();
 sg13g2_fill_1 FILLER_78_1127 ();
 sg13g2_fill_2 FILLER_78_1162 ();
 sg13g2_fill_1 FILLER_78_1164 ();
 sg13g2_fill_2 FILLER_78_1195 ();
 sg13g2_fill_1 FILLER_78_1197 ();
 sg13g2_fill_2 FILLER_78_1244 ();
 sg13g2_fill_1 FILLER_78_1246 ();
 sg13g2_decap_4 FILLER_78_1260 ();
 sg13g2_fill_2 FILLER_78_1264 ();
 sg13g2_fill_2 FILLER_78_1312 ();
 sg13g2_fill_1 FILLER_78_1314 ();
 sg13g2_fill_1 FILLER_78_1367 ();
 sg13g2_decap_8 FILLER_78_1420 ();
 sg13g2_decap_4 FILLER_78_1427 ();
 sg13g2_fill_2 FILLER_78_1431 ();
 sg13g2_decap_8 FILLER_78_1437 ();
 sg13g2_fill_2 FILLER_78_1444 ();
 sg13g2_fill_1 FILLER_78_1450 ();
 sg13g2_fill_2 FILLER_78_1498 ();
 sg13g2_fill_1 FILLER_78_1505 ();
 sg13g2_decap_4 FILLER_78_1552 ();
 sg13g2_fill_1 FILLER_78_1591 ();
 sg13g2_fill_1 FILLER_78_1596 ();
 sg13g2_decap_4 FILLER_78_1629 ();
 sg13g2_fill_1 FILLER_78_1648 ();
 sg13g2_fill_2 FILLER_78_1653 ();
 sg13g2_fill_1 FILLER_78_1676 ();
 sg13g2_fill_1 FILLER_78_1682 ();
 sg13g2_fill_1 FILLER_78_1688 ();
 sg13g2_fill_2 FILLER_78_1694 ();
 sg13g2_fill_2 FILLER_78_1701 ();
 sg13g2_fill_1 FILLER_78_1734 ();
 sg13g2_fill_1 FILLER_78_1741 ();
 sg13g2_fill_1 FILLER_78_1746 ();
 sg13g2_fill_2 FILLER_78_1760 ();
 sg13g2_fill_2 FILLER_78_1765 ();
 sg13g2_fill_1 FILLER_78_1767 ();
 sg13g2_decap_8 FILLER_78_1776 ();
 sg13g2_decap_8 FILLER_78_1783 ();
 sg13g2_fill_2 FILLER_78_1790 ();
 sg13g2_fill_1 FILLER_78_1792 ();
 sg13g2_fill_2 FILLER_78_1797 ();
 sg13g2_fill_2 FILLER_78_1807 ();
 sg13g2_fill_1 FILLER_78_1809 ();
 sg13g2_fill_2 FILLER_78_1828 ();
 sg13g2_fill_1 FILLER_78_1842 ();
 sg13g2_fill_2 FILLER_78_1852 ();
 sg13g2_fill_1 FILLER_78_1881 ();
 sg13g2_fill_1 FILLER_78_1917 ();
 sg13g2_fill_2 FILLER_78_1927 ();
 sg13g2_fill_1 FILLER_78_1929 ();
 sg13g2_fill_1 FILLER_78_1956 ();
 sg13g2_fill_1 FILLER_78_1975 ();
 sg13g2_decap_8 FILLER_78_2012 ();
 sg13g2_decap_8 FILLER_78_2019 ();
 sg13g2_decap_8 FILLER_78_2026 ();
 sg13g2_decap_8 FILLER_78_2033 ();
 sg13g2_decap_8 FILLER_78_2040 ();
 sg13g2_decap_8 FILLER_78_2047 ();
 sg13g2_decap_8 FILLER_78_2054 ();
 sg13g2_decap_8 FILLER_78_2061 ();
 sg13g2_decap_8 FILLER_78_2068 ();
 sg13g2_decap_4 FILLER_78_2075 ();
 sg13g2_fill_1 FILLER_78_2079 ();
 sg13g2_fill_2 FILLER_78_2084 ();
 sg13g2_fill_1 FILLER_78_2086 ();
 sg13g2_fill_1 FILLER_78_2177 ();
 sg13g2_fill_1 FILLER_78_2188 ();
 sg13g2_fill_1 FILLER_78_2215 ();
 sg13g2_fill_2 FILLER_78_2282 ();
 sg13g2_decap_4 FILLER_78_2410 ();
 sg13g2_fill_2 FILLER_78_2414 ();
 sg13g2_decap_8 FILLER_78_2442 ();
 sg13g2_decap_4 FILLER_78_2449 ();
 sg13g2_fill_2 FILLER_78_2483 ();
 sg13g2_fill_1 FILLER_78_2485 ();
 sg13g2_fill_1 FILLER_78_2522 ();
 sg13g2_fill_2 FILLER_78_2559 ();
 sg13g2_fill_1 FILLER_78_2561 ();
 sg13g2_fill_2 FILLER_78_2572 ();
 sg13g2_fill_1 FILLER_78_2574 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_8 FILLER_78_2586 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_fill_1 FILLER_79_85 ();
 sg13g2_fill_1 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_117 ();
 sg13g2_fill_1 FILLER_79_128 ();
 sg13g2_fill_1 FILLER_79_210 ();
 sg13g2_fill_1 FILLER_79_225 ();
 sg13g2_fill_1 FILLER_79_263 ();
 sg13g2_decap_8 FILLER_79_306 ();
 sg13g2_decap_8 FILLER_79_313 ();
 sg13g2_decap_8 FILLER_79_320 ();
 sg13g2_decap_4 FILLER_79_327 ();
 sg13g2_fill_2 FILLER_79_335 ();
 sg13g2_fill_1 FILLER_79_337 ();
 sg13g2_fill_2 FILLER_79_343 ();
 sg13g2_fill_1 FILLER_79_345 ();
 sg13g2_fill_2 FILLER_79_372 ();
 sg13g2_fill_2 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_4 FILLER_79_391 ();
 sg13g2_fill_2 FILLER_79_445 ();
 sg13g2_decap_4 FILLER_79_459 ();
 sg13g2_fill_1 FILLER_79_463 ();
 sg13g2_fill_2 FILLER_79_470 ();
 sg13g2_decap_8 FILLER_79_498 ();
 sg13g2_decap_4 FILLER_79_505 ();
 sg13g2_fill_2 FILLER_79_509 ();
 sg13g2_decap_4 FILLER_79_623 ();
 sg13g2_fill_2 FILLER_79_670 ();
 sg13g2_fill_1 FILLER_79_712 ();
 sg13g2_fill_2 FILLER_79_718 ();
 sg13g2_fill_2 FILLER_79_762 ();
 sg13g2_fill_1 FILLER_79_764 ();
 sg13g2_fill_2 FILLER_79_773 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_831 ();
 sg13g2_decap_4 FILLER_79_838 ();
 sg13g2_decap_8 FILLER_79_864 ();
 sg13g2_decap_8 FILLER_79_871 ();
 sg13g2_decap_8 FILLER_79_878 ();
 sg13g2_decap_8 FILLER_79_885 ();
 sg13g2_decap_8 FILLER_79_892 ();
 sg13g2_decap_8 FILLER_79_899 ();
 sg13g2_fill_1 FILLER_79_906 ();
 sg13g2_decap_4 FILLER_79_954 ();
 sg13g2_fill_2 FILLER_79_968 ();
 sg13g2_fill_1 FILLER_79_970 ();
 sg13g2_decap_8 FILLER_79_975 ();
 sg13g2_fill_1 FILLER_79_992 ();
 sg13g2_fill_2 FILLER_79_1019 ();
 sg13g2_decap_4 FILLER_79_1045 ();
 sg13g2_fill_2 FILLER_79_1049 ();
 sg13g2_decap_8 FILLER_79_1078 ();
 sg13g2_decap_8 FILLER_79_1085 ();
 sg13g2_decap_8 FILLER_79_1092 ();
 sg13g2_decap_4 FILLER_79_1099 ();
 sg13g2_fill_2 FILLER_79_1103 ();
 sg13g2_fill_1 FILLER_79_1109 ();
 sg13g2_decap_4 FILLER_79_1150 ();
 sg13g2_fill_2 FILLER_79_1167 ();
 sg13g2_fill_2 FILLER_79_1215 ();
 sg13g2_fill_2 FILLER_79_1263 ();
 sg13g2_fill_1 FILLER_79_1265 ();
 sg13g2_fill_2 FILLER_79_1292 ();
 sg13g2_fill_1 FILLER_79_1294 ();
 sg13g2_decap_4 FILLER_79_1325 ();
 sg13g2_fill_2 FILLER_79_1369 ();
 sg13g2_decap_8 FILLER_79_1427 ();
 sg13g2_decap_8 FILLER_79_1434 ();
 sg13g2_decap_8 FILLER_79_1441 ();
 sg13g2_decap_8 FILLER_79_1448 ();
 sg13g2_decap_8 FILLER_79_1455 ();
 sg13g2_fill_2 FILLER_79_1462 ();
 sg13g2_fill_2 FILLER_79_1468 ();
 sg13g2_fill_1 FILLER_79_1470 ();
 sg13g2_decap_8 FILLER_79_1474 ();
 sg13g2_decap_8 FILLER_79_1481 ();
 sg13g2_fill_1 FILLER_79_1496 ();
 sg13g2_fill_1 FILLER_79_1512 ();
 sg13g2_decap_4 FILLER_79_1517 ();
 sg13g2_fill_2 FILLER_79_1525 ();
 sg13g2_fill_1 FILLER_79_1527 ();
 sg13g2_fill_2 FILLER_79_1535 ();
 sg13g2_fill_1 FILLER_79_1569 ();
 sg13g2_fill_2 FILLER_79_1575 ();
 sg13g2_fill_1 FILLER_79_1577 ();
 sg13g2_fill_2 FILLER_79_1583 ();
 sg13g2_decap_4 FILLER_79_1589 ();
 sg13g2_decap_4 FILLER_79_1598 ();
 sg13g2_fill_1 FILLER_79_1602 ();
 sg13g2_decap_4 FILLER_79_1607 ();
 sg13g2_fill_1 FILLER_79_1611 ();
 sg13g2_decap_8 FILLER_79_1616 ();
 sg13g2_decap_8 FILLER_79_1623 ();
 sg13g2_fill_2 FILLER_79_1630 ();
 sg13g2_fill_1 FILLER_79_1632 ();
 sg13g2_fill_2 FILLER_79_1712 ();
 sg13g2_fill_1 FILLER_79_1714 ();
 sg13g2_decap_4 FILLER_79_1745 ();
 sg13g2_fill_1 FILLER_79_1749 ();
 sg13g2_decap_8 FILLER_79_1780 ();
 sg13g2_decap_8 FILLER_79_1787 ();
 sg13g2_decap_8 FILLER_79_1794 ();
 sg13g2_decap_8 FILLER_79_1801 ();
 sg13g2_decap_4 FILLER_79_1808 ();
 sg13g2_fill_2 FILLER_79_1812 ();
 sg13g2_fill_1 FILLER_79_1818 ();
 sg13g2_fill_2 FILLER_79_1824 ();
 sg13g2_fill_2 FILLER_79_1834 ();
 sg13g2_fill_1 FILLER_79_1836 ();
 sg13g2_fill_1 FILLER_79_1881 ();
 sg13g2_fill_1 FILLER_79_1901 ();
 sg13g2_decap_4 FILLER_79_1907 ();
 sg13g2_fill_2 FILLER_79_1911 ();
 sg13g2_fill_2 FILLER_79_1939 ();
 sg13g2_fill_2 FILLER_79_1945 ();
 sg13g2_fill_2 FILLER_79_1951 ();
 sg13g2_decap_4 FILLER_79_1957 ();
 sg13g2_fill_1 FILLER_79_1961 ();
 sg13g2_decap_4 FILLER_79_1988 ();
 sg13g2_fill_1 FILLER_79_1992 ();
 sg13g2_decap_8 FILLER_79_1997 ();
 sg13g2_decap_8 FILLER_79_2004 ();
 sg13g2_decap_8 FILLER_79_2011 ();
 sg13g2_decap_8 FILLER_79_2018 ();
 sg13g2_decap_8 FILLER_79_2025 ();
 sg13g2_decap_8 FILLER_79_2032 ();
 sg13g2_decap_8 FILLER_79_2039 ();
 sg13g2_decap_8 FILLER_79_2046 ();
 sg13g2_decap_8 FILLER_79_2053 ();
 sg13g2_decap_8 FILLER_79_2060 ();
 sg13g2_decap_8 FILLER_79_2067 ();
 sg13g2_decap_4 FILLER_79_2100 ();
 sg13g2_fill_1 FILLER_79_2104 ();
 sg13g2_fill_1 FILLER_79_2109 ();
 sg13g2_fill_1 FILLER_79_2114 ();
 sg13g2_fill_1 FILLER_79_2155 ();
 sg13g2_decap_8 FILLER_79_2160 ();
 sg13g2_decap_4 FILLER_79_2167 ();
 sg13g2_fill_2 FILLER_79_2176 ();
 sg13g2_fill_2 FILLER_79_2217 ();
 sg13g2_fill_1 FILLER_79_2245 ();
 sg13g2_fill_1 FILLER_79_2282 ();
 sg13g2_fill_1 FILLER_79_2288 ();
 sg13g2_fill_1 FILLER_79_2293 ();
 sg13g2_fill_2 FILLER_79_2320 ();
 sg13g2_fill_1 FILLER_79_2348 ();
 sg13g2_fill_1 FILLER_79_2375 ();
 sg13g2_decap_4 FILLER_79_2415 ();
 sg13g2_fill_1 FILLER_79_2419 ();
 sg13g2_decap_4 FILLER_79_2472 ();
 sg13g2_fill_1 FILLER_79_2480 ();
 sg13g2_decap_8 FILLER_79_2517 ();
 sg13g2_decap_4 FILLER_79_2524 ();
 sg13g2_fill_2 FILLER_79_2528 ();
 sg13g2_decap_8 FILLER_79_2534 ();
 sg13g2_decap_8 FILLER_79_2541 ();
 sg13g2_decap_8 FILLER_79_2574 ();
 sg13g2_decap_8 FILLER_79_2581 ();
 sg13g2_decap_8 FILLER_79_2588 ();
 sg13g2_decap_8 FILLER_79_2595 ();
 sg13g2_decap_8 FILLER_79_2602 ();
 sg13g2_decap_8 FILLER_79_2609 ();
 sg13g2_decap_8 FILLER_79_2616 ();
 sg13g2_decap_8 FILLER_79_2623 ();
 sg13g2_decap_8 FILLER_79_2630 ();
 sg13g2_decap_8 FILLER_79_2637 ();
 sg13g2_decap_8 FILLER_79_2644 ();
 sg13g2_decap_8 FILLER_79_2651 ();
 sg13g2_decap_8 FILLER_79_2658 ();
 sg13g2_decap_4 FILLER_79_2665 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_fill_1 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_89 ();
 sg13g2_fill_2 FILLER_80_95 ();
 sg13g2_fill_2 FILLER_80_101 ();
 sg13g2_fill_2 FILLER_80_121 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_143 ();
 sg13g2_fill_1 FILLER_80_163 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_182 ();
 sg13g2_fill_2 FILLER_80_195 ();
 sg13g2_fill_1 FILLER_80_197 ();
 sg13g2_decap_4 FILLER_80_206 ();
 sg13g2_fill_1 FILLER_80_210 ();
 sg13g2_decap_4 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_223 ();
 sg13g2_fill_1 FILLER_80_225 ();
 sg13g2_fill_1 FILLER_80_259 ();
 sg13g2_fill_1 FILLER_80_269 ();
 sg13g2_fill_2 FILLER_80_279 ();
 sg13g2_fill_1 FILLER_80_281 ();
 sg13g2_fill_2 FILLER_80_291 ();
 sg13g2_fill_1 FILLER_80_293 ();
 sg13g2_decap_4 FILLER_80_313 ();
 sg13g2_fill_1 FILLER_80_317 ();
 sg13g2_fill_2 FILLER_80_333 ();
 sg13g2_fill_2 FILLER_80_340 ();
 sg13g2_fill_2 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_363 ();
 sg13g2_decap_8 FILLER_80_370 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_fill_1 FILLER_80_379 ();
 sg13g2_fill_1 FILLER_80_417 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_fill_2 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_fill_1 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_497 ();
 sg13g2_decap_8 FILLER_80_504 ();
 sg13g2_decap_4 FILLER_80_511 ();
 sg13g2_fill_2 FILLER_80_515 ();
 sg13g2_fill_2 FILLER_80_529 ();
 sg13g2_decap_4 FILLER_80_535 ();
 sg13g2_fill_2 FILLER_80_545 ();
 sg13g2_fill_1 FILLER_80_584 ();
 sg13g2_fill_2 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_fill_1 FILLER_80_630 ();
 sg13g2_fill_2 FILLER_80_638 ();
 sg13g2_fill_2 FILLER_80_684 ();
 sg13g2_decap_4 FILLER_80_722 ();
 sg13g2_fill_1 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_fill_1 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_4 FILLER_80_826 ();
 sg13g2_fill_1 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_fill_1 FILLER_80_917 ();
 sg13g2_decap_4 FILLER_80_922 ();
 sg13g2_decap_8 FILLER_80_930 ();
 sg13g2_decap_8 FILLER_80_937 ();
 sg13g2_decap_8 FILLER_80_944 ();
 sg13g2_decap_8 FILLER_80_951 ();
 sg13g2_decap_8 FILLER_80_958 ();
 sg13g2_decap_8 FILLER_80_965 ();
 sg13g2_decap_8 FILLER_80_972 ();
 sg13g2_decap_8 FILLER_80_979 ();
 sg13g2_decap_8 FILLER_80_986 ();
 sg13g2_decap_4 FILLER_80_993 ();
 sg13g2_fill_1 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1006 ();
 sg13g2_decap_8 FILLER_80_1013 ();
 sg13g2_decap_8 FILLER_80_1020 ();
 sg13g2_decap_8 FILLER_80_1027 ();
 sg13g2_decap_4 FILLER_80_1034 ();
 sg13g2_fill_1 FILLER_80_1038 ();
 sg13g2_decap_8 FILLER_80_1073 ();
 sg13g2_decap_8 FILLER_80_1080 ();
 sg13g2_decap_8 FILLER_80_1087 ();
 sg13g2_decap_8 FILLER_80_1094 ();
 sg13g2_decap_8 FILLER_80_1101 ();
 sg13g2_decap_8 FILLER_80_1108 ();
 sg13g2_decap_8 FILLER_80_1115 ();
 sg13g2_decap_8 FILLER_80_1122 ();
 sg13g2_decap_4 FILLER_80_1129 ();
 sg13g2_decap_8 FILLER_80_1141 ();
 sg13g2_decap_8 FILLER_80_1148 ();
 sg13g2_decap_8 FILLER_80_1155 ();
 sg13g2_fill_2 FILLER_80_1162 ();
 sg13g2_fill_1 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_4 FILLER_80_1194 ();
 sg13g2_fill_2 FILLER_80_1227 ();
 sg13g2_fill_1 FILLER_80_1233 ();
 sg13g2_fill_2 FILLER_80_1242 ();
 sg13g2_decap_8 FILLER_80_1260 ();
 sg13g2_decap_4 FILLER_80_1267 ();
 sg13g2_fill_1 FILLER_80_1271 ();
 sg13g2_fill_1 FILLER_80_1276 ();
 sg13g2_fill_1 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1286 ();
 sg13g2_decap_8 FILLER_80_1293 ();
 sg13g2_fill_2 FILLER_80_1300 ();
 sg13g2_decap_4 FILLER_80_1306 ();
 sg13g2_decap_8 FILLER_80_1314 ();
 sg13g2_decap_8 FILLER_80_1321 ();
 sg13g2_decap_8 FILLER_80_1328 ();
 sg13g2_fill_2 FILLER_80_1335 ();
 sg13g2_decap_4 FILLER_80_1341 ();
 sg13g2_decap_8 FILLER_80_1349 ();
 sg13g2_decap_8 FILLER_80_1356 ();
 sg13g2_decap_8 FILLER_80_1363 ();
 sg13g2_decap_8 FILLER_80_1370 ();
 sg13g2_decap_8 FILLER_80_1377 ();
 sg13g2_fill_1 FILLER_80_1384 ();
 sg13g2_decap_8 FILLER_80_1389 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_fill_1 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1440 ();
 sg13g2_decap_8 FILLER_80_1447 ();
 sg13g2_decap_8 FILLER_80_1454 ();
 sg13g2_decap_8 FILLER_80_1461 ();
 sg13g2_decap_8 FILLER_80_1468 ();
 sg13g2_decap_8 FILLER_80_1475 ();
 sg13g2_decap_8 FILLER_80_1482 ();
 sg13g2_decap_4 FILLER_80_1489 ();
 sg13g2_fill_1 FILLER_80_1493 ();
 sg13g2_decap_8 FILLER_80_1498 ();
 sg13g2_decap_8 FILLER_80_1505 ();
 sg13g2_decap_8 FILLER_80_1512 ();
 sg13g2_decap_8 FILLER_80_1519 ();
 sg13g2_fill_2 FILLER_80_1526 ();
 sg13g2_fill_1 FILLER_80_1565 ();
 sg13g2_decap_8 FILLER_80_1570 ();
 sg13g2_decap_8 FILLER_80_1577 ();
 sg13g2_decap_8 FILLER_80_1584 ();
 sg13g2_decap_8 FILLER_80_1591 ();
 sg13g2_decap_8 FILLER_80_1598 ();
 sg13g2_decap_8 FILLER_80_1605 ();
 sg13g2_decap_8 FILLER_80_1612 ();
 sg13g2_decap_8 FILLER_80_1619 ();
 sg13g2_decap_8 FILLER_80_1626 ();
 sg13g2_decap_8 FILLER_80_1633 ();
 sg13g2_decap_8 FILLER_80_1640 ();
 sg13g2_fill_2 FILLER_80_1647 ();
 sg13g2_fill_1 FILLER_80_1649 ();
 sg13g2_decap_4 FILLER_80_1654 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_4 FILLER_80_1677 ();
 sg13g2_fill_1 FILLER_80_1681 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_4 FILLER_80_1711 ();
 sg13g2_decap_4 FILLER_80_1719 ();
 sg13g2_fill_2 FILLER_80_1723 ();
 sg13g2_decap_8 FILLER_80_1729 ();
 sg13g2_fill_2 FILLER_80_1736 ();
 sg13g2_decap_8 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1749 ();
 sg13g2_decap_4 FILLER_80_1756 ();
 sg13g2_fill_2 FILLER_80_1760 ();
 sg13g2_decap_8 FILLER_80_1766 ();
 sg13g2_decap_8 FILLER_80_1773 ();
 sg13g2_decap_8 FILLER_80_1780 ();
 sg13g2_decap_8 FILLER_80_1787 ();
 sg13g2_decap_8 FILLER_80_1794 ();
 sg13g2_decap_8 FILLER_80_1801 ();
 sg13g2_decap_8 FILLER_80_1808 ();
 sg13g2_decap_8 FILLER_80_1815 ();
 sg13g2_decap_8 FILLER_80_1822 ();
 sg13g2_decap_8 FILLER_80_1829 ();
 sg13g2_decap_8 FILLER_80_1836 ();
 sg13g2_decap_8 FILLER_80_1843 ();
 sg13g2_fill_1 FILLER_80_1850 ();
 sg13g2_decap_8 FILLER_80_1863 ();
 sg13g2_decap_8 FILLER_80_1870 ();
 sg13g2_decap_8 FILLER_80_1877 ();
 sg13g2_decap_8 FILLER_80_1884 ();
 sg13g2_decap_8 FILLER_80_1891 ();
 sg13g2_decap_8 FILLER_80_1898 ();
 sg13g2_decap_8 FILLER_80_1905 ();
 sg13g2_decap_8 FILLER_80_1912 ();
 sg13g2_fill_1 FILLER_80_1919 ();
 sg13g2_decap_8 FILLER_80_1924 ();
 sg13g2_decap_8 FILLER_80_1931 ();
 sg13g2_decap_8 FILLER_80_1938 ();
 sg13g2_decap_8 FILLER_80_1945 ();
 sg13g2_decap_8 FILLER_80_1952 ();
 sg13g2_decap_8 FILLER_80_1959 ();
 sg13g2_fill_1 FILLER_80_1966 ();
 sg13g2_decap_8 FILLER_80_1975 ();
 sg13g2_decap_8 FILLER_80_1982 ();
 sg13g2_decap_8 FILLER_80_1989 ();
 sg13g2_decap_8 FILLER_80_1996 ();
 sg13g2_decap_8 FILLER_80_2003 ();
 sg13g2_decap_8 FILLER_80_2010 ();
 sg13g2_decap_8 FILLER_80_2017 ();
 sg13g2_decap_8 FILLER_80_2024 ();
 sg13g2_decap_8 FILLER_80_2031 ();
 sg13g2_decap_8 FILLER_80_2038 ();
 sg13g2_decap_8 FILLER_80_2045 ();
 sg13g2_decap_8 FILLER_80_2052 ();
 sg13g2_decap_8 FILLER_80_2059 ();
 sg13g2_decap_8 FILLER_80_2066 ();
 sg13g2_decap_8 FILLER_80_2073 ();
 sg13g2_decap_8 FILLER_80_2080 ();
 sg13g2_decap_8 FILLER_80_2087 ();
 sg13g2_decap_8 FILLER_80_2094 ();
 sg13g2_decap_8 FILLER_80_2101 ();
 sg13g2_decap_8 FILLER_80_2108 ();
 sg13g2_decap_4 FILLER_80_2115 ();
 sg13g2_fill_2 FILLER_80_2119 ();
 sg13g2_decap_8 FILLER_80_2125 ();
 sg13g2_decap_8 FILLER_80_2132 ();
 sg13g2_decap_8 FILLER_80_2139 ();
 sg13g2_fill_2 FILLER_80_2146 ();
 sg13g2_fill_1 FILLER_80_2148 ();
 sg13g2_fill_2 FILLER_80_2175 ();
 sg13g2_decap_8 FILLER_80_2191 ();
 sg13g2_fill_2 FILLER_80_2198 ();
 sg13g2_fill_1 FILLER_80_2213 ();
 sg13g2_decap_8 FILLER_80_2219 ();
 sg13g2_fill_2 FILLER_80_2263 ();
 sg13g2_fill_1 FILLER_80_2301 ();
 sg13g2_fill_1 FILLER_80_2309 ();
 sg13g2_fill_2 FILLER_80_2326 ();
 sg13g2_fill_1 FILLER_80_2332 ();
 sg13g2_fill_1 FILLER_80_2349 ();
 sg13g2_fill_1 FILLER_80_2357 ();
 sg13g2_fill_2 FILLER_80_2380 ();
 sg13g2_fill_2 FILLER_80_2404 ();
 sg13g2_fill_2 FILLER_80_2416 ();
 sg13g2_decap_4 FILLER_80_2435 ();
 sg13g2_fill_2 FILLER_80_2439 ();
 sg13g2_fill_2 FILLER_80_2451 ();
 sg13g2_decap_8 FILLER_80_2457 ();
 sg13g2_decap_8 FILLER_80_2464 ();
 sg13g2_decap_8 FILLER_80_2471 ();
 sg13g2_decap_4 FILLER_80_2478 ();
 sg13g2_fill_1 FILLER_80_2482 ();
 sg13g2_decap_4 FILLER_80_2493 ();
 sg13g2_fill_1 FILLER_80_2497 ();
 sg13g2_fill_1 FILLER_80_2502 ();
 sg13g2_decap_8 FILLER_80_2507 ();
 sg13g2_decap_8 FILLER_80_2514 ();
 sg13g2_decap_8 FILLER_80_2521 ();
 sg13g2_decap_8 FILLER_80_2528 ();
 sg13g2_decap_8 FILLER_80_2535 ();
 sg13g2_decap_8 FILLER_80_2542 ();
 sg13g2_decap_8 FILLER_80_2549 ();
 sg13g2_decap_8 FILLER_80_2560 ();
 sg13g2_decap_8 FILLER_80_2567 ();
 sg13g2_decap_8 FILLER_80_2574 ();
 sg13g2_decap_8 FILLER_80_2581 ();
 sg13g2_decap_8 FILLER_80_2588 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_4 FILLER_80_2665 ();
 sg13g2_fill_1 FILLER_80_2669 ();
endmodule
