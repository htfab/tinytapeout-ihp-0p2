module tt_um_tinytapeout_logo_screensaver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire clknet_0_clk;
 wire net217;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire \palette_inst.rrggbb[0] ;
 wire \palette_inst.rrggbb[1] ;
 wire \palette_inst.rrggbb[2] ;
 wire \palette_inst.rrggbb[3] ;
 wire \palette_inst.rrggbb[4] ;
 wire \palette_inst.rrggbb[5] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire \vga_sync_gen.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_dfrbp_1 \B[0]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net217),
    .D(_0015_),
    .Q_N(_2038_),
    .Q(net9));
 sg13g2_dfrbp_1 \B[1]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net218),
    .D(_0016_),
    .Q_N(_2037_),
    .Q(net5));
 sg13g2_dfrbp_1 \G[0]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net219),
    .D(_0017_),
    .Q_N(_2036_),
    .Q(net8));
 sg13g2_dfrbp_1 \G[1]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net220),
    .D(_0018_),
    .Q_N(_2035_),
    .Q(net4));
 sg13g2_dfrbp_1 \R[0]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net221),
    .D(_0019_),
    .Q_N(_2034_),
    .Q(net7));
 sg13g2_dfrbp_1 \R[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net222),
    .D(_0020_),
    .Q_N(_2033_),
    .Q(net3));
 sg13g2_buf_1 _2047_ (.A(\pix_y[1] ),
    .X(_0508_));
 sg13g2_inv_1 _2048_ (.Y(_0519_),
    .A(_0508_));
 sg13g2_buf_1 _2049_ (.A(\pix_y[5] ),
    .X(_0530_));
 sg13g2_buf_1 _2050_ (.A(_0530_),
    .X(_0541_));
 sg13g2_buf_1 _2051_ (.A(\pix_y[7] ),
    .X(_0552_));
 sg13g2_buf_1 _2052_ (.A(\pix_y[6] ),
    .X(_0563_));
 sg13g2_buf_1 _2053_ (.A(\pix_y[8] ),
    .X(_0574_));
 sg13g2_nand4_1 _2054_ (.B(_0552_),
    .C(net198),
    .A(net182),
    .Y(_0585_),
    .D(_0574_));
 sg13g2_buf_1 _2055_ (.A(\pix_y[2] ),
    .X(_0596_));
 sg13g2_buf_2 _2056_ (.A(\pix_y[9] ),
    .X(_0607_));
 sg13g2_or2_1 _2057_ (.X(_0618_),
    .B(_0607_),
    .A(net196));
 sg13g2_buf_1 _2058_ (.A(\pix_y[3] ),
    .X(_0629_));
 sg13g2_buf_1 _2059_ (.A(\pix_y[4] ),
    .X(_0640_));
 sg13g2_inv_1 _2060_ (.Y(_0651_),
    .A(net194));
 sg13g2_nand2_1 _2061_ (.Y(_0662_),
    .A(net195),
    .B(_0651_));
 sg13g2_nor4_1 _2062_ (.A(_0519_),
    .B(_0585_),
    .C(_0618_),
    .D(_0662_),
    .Y(_0005_));
 sg13g2_buf_1 _2063_ (.A(\pix_x[9] ),
    .X(_0683_));
 sg13g2_buf_1 _2064_ (.A(\pix_x[8] ),
    .X(_0694_));
 sg13g2_buf_2 _2065_ (.A(\pix_x[7] ),
    .X(_0705_));
 sg13g2_inv_1 _2066_ (.Y(_0716_),
    .A(_0705_));
 sg13g2_nor2_1 _2067_ (.A(net193),
    .B(_0716_),
    .Y(_0727_));
 sg13g2_buf_2 _2068_ (.A(\pix_x[6] ),
    .X(_0738_));
 sg13g2_buf_1 _2069_ (.A(\pix_x[5] ),
    .X(_0749_));
 sg13g2_buf_1 _2070_ (.A(_0749_),
    .X(_0760_));
 sg13g2_buf_1 _2071_ (.A(\pix_x[4] ),
    .X(_0771_));
 sg13g2_nand3_1 _2072_ (.B(net181),
    .C(net192),
    .A(_0738_),
    .Y(_0782_));
 sg13g2_inv_2 _2073_ (.Y(_0793_),
    .A(_0738_));
 sg13g2_inv_1 _2074_ (.Y(_0804_),
    .A(_0749_));
 sg13g2_inv_1 _2075_ (.Y(_0815_),
    .A(_0771_));
 sg13g2_nand3_1 _2076_ (.B(_0804_),
    .C(_0815_),
    .A(_0793_),
    .Y(_0826_));
 sg13g2_and4_1 _2077_ (.A(_0683_),
    .B(_0727_),
    .C(_0782_),
    .D(_0826_),
    .X(_0004_));
 sg13g2_buf_2 _2078_ (.A(rst_n),
    .X(_0847_));
 sg13g2_buf_1 _2079_ (.A(_0847_),
    .X(_0858_));
 sg13g2_buf_2 _2080_ (.A(dir_y),
    .X(_0869_));
 sg13g2_buf_2 _2081_ (.A(\logo_top[6] ),
    .X(_0880_));
 sg13g2_buf_1 _2082_ (.A(\logo_top[5] ),
    .X(_0891_));
 sg13g2_buf_1 _2083_ (.A(_0891_),
    .X(_0902_));
 sg13g2_buf_1 _2084_ (.A(_0012_),
    .X(_0913_));
 sg13g2_nor2_1 _2085_ (.A(net180),
    .B(_0913_),
    .Y(_0924_));
 sg13g2_nor2b_1 _2086_ (.A(_0880_),
    .B_N(net180),
    .Y(_0935_));
 sg13g2_a22oi_1 _2087_ (.Y(_0946_),
    .B1(_0935_),
    .B2(_0913_),
    .A2(_0924_),
    .A1(_0880_));
 sg13g2_buf_1 _2088_ (.A(\logo_top[9] ),
    .X(_0957_));
 sg13g2_buf_1 _2089_ (.A(\logo_top[8] ),
    .X(_0968_));
 sg13g2_inv_2 _2090_ (.Y(_0979_),
    .A(_0968_));
 sg13g2_buf_2 _2091_ (.A(\logo_top[7] ),
    .X(_0990_));
 sg13g2_buf_1 _2092_ (.A(\logo_top[4] ),
    .X(_1001_));
 sg13g2_inv_1 _2093_ (.Y(_1012_),
    .A(_1001_));
 sg13g2_nor4_1 _2094_ (.A(_0957_),
    .B(_0979_),
    .C(_0990_),
    .D(_1012_),
    .Y(_1023_));
 sg13g2_buf_1 _2095_ (.A(\logo_top[3] ),
    .X(_1034_));
 sg13g2_buf_2 _2096_ (.A(\logo_top[2] ),
    .X(_1045_));
 sg13g2_buf_1 _2097_ (.A(\logo_top[1] ),
    .X(_1055_));
 sg13g2_buf_1 _2098_ (.A(\logo_top[0] ),
    .X(_1065_));
 sg13g2_nand4_1 _2099_ (.B(_1045_),
    .C(_1055_),
    .A(net190),
    .Y(_1076_),
    .D(net188));
 sg13g2_inv_1 _2100_ (.Y(_1086_),
    .A(_1076_));
 sg13g2_nand3b_1 _2101_ (.B(_1023_),
    .C(_1086_),
    .Y(_1096_),
    .A_N(_0946_));
 sg13g2_inv_1 _2102_ (.Y(_1107_),
    .A(net188));
 sg13g2_nor4_1 _2103_ (.A(_0957_),
    .B(_0968_),
    .C(_0990_),
    .D(_1107_),
    .Y(_1115_));
 sg13g2_nor3_1 _2104_ (.A(_0880_),
    .B(net180),
    .C(_1001_),
    .Y(_1124_));
 sg13g2_nor3_1 _2105_ (.A(_1034_),
    .B(_1045_),
    .C(net189),
    .Y(_1133_));
 sg13g2_and3_1 _2106_ (.X(_1141_),
    .A(_1115_),
    .B(_1124_),
    .C(_1133_));
 sg13g2_nor2_1 _2107_ (.A(_0869_),
    .B(_1141_),
    .Y(_1151_));
 sg13g2_a21oi_1 _2108_ (.A1(_0869_),
    .A2(_1096_),
    .Y(_1161_),
    .B1(_1151_));
 sg13g2_buf_1 _2109_ (.A(dir_x),
    .X(_1170_));
 sg13g2_buf_1 _2110_ (.A(\logo_left[3] ),
    .X(_1179_));
 sg13g2_buf_1 _2111_ (.A(_1179_),
    .X(_1187_));
 sg13g2_buf_2 _2112_ (.A(\logo_left[2] ),
    .X(_1197_));
 sg13g2_buf_1 _2113_ (.A(\logo_left[1] ),
    .X(_1206_));
 sg13g2_buf_8 _2114_ (.A(\logo_left[0] ),
    .X(_1215_));
 sg13g2_and2_1 _2115_ (.A(net187),
    .B(net186),
    .X(_1225_));
 sg13g2_buf_1 _2116_ (.A(_1225_),
    .X(_1233_));
 sg13g2_nand3_1 _2117_ (.B(_1197_),
    .C(_1233_),
    .A(net179),
    .Y(_1234_));
 sg13g2_buf_1 _2118_ (.A(_1234_),
    .X(_1235_));
 sg13g2_buf_1 _2119_ (.A(\logo_left[9] ),
    .X(_1236_));
 sg13g2_buf_2 _2120_ (.A(\logo_left[4] ),
    .X(_1237_));
 sg13g2_buf_1 _2121_ (.A(_1237_),
    .X(_1238_));
 sg13g2_inv_1 _2122_ (.Y(_1239_),
    .A(net178));
 sg13g2_nor3_1 _2123_ (.A(_1236_),
    .B(_1239_),
    .C(_0011_),
    .Y(_1240_));
 sg13g2_buf_2 _2124_ (.A(\logo_left[6] ),
    .X(_1241_));
 sg13g2_buf_1 _2125_ (.A(\logo_left[5] ),
    .X(_1242_));
 sg13g2_buf_1 _2126_ (.A(net185),
    .X(_1243_));
 sg13g2_buf_1 _2127_ (.A(\logo_left[8] ),
    .X(_1244_));
 sg13g2_buf_1 _2128_ (.A(\logo_left[7] ),
    .X(_1245_));
 sg13g2_and2_1 _2129_ (.A(_1244_),
    .B(_1245_),
    .X(_1246_));
 sg13g2_and3_1 _2130_ (.X(_1247_),
    .A(_1241_),
    .B(net177),
    .C(_1246_));
 sg13g2_nand2_1 _2131_ (.Y(_1248_),
    .A(_1240_),
    .B(_1247_));
 sg13g2_nor2_1 _2132_ (.A(_1235_),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_inv_2 _2133_ (.Y(_1250_),
    .A(net179));
 sg13g2_nor3_1 _2134_ (.A(_1241_),
    .B(net185),
    .C(_1170_),
    .Y(_1251_));
 sg13g2_nand3_1 _2135_ (.B(_1250_),
    .C(_1251_),
    .A(_1239_),
    .Y(_1252_));
 sg13g2_nor2_1 _2136_ (.A(_1244_),
    .B(_1245_),
    .Y(_1253_));
 sg13g2_nand3b_1 _2137_ (.B(net186),
    .C(_1253_),
    .Y(_1254_),
    .A_N(net187));
 sg13g2_nor4_1 _2138_ (.A(_1236_),
    .B(_1197_),
    .C(_1252_),
    .D(_1254_),
    .Y(_1255_));
 sg13g2_a21o_1 _2139_ (.A2(_1249_),
    .A1(_1170_),
    .B1(_1255_),
    .X(_1256_));
 sg13g2_xnor2_1 _2140_ (.Y(_1257_),
    .A(_0541_),
    .B(\prev_y[5] ));
 sg13g2_xnor2_1 _2141_ (.Y(_1258_),
    .A(net194),
    .B(\prev_y[4] ));
 sg13g2_xnor2_1 _2142_ (.Y(_1259_),
    .A(\pix_y[8] ),
    .B(\prev_y[8] ));
 sg13g2_xnor2_1 _2143_ (.Y(_1260_),
    .A(\pix_y[7] ),
    .B(\prev_y[7] ));
 sg13g2_nand4_1 _2144_ (.B(_1258_),
    .C(_1259_),
    .A(_1257_),
    .Y(_1261_),
    .D(_1260_));
 sg13g2_xor2_1 _2145_ (.B(\prev_y[9] ),
    .A(_0607_),
    .X(_1262_));
 sg13g2_xor2_1 _2146_ (.B(\prev_y[3] ),
    .A(net195),
    .X(_1263_));
 sg13g2_buf_1 _2147_ (.A(_0508_),
    .X(_1264_));
 sg13g2_xnor2_1 _2148_ (.Y(_1265_),
    .A(_1264_),
    .B(\prev_y[1] ));
 sg13g2_buf_1 _2149_ (.A(\pix_y[0] ),
    .X(_1266_));
 sg13g2_buf_1 _2150_ (.A(_1266_),
    .X(_1267_));
 sg13g2_xnor2_1 _2151_ (.Y(_1268_),
    .A(_1267_),
    .B(\prev_y[0] ));
 sg13g2_xnor2_1 _2152_ (.Y(_1269_),
    .A(net198),
    .B(\prev_y[6] ));
 sg13g2_xnor2_1 _2153_ (.Y(_1270_),
    .A(net196),
    .B(\prev_y[2] ));
 sg13g2_nand4_1 _2154_ (.B(_1268_),
    .C(_1269_),
    .A(_1265_),
    .Y(_1271_),
    .D(_1270_));
 sg13g2_nor4_1 _2155_ (.A(_1261_),
    .B(_1262_),
    .C(_1263_),
    .D(_1271_),
    .Y(_1272_));
 sg13g2_nor4_1 _2156_ (.A(_1264_),
    .B(_1267_),
    .C(net182),
    .D(net194),
    .Y(_1273_));
 sg13g2_nor3_1 _2157_ (.A(_0552_),
    .B(net198),
    .C(\pix_y[8] ),
    .Y(_1274_));
 sg13g2_nand2_1 _2158_ (.Y(_1275_),
    .A(_1273_),
    .B(_1274_));
 sg13g2_nor4_2 _2159_ (.A(_0629_),
    .B(_0618_),
    .C(_1272_),
    .Y(_1276_),
    .D(_1275_));
 sg13g2_o21ai_1 _2160_ (.B1(_1276_),
    .Y(_1277_),
    .A1(_1161_),
    .A2(_1256_));
 sg13g2_buf_2 _2161_ (.A(_1277_),
    .X(_1278_));
 sg13g2_nand2_1 _2162_ (.Y(_1279_),
    .A(\color_index[1] ),
    .B(\color_index[0] ));
 sg13g2_nor2_1 _2163_ (.A(_1278_),
    .B(_1279_),
    .Y(_1280_));
 sg13g2_xnor2_1 _2164_ (.Y(_1281_),
    .A(_0007_),
    .B(_1280_));
 sg13g2_or2_1 _2165_ (.X(_1282_),
    .B(\color_index[0] ),
    .A(\color_index[1] ));
 sg13g2_a21oi_1 _2166_ (.A1(_1279_),
    .A2(_1282_),
    .Y(_1283_),
    .B1(_1278_));
 sg13g2_a21o_1 _2167_ (.A2(_1278_),
    .A1(_0008_),
    .B1(_1283_),
    .X(_1284_));
 sg13g2_buf_1 _2168_ (.A(_1284_),
    .X(_1285_));
 sg13g2_inv_1 _2169_ (.Y(_1286_),
    .A(_1285_));
 sg13g2_nand2_1 _2170_ (.Y(_1287_),
    .A(_1281_),
    .B(_1286_));
 sg13g2_xor2_1 _2171_ (.B(_1278_),
    .A(_0013_),
    .X(_1288_));
 sg13g2_nand3_1 _2172_ (.B(_1287_),
    .C(_1288_),
    .A(net191),
    .Y(_0000_));
 sg13g2_nand2_1 _2173_ (.Y(_1289_),
    .A(_1281_),
    .B(_1288_));
 sg13g2_xnor2_1 _2174_ (.Y(_1290_),
    .A(_1286_),
    .B(_1289_));
 sg13g2_nand2_1 _2175_ (.Y(_0001_),
    .A(_0858_),
    .B(_1290_));
 sg13g2_inv_1 _2176_ (.Y(_1291_),
    .A(_0847_));
 sg13g2_buf_1 _2177_ (.A(_1291_),
    .X(_1292_));
 sg13g2_nor2_1 _2178_ (.A(_1281_),
    .B(_1285_),
    .Y(_1293_));
 sg13g2_xnor2_1 _2179_ (.Y(_1294_),
    .A(_1288_),
    .B(_1293_));
 sg13g2_nor2_1 _2180_ (.A(_1292_),
    .B(_1294_),
    .Y(_0002_));
 sg13g2_nand2_1 _2181_ (.Y(_1295_),
    .A(_1285_),
    .B(_1288_));
 sg13g2_nor2_1 _2182_ (.A(_1281_),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_nor2b_1 _2183_ (.A(_1288_),
    .B_N(_1281_),
    .Y(_1297_));
 sg13g2_o21ai_1 _2184_ (.B1(_0858_),
    .Y(_0003_),
    .A1(_1296_),
    .A2(_1297_));
 sg13g2_buf_1 _2185_ (.A(_0847_),
    .X(_1298_));
 sg13g2_mux2_1 _2186_ (.A0(\prev_y[0] ),
    .A1(net175),
    .S(net183),
    .X(_0048_));
 sg13g2_mux2_1 _2187_ (.A0(\prev_y[1] ),
    .A1(net176),
    .S(_1298_),
    .X(_0049_));
 sg13g2_mux2_1 _2188_ (.A0(\prev_y[2] ),
    .A1(_0596_),
    .S(net183),
    .X(_0050_));
 sg13g2_mux2_1 _2189_ (.A0(\prev_y[3] ),
    .A1(net195),
    .S(net183),
    .X(_0051_));
 sg13g2_mux2_1 _2190_ (.A0(\prev_y[4] ),
    .A1(_0640_),
    .S(net183),
    .X(_0052_));
 sg13g2_mux2_1 _2191_ (.A0(\prev_y[5] ),
    .A1(_0541_),
    .S(net183),
    .X(_0053_));
 sg13g2_mux2_1 _2192_ (.A0(\prev_y[6] ),
    .A1(_0563_),
    .S(net183),
    .X(_0054_));
 sg13g2_mux2_1 _2193_ (.A0(\prev_y[7] ),
    .A1(net199),
    .S(net183),
    .X(_0055_));
 sg13g2_mux2_1 _2194_ (.A0(\prev_y[8] ),
    .A1(_0574_),
    .S(net183),
    .X(_0056_));
 sg13g2_mux2_1 _2195_ (.A0(\prev_y[9] ),
    .A1(_0607_),
    .S(_0847_),
    .X(_0057_));
 sg13g2_buf_2 _2196_ (.A(\pix_x[3] ),
    .X(_1299_));
 sg13g2_inv_2 _2197_ (.Y(_1300_),
    .A(_1299_));
 sg13g2_buf_8 _2198_ (.A(\pix_x[2] ),
    .X(_1301_));
 sg13g2_buf_2 _2199_ (.A(\pix_x[1] ),
    .X(_1302_));
 sg13g2_buf_2 _2200_ (.A(\pix_x[0] ),
    .X(_1303_));
 sg13g2_nand3_1 _2201_ (.B(_1302_),
    .C(_1303_),
    .A(_1301_),
    .Y(_1304_));
 sg13g2_buf_1 _2202_ (.A(_1304_),
    .X(_1305_));
 sg13g2_nor3_2 _2203_ (.A(_0815_),
    .B(_1300_),
    .C(_1305_),
    .Y(_1306_));
 sg13g2_nand2_1 _2204_ (.Y(_1307_),
    .A(net193),
    .B(_0683_));
 sg13g2_nor4_1 _2205_ (.A(_0705_),
    .B(_0738_),
    .C(net181),
    .D(_1307_),
    .Y(_1308_));
 sg13g2_and2_1 _2206_ (.A(_1306_),
    .B(_1308_),
    .X(_1309_));
 sg13g2_buf_1 _2207_ (.A(_1309_),
    .X(_1310_));
 sg13g2_nor2_1 _2208_ (.A(net184),
    .B(_1310_),
    .Y(_1311_));
 sg13g2_buf_2 _2209_ (.A(_1311_),
    .X(_1312_));
 sg13g2_nand3_1 _2210_ (.B(_0596_),
    .C(_0607_),
    .A(_0629_),
    .Y(_1313_));
 sg13g2_o21ai_1 _2211_ (.B1(_0847_),
    .Y(_1314_),
    .A1(_1275_),
    .A2(_1313_));
 sg13g2_buf_1 _2212_ (.A(_1314_),
    .X(_1315_));
 sg13g2_inv_1 _2213_ (.Y(_1316_),
    .A(_1315_));
 sg13g2_and2_1 _2214_ (.A(_1310_),
    .B(_1316_),
    .X(_1317_));
 sg13g2_buf_1 _2215_ (.A(_1317_),
    .X(_1318_));
 sg13g2_a22oi_1 _2216_ (.Y(_1319_),
    .B1(net133),
    .B2(_0010_),
    .A2(_1312_),
    .A1(net175));
 sg13g2_inv_1 _2217_ (.Y(_0068_),
    .A(_1319_));
 sg13g2_nand2_1 _2218_ (.Y(_1320_),
    .A(net175),
    .B(_1310_));
 sg13g2_xnor2_1 _2219_ (.Y(_1321_),
    .A(_0519_),
    .B(_1320_));
 sg13g2_nor2_1 _2220_ (.A(_1292_),
    .B(_1321_),
    .Y(_0069_));
 sg13g2_nand2_1 _2221_ (.Y(_1322_),
    .A(net176),
    .B(net175));
 sg13g2_xnor2_1 _2222_ (.Y(_1323_),
    .A(net196),
    .B(_1322_));
 sg13g2_a22oi_1 _2223_ (.Y(_1324_),
    .B1(net133),
    .B2(_1323_),
    .A2(_1312_),
    .A1(net196));
 sg13g2_inv_1 _2224_ (.Y(_0070_),
    .A(_1324_));
 sg13g2_and3_1 _2225_ (.X(_1325_),
    .A(net176),
    .B(net175),
    .C(net196));
 sg13g2_buf_1 _2226_ (.A(_1325_),
    .X(_1326_));
 sg13g2_nand2_1 _2227_ (.Y(_1327_),
    .A(net133),
    .B(_1326_));
 sg13g2_nor2_1 _2228_ (.A(_1315_),
    .B(_1326_),
    .Y(_1328_));
 sg13g2_o21ai_1 _2229_ (.B1(net195),
    .Y(_1329_),
    .A1(_1312_),
    .A2(_1328_));
 sg13g2_o21ai_1 _2230_ (.B1(_1329_),
    .Y(_0071_),
    .A1(net195),
    .A2(_1327_));
 sg13g2_and2_1 _2231_ (.A(net195),
    .B(_1326_),
    .X(_1330_));
 sg13g2_nand2_1 _2232_ (.Y(_1331_),
    .A(net133),
    .B(_1330_));
 sg13g2_nor2_1 _2233_ (.A(_1315_),
    .B(_1330_),
    .Y(_1332_));
 sg13g2_o21ai_1 _2234_ (.B1(net194),
    .Y(_1333_),
    .A1(_1312_),
    .A2(_1332_));
 sg13g2_o21ai_1 _2235_ (.B1(_1333_),
    .Y(_0072_),
    .A1(net194),
    .A2(_1331_));
 sg13g2_and2_1 _2236_ (.A(net194),
    .B(_1330_),
    .X(_1334_));
 sg13g2_nand2_1 _2237_ (.Y(_1335_),
    .A(net133),
    .B(_1334_));
 sg13g2_nor2_1 _2238_ (.A(_1315_),
    .B(_1334_),
    .Y(_1336_));
 sg13g2_o21ai_1 _2239_ (.B1(net182),
    .Y(_1337_),
    .A1(_1312_),
    .A2(_1336_));
 sg13g2_o21ai_1 _2240_ (.B1(_1337_),
    .Y(_0073_),
    .A1(net182),
    .A2(_1335_));
 sg13g2_and2_1 _2241_ (.A(net182),
    .B(_1334_),
    .X(_1338_));
 sg13g2_nand2_1 _2242_ (.Y(_1339_),
    .A(_1318_),
    .B(_1338_));
 sg13g2_nor2_1 _2243_ (.A(_1315_),
    .B(_1338_),
    .Y(_1340_));
 sg13g2_o21ai_1 _2244_ (.B1(net198),
    .Y(_1341_),
    .A1(_1312_),
    .A2(_1340_));
 sg13g2_o21ai_1 _2245_ (.B1(_1341_),
    .Y(_0074_),
    .A1(net198),
    .A2(_1339_));
 sg13g2_and2_1 _2246_ (.A(net198),
    .B(_1338_),
    .X(_1342_));
 sg13g2_buf_1 _2247_ (.A(_1342_),
    .X(_1343_));
 sg13g2_nand2_1 _2248_ (.Y(_1344_),
    .A(net133),
    .B(_1343_));
 sg13g2_nand2b_1 _2249_ (.Y(_1345_),
    .B(_0847_),
    .A_N(_1310_));
 sg13g2_buf_1 _2250_ (.A(_1345_),
    .X(_1346_));
 sg13g2_o21ai_1 _2251_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1315_),
    .A2(_1343_));
 sg13g2_nand2_1 _2252_ (.Y(_1348_),
    .A(net199),
    .B(_1347_));
 sg13g2_o21ai_1 _2253_ (.B1(_1348_),
    .Y(_0075_),
    .A1(net199),
    .A2(_1344_));
 sg13g2_and2_1 _2254_ (.A(net199),
    .B(_1343_),
    .X(_1349_));
 sg13g2_buf_1 _2255_ (.A(_1349_),
    .X(_1350_));
 sg13g2_nand2_1 _2256_ (.Y(_1351_),
    .A(net133),
    .B(_1350_));
 sg13g2_nand2_1 _2257_ (.Y(_1352_),
    .A(_1310_),
    .B(_1316_));
 sg13g2_o21ai_1 _2258_ (.B1(_1346_),
    .Y(_1353_),
    .A1(_1352_),
    .A2(_1350_));
 sg13g2_nand2_1 _2259_ (.Y(_1354_),
    .A(net197),
    .B(_1353_));
 sg13g2_o21ai_1 _2260_ (.B1(_1354_),
    .Y(_0076_),
    .A1(net197),
    .A2(_1351_));
 sg13g2_nand3_1 _2261_ (.B(net133),
    .C(_1350_),
    .A(net197),
    .Y(_1355_));
 sg13g2_a21oi_1 _2262_ (.A1(net197),
    .A2(_1350_),
    .Y(_1356_),
    .B1(_1352_));
 sg13g2_o21ai_1 _2263_ (.B1(_0607_),
    .Y(_1357_),
    .A1(_1312_),
    .A2(_1356_));
 sg13g2_o21ai_1 _2264_ (.B1(_1357_),
    .Y(_0077_),
    .A1(_0607_),
    .A2(_1355_));
 sg13g2_o21ai_1 _2265_ (.B1(_0847_),
    .Y(_1358_),
    .A1(_1281_),
    .A2(_1288_));
 sg13g2_inv_1 _2266_ (.Y(_0046_),
    .A(_1358_));
 sg13g2_o21ai_1 _2267_ (.B1(_1358_),
    .Y(_0047_),
    .A1(net184),
    .A2(_1285_));
 sg13g2_and2_1 _2268_ (.A(_0014_),
    .B(_1312_),
    .X(_0058_));
 sg13g2_xnor2_1 _2269_ (.Y(_1359_),
    .A(_1302_),
    .B(_1303_));
 sg13g2_nor2_1 _2270_ (.A(net174),
    .B(_1359_),
    .Y(_0059_));
 sg13g2_inv_1 _2271_ (.Y(_1360_),
    .A(_1301_));
 sg13g2_nand2_1 _2272_ (.Y(_1361_),
    .A(_1302_),
    .B(_1303_));
 sg13g2_xnor2_1 _2273_ (.Y(_1362_),
    .A(_1360_),
    .B(_1361_));
 sg13g2_nor2_1 _2274_ (.A(net174),
    .B(_1362_),
    .Y(_0060_));
 sg13g2_xnor2_1 _2275_ (.Y(_1363_),
    .A(_1300_),
    .B(_1305_));
 sg13g2_nor2_1 _2276_ (.A(net174),
    .B(_1363_),
    .Y(_0061_));
 sg13g2_nor2_1 _2277_ (.A(_1300_),
    .B(_1305_),
    .Y(_1364_));
 sg13g2_xnor2_1 _2278_ (.Y(_1365_),
    .A(net192),
    .B(_1364_));
 sg13g2_nor2_1 _2279_ (.A(net174),
    .B(_1365_),
    .Y(_0062_));
 sg13g2_xnor2_1 _2280_ (.Y(_1366_),
    .A(net181),
    .B(_1306_));
 sg13g2_nor2_1 _2281_ (.A(_1346_),
    .B(_1366_),
    .Y(_0063_));
 sg13g2_nand2_1 _2282_ (.Y(_1367_),
    .A(_0760_),
    .B(_1306_));
 sg13g2_xnor2_1 _2283_ (.Y(_1368_),
    .A(_0793_),
    .B(_1367_));
 sg13g2_nor2_1 _2284_ (.A(net174),
    .B(_1368_),
    .Y(_0064_));
 sg13g2_nand3_1 _2285_ (.B(net181),
    .C(_1306_),
    .A(_0738_),
    .Y(_1369_));
 sg13g2_xnor2_1 _2286_ (.Y(_1370_),
    .A(_0716_),
    .B(_1369_));
 sg13g2_nor2_1 _2287_ (.A(net174),
    .B(_1370_),
    .Y(_0065_));
 sg13g2_nor2_1 _2288_ (.A(_0716_),
    .B(_1369_),
    .Y(_1371_));
 sg13g2_xnor2_1 _2289_ (.Y(_1372_),
    .A(net193),
    .B(_1371_));
 sg13g2_nor2_1 _2290_ (.A(_1346_),
    .B(_1372_),
    .Y(_0066_));
 sg13g2_nand2_1 _2291_ (.Y(_1373_),
    .A(_0694_),
    .B(_1371_));
 sg13g2_xor2_1 _2292_ (.B(_1373_),
    .A(_0683_),
    .X(_1374_));
 sg13g2_nor2_1 _2293_ (.A(_1346_),
    .B(_1374_),
    .Y(_0067_));
 sg13g2_nor2b_1 _2294_ (.A(_1045_),
    .B_N(net196),
    .Y(_1375_));
 sg13g2_nand2b_1 _2295_ (.Y(_1376_),
    .B(net190),
    .A_N(net195));
 sg13g2_nor2b_1 _2296_ (.A(net190),
    .B_N(net195),
    .Y(_1377_));
 sg13g2_a21oi_2 _2297_ (.B1(_1377_),
    .Y(_1378_),
    .A2(_1376_),
    .A1(_1375_));
 sg13g2_nor2b_1 _2298_ (.A(_1266_),
    .B_N(net188),
    .Y(_1379_));
 sg13g2_buf_2 _2299_ (.A(_1379_),
    .X(_1380_));
 sg13g2_nand2_1 _2300_ (.Y(_1381_),
    .A(net189),
    .B(_1380_));
 sg13g2_o21ai_1 _2301_ (.B1(_0519_),
    .Y(_1382_),
    .A1(net189),
    .A2(_1380_));
 sg13g2_nand2b_1 _2302_ (.Y(_1383_),
    .B(_1045_),
    .A_N(net196));
 sg13g2_nand4_1 _2303_ (.B(_1381_),
    .C(_1382_),
    .A(_1376_),
    .Y(_1384_),
    .D(_1383_));
 sg13g2_nand2_1 _2304_ (.Y(_1385_),
    .A(_1378_),
    .B(_1384_));
 sg13g2_nor2_1 _2305_ (.A(net194),
    .B(_1012_),
    .Y(_1386_));
 sg13g2_nand2_1 _2306_ (.Y(_1387_),
    .A(net194),
    .B(_1012_));
 sg13g2_nand2b_1 _2307_ (.Y(_1388_),
    .B(_1387_),
    .A_N(_1386_));
 sg13g2_xor2_1 _2308_ (.B(_1388_),
    .A(_1385_),
    .X(_1389_));
 sg13g2_buf_2 _2309_ (.A(_1389_),
    .X(_1390_));
 sg13g2_buf_1 _2310_ (.A(_1390_),
    .X(_1391_));
 sg13g2_buf_1 _2311_ (.A(net132),
    .X(_1392_));
 sg13g2_inv_1 _2312_ (.Y(_1393_),
    .A(\logo_top[1] ));
 sg13g2_nand2b_2 _2313_ (.Y(_1394_),
    .B(net188),
    .A_N(_1266_));
 sg13g2_nor2_1 _2314_ (.A(_1393_),
    .B(_1394_),
    .Y(_1395_));
 sg13g2_a21oi_1 _2315_ (.A1(_1393_),
    .A2(_1394_),
    .Y(_1396_),
    .B1(_0508_));
 sg13g2_xnor2_1 _2316_ (.Y(_1397_),
    .A(\pix_y[3] ),
    .B(net190));
 sg13g2_nor2_1 _2317_ (.A(_1375_),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_o21ai_1 _2318_ (.B1(_1398_),
    .Y(_1399_),
    .A1(_1395_),
    .A2(_1396_));
 sg13g2_nand4_1 _2319_ (.B(_1382_),
    .C(_1383_),
    .A(_1381_),
    .Y(_1400_),
    .D(_1397_));
 sg13g2_nor2_1 _2320_ (.A(_1383_),
    .B(_1397_),
    .Y(_1401_));
 sg13g2_a21oi_1 _2321_ (.A1(_1375_),
    .A2(_1397_),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_and3_1 _2322_ (.X(_1403_),
    .A(_1399_),
    .B(_1400_),
    .C(_1402_));
 sg13g2_buf_2 _2323_ (.A(_1403_),
    .X(_1404_));
 sg13g2_xnor2_1 _2324_ (.Y(_1405_),
    .A(_0508_),
    .B(net189));
 sg13g2_xnor2_1 _2325_ (.Y(_1406_),
    .A(_1394_),
    .B(_1405_));
 sg13g2_buf_1 _2326_ (.A(_1406_),
    .X(_1407_));
 sg13g2_xnor2_1 _2327_ (.Y(_1408_),
    .A(net196),
    .B(_1045_));
 sg13g2_nand3_1 _2328_ (.B(_1382_),
    .C(_1408_),
    .A(_1381_),
    .Y(_1409_));
 sg13g2_buf_2 _2329_ (.A(_1409_),
    .X(_1410_));
 sg13g2_nand2b_1 _2330_ (.Y(_1411_),
    .B(_1383_),
    .A_N(_1375_));
 sg13g2_o21ai_1 _2331_ (.B1(_1411_),
    .Y(_1412_),
    .A1(_1395_),
    .A2(_1396_));
 sg13g2_buf_1 _2332_ (.A(_1412_),
    .X(_1413_));
 sg13g2_and2_1 _2333_ (.A(_1410_),
    .B(_1413_),
    .X(_1414_));
 sg13g2_buf_1 _2334_ (.A(_1414_),
    .X(_1415_));
 sg13g2_nor2_1 _2335_ (.A(_1407_),
    .B(_1415_),
    .Y(_1416_));
 sg13g2_nand2_1 _2336_ (.Y(_1417_),
    .A(_1404_),
    .B(_1416_));
 sg13g2_nor2b_1 _2337_ (.A(net188),
    .B_N(_1266_),
    .Y(_1418_));
 sg13g2_nor2_1 _2338_ (.A(_1380_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_buf_1 _2339_ (.A(_1419_),
    .X(_1420_));
 sg13g2_buf_1 _2340_ (.A(_1420_),
    .X(_1421_));
 sg13g2_nor2b_1 _2341_ (.A(_1197_),
    .B_N(_1301_),
    .Y(_1422_));
 sg13g2_buf_1 _2342_ (.A(_1422_),
    .X(_1423_));
 sg13g2_nor2b_1 _2343_ (.A(_1303_),
    .B_N(net186),
    .Y(_1424_));
 sg13g2_nand2b_1 _2344_ (.Y(_1425_),
    .B(_1302_),
    .A_N(net187));
 sg13g2_nor2b_1 _2345_ (.A(_1302_),
    .B_N(net187),
    .Y(_1426_));
 sg13g2_a221oi_1 _2346_ (.B2(_1425_),
    .C1(_1426_),
    .B1(_1424_),
    .A1(_1197_),
    .Y(_1427_),
    .A2(_1360_));
 sg13g2_buf_2 _2347_ (.A(_1427_),
    .X(_1428_));
 sg13g2_o21ai_1 _2348_ (.B1(_1299_),
    .Y(_1429_),
    .A1(net170),
    .A2(_1428_));
 sg13g2_buf_1 _2349_ (.A(_1429_),
    .X(_1430_));
 sg13g2_or2_1 _2350_ (.X(_1431_),
    .B(net170),
    .A(_1299_));
 sg13g2_buf_1 _2351_ (.A(_1431_),
    .X(_1432_));
 sg13g2_o21ai_1 _2352_ (.B1(_1250_),
    .Y(_1433_),
    .A1(_1428_),
    .A2(_1432_));
 sg13g2_buf_2 _2353_ (.A(_1433_),
    .X(_1434_));
 sg13g2_xnor2_1 _2354_ (.Y(_1435_),
    .A(net185),
    .B(net181));
 sg13g2_buf_1 _2355_ (.A(_1435_),
    .X(_1436_));
 sg13g2_nand3_1 _2356_ (.B(_0815_),
    .C(_1436_),
    .A(_1239_),
    .Y(_1437_));
 sg13g2_nand3_1 _2357_ (.B(net192),
    .C(_1436_),
    .A(_1238_),
    .Y(_1438_));
 sg13g2_a22oi_1 _2358_ (.Y(_1439_),
    .B1(_1437_),
    .B2(_1438_),
    .A2(_1434_),
    .A1(net160));
 sg13g2_a21o_1 _2359_ (.A2(_1425_),
    .A1(_1424_),
    .B1(_1426_),
    .X(_1440_));
 sg13g2_a221oi_1 _2360_ (.B2(_1440_),
    .C1(_1197_),
    .B1(_1360_),
    .A1(net179),
    .Y(_1441_),
    .A2(_1300_));
 sg13g2_buf_2 _2361_ (.A(_1441_),
    .X(_1442_));
 sg13g2_inv_1 _2362_ (.Y(_1443_),
    .A(_1302_));
 sg13g2_o21ai_1 _2363_ (.B1(net187),
    .Y(_1444_),
    .A1(_1443_),
    .A2(_1424_));
 sg13g2_a221oi_1 _2364_ (.B2(_1424_),
    .C1(_1360_),
    .B1(_1443_),
    .A1(_1179_),
    .Y(_1445_),
    .A2(_1300_));
 sg13g2_nor2b_1 _2365_ (.A(_1179_),
    .B_N(_1299_),
    .Y(_1446_));
 sg13g2_a21o_1 _2366_ (.A2(_1445_),
    .A1(_1444_),
    .B1(_1446_),
    .X(_1447_));
 sg13g2_buf_2 _2367_ (.A(_1447_),
    .X(_1448_));
 sg13g2_nand2b_1 _2368_ (.Y(_1449_),
    .B(net178),
    .A_N(net192));
 sg13g2_nor4_1 _2369_ (.A(_1442_),
    .B(_1448_),
    .C(_1436_),
    .D(_1449_),
    .Y(_1450_));
 sg13g2_xor2_1 _2370_ (.B(net181),
    .A(net185),
    .X(_1451_));
 sg13g2_nand2b_1 _2371_ (.Y(_1452_),
    .B(\pix_x[4] ),
    .A_N(_1237_));
 sg13g2_buf_2 _2372_ (.A(_1452_),
    .X(_1453_));
 sg13g2_nor4_1 _2373_ (.A(_1442_),
    .B(_1448_),
    .C(_1451_),
    .D(_1453_),
    .Y(_1454_));
 sg13g2_nor3_1 _2374_ (.A(_1439_),
    .B(_1450_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_buf_2 _2375_ (.A(_1455_),
    .X(_1456_));
 sg13g2_nor2_1 _2376_ (.A(net161),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_buf_8 _2377_ (.A(_1428_),
    .X(_1458_));
 sg13g2_nor2b_1 _2378_ (.A(_1299_),
    .B_N(net179),
    .Y(_1459_));
 sg13g2_xor2_1 _2379_ (.B(net192),
    .A(_1237_),
    .X(_1460_));
 sg13g2_buf_2 _2380_ (.A(_1460_),
    .X(_1461_));
 sg13g2_nor2_1 _2381_ (.A(_1459_),
    .B(_1461_),
    .Y(_1462_));
 sg13g2_o21ai_1 _2382_ (.B1(_1462_),
    .Y(_1463_),
    .A1(_1423_),
    .A2(_1458_));
 sg13g2_xnor2_1 _2383_ (.Y(_1464_),
    .A(_1241_),
    .B(_0738_));
 sg13g2_nand3b_1 _2384_ (.B(_0749_),
    .C(net192),
    .Y(_1465_),
    .A_N(_1237_));
 sg13g2_and2_1 _2385_ (.A(_1464_),
    .B(_1465_),
    .X(_1466_));
 sg13g2_a21o_1 _2386_ (.A2(_1453_),
    .A1(_0804_),
    .B1(net185),
    .X(_1467_));
 sg13g2_a21oi_1 _2387_ (.A1(net185),
    .A2(_1453_),
    .Y(_1468_),
    .B1(_1464_));
 sg13g2_o21ai_1 _2388_ (.B1(_0804_),
    .Y(_1469_),
    .A1(net185),
    .A2(_1453_));
 sg13g2_nand2b_1 _2389_ (.Y(_1470_),
    .B(_1299_),
    .A_N(net179));
 sg13g2_nor2_1 _2390_ (.A(_1470_),
    .B(_1461_),
    .Y(_1471_));
 sg13g2_a221oi_1 _2391_ (.B2(_1469_),
    .C1(_1471_),
    .B1(_1468_),
    .A1(_1466_),
    .Y(_1472_),
    .A2(_1467_));
 sg13g2_nand2_1 _2392_ (.Y(_1473_),
    .A(_1463_),
    .B(_1472_));
 sg13g2_nor2b_1 _2393_ (.A(_0749_),
    .B_N(net185),
    .Y(_1474_));
 sg13g2_xnor2_1 _2394_ (.Y(_1475_),
    .A(_1474_),
    .B(_1464_));
 sg13g2_and2_1 _2395_ (.A(_1453_),
    .B(_1449_),
    .X(_1476_));
 sg13g2_buf_1 _2396_ (.A(_1476_),
    .X(_1477_));
 sg13g2_nand2b_1 _2397_ (.Y(_1478_),
    .B(net164),
    .A_N(_1475_));
 sg13g2_a21o_1 _2398_ (.A2(_1434_),
    .A1(net160),
    .B1(_1478_),
    .X(_1479_));
 sg13g2_buf_2 _2399_ (.A(_1479_),
    .X(_1480_));
 sg13g2_nand2_1 _2400_ (.Y(_1481_),
    .A(_1473_),
    .B(_1480_));
 sg13g2_buf_1 _2401_ (.A(_1481_),
    .X(_1482_));
 sg13g2_buf_1 _2402_ (.A(net85),
    .X(_1483_));
 sg13g2_buf_1 _2403_ (.A(net60),
    .X(_1484_));
 sg13g2_and2_1 _2404_ (.A(net179),
    .B(_1453_),
    .X(_1485_));
 sg13g2_o21ai_1 _2405_ (.B1(net192),
    .Y(_1486_),
    .A1(_1428_),
    .A2(_1432_));
 sg13g2_nor4_1 _2406_ (.A(net192),
    .B(_1299_),
    .C(net170),
    .D(net165),
    .Y(_1487_));
 sg13g2_a221oi_1 _2407_ (.B2(net178),
    .C1(_1487_),
    .B1(_1486_),
    .A1(_1429_),
    .Y(_1488_),
    .A2(_1485_));
 sg13g2_buf_2 _2408_ (.A(_1488_),
    .X(_1489_));
 sg13g2_xnor2_1 _2409_ (.Y(_1490_),
    .A(_1451_),
    .B(_1489_));
 sg13g2_buf_8 _2410_ (.A(_1490_),
    .X(_1491_));
 sg13g2_buf_8 _2411_ (.A(_1491_),
    .X(_1492_));
 sg13g2_buf_1 _2412_ (.A(net84),
    .X(_1493_));
 sg13g2_nor2_1 _2413_ (.A(net165),
    .B(_1432_),
    .Y(_1494_));
 sg13g2_or2_1 _2414_ (.X(_1495_),
    .B(net165),
    .A(_1423_));
 sg13g2_a22oi_1 _2415_ (.Y(_1496_),
    .B1(_1446_),
    .B2(_1495_),
    .A2(_1494_),
    .A1(net179));
 sg13g2_xnor2_1 _2416_ (.Y(_1497_),
    .A(_1461_),
    .B(_1496_));
 sg13g2_buf_1 _2417_ (.A(_1497_),
    .X(_1498_));
 sg13g2_and2_1 _2418_ (.A(_1493_),
    .B(_1498_),
    .X(_1499_));
 sg13g2_nor4_1 _2419_ (.A(_1417_),
    .B(_1457_),
    .C(net36),
    .D(_1499_),
    .Y(_1500_));
 sg13g2_and2_1 _2420_ (.A(_1463_),
    .B(_1472_),
    .X(_1501_));
 sg13g2_buf_2 _2421_ (.A(_1501_),
    .X(_1502_));
 sg13g2_a21oi_1 _2422_ (.A1(net160),
    .A2(_1434_),
    .Y(_1503_),
    .B1(_1478_));
 sg13g2_buf_2 _2423_ (.A(_1503_),
    .X(_1504_));
 sg13g2_nor2_1 _2424_ (.A(_1502_),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_buf_2 _2425_ (.A(_1505_),
    .X(_1506_));
 sg13g2_buf_1 _2426_ (.A(_1506_),
    .X(_1507_));
 sg13g2_buf_1 _2427_ (.A(net58),
    .X(_1508_));
 sg13g2_buf_8 _2428_ (.A(_1491_),
    .X(_1509_));
 sg13g2_o21ai_1 _2429_ (.B1(net164),
    .Y(_1510_),
    .A1(_1442_),
    .A2(_1448_));
 sg13g2_buf_1 _2430_ (.A(_1510_),
    .X(_1511_));
 sg13g2_nand3_1 _2431_ (.B(_1434_),
    .C(_1461_),
    .A(net160),
    .Y(_1512_));
 sg13g2_buf_2 _2432_ (.A(_1512_),
    .X(_1513_));
 sg13g2_nand2_1 _2433_ (.Y(_1514_),
    .A(net155),
    .B(_1513_));
 sg13g2_buf_2 _2434_ (.A(_1514_),
    .X(_1515_));
 sg13g2_nor2_1 _2435_ (.A(net83),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_buf_1 _2436_ (.A(_1516_),
    .X(_1517_));
 sg13g2_xnor2_1 _2437_ (.Y(_1518_),
    .A(_1436_),
    .B(_1489_));
 sg13g2_buf_8 _2438_ (.A(_1518_),
    .X(_1519_));
 sg13g2_buf_1 _2439_ (.A(net113),
    .X(_1520_));
 sg13g2_nor2_1 _2440_ (.A(_1421_),
    .B(net82),
    .Y(_1521_));
 sg13g2_nor4_1 _2441_ (.A(_1417_),
    .B(_1508_),
    .C(net34),
    .D(_1521_),
    .Y(_1522_));
 sg13g2_nor3_1 _2442_ (.A(net114),
    .B(_1500_),
    .C(_1522_),
    .Y(_1523_));
 sg13g2_nor2_1 _2443_ (.A(_1519_),
    .B(net85),
    .Y(_1524_));
 sg13g2_buf_1 _2444_ (.A(_1524_),
    .X(_1525_));
 sg13g2_xnor2_1 _2445_ (.Y(_1526_),
    .A(_1187_),
    .B(_1299_));
 sg13g2_o21ai_1 _2446_ (.B1(_1526_),
    .Y(_1527_),
    .A1(net170),
    .A2(net165));
 sg13g2_buf_1 _2447_ (.A(_1527_),
    .X(_1528_));
 sg13g2_or3_1 _2448_ (.A(net170),
    .B(net165),
    .C(_1526_),
    .X(_1529_));
 sg13g2_buf_2 _2449_ (.A(_1529_),
    .X(_1530_));
 sg13g2_nand2_1 _2450_ (.Y(_1531_),
    .A(_1528_),
    .B(_1530_));
 sg13g2_buf_1 _2451_ (.A(_1531_),
    .X(_1532_));
 sg13g2_nand3_1 _2452_ (.B(_1513_),
    .C(net131),
    .A(_1511_),
    .Y(_1533_));
 sg13g2_buf_2 _2453_ (.A(_1533_),
    .X(_1534_));
 sg13g2_mux2_1 _2454_ (.A0(_1446_),
    .A1(_1459_),
    .S(_1461_),
    .X(_1535_));
 sg13g2_o21ai_1 _2455_ (.B1(_1535_),
    .Y(_1536_),
    .A1(net170),
    .A2(_1458_));
 sg13g2_inv_1 _2456_ (.Y(_1537_),
    .A(_1526_));
 sg13g2_or4_1 _2457_ (.A(net170),
    .B(net165),
    .C(net164),
    .D(_1537_),
    .X(_1538_));
 sg13g2_and2_1 _2458_ (.A(_1536_),
    .B(_1538_),
    .X(_1539_));
 sg13g2_buf_1 _2459_ (.A(_1539_),
    .X(_1540_));
 sg13g2_o21ai_1 _2460_ (.B1(net145),
    .Y(_1541_),
    .A1(net161),
    .A2(_1534_));
 sg13g2_nand2_1 _2461_ (.Y(_1542_),
    .A(net33),
    .B(_1541_));
 sg13g2_buf_1 _2462_ (.A(_1518_),
    .X(_1543_));
 sg13g2_a221oi_1 _2463_ (.B2(_1469_),
    .C1(_1477_),
    .B1(_1468_),
    .A1(_1466_),
    .Y(_1544_),
    .A2(_1467_));
 sg13g2_o21ai_1 _2464_ (.B1(_1544_),
    .Y(_1545_),
    .A1(_1442_),
    .A2(_1448_));
 sg13g2_a22oi_1 _2465_ (.Y(_1546_),
    .B1(_1468_),
    .B2(_1469_),
    .A2(_1467_),
    .A1(_1466_));
 sg13g2_buf_1 _2466_ (.A(_1546_),
    .X(_1547_));
 sg13g2_nand4_1 _2467_ (.B(_1434_),
    .C(net164),
    .A(net160),
    .Y(_1548_),
    .D(_1547_));
 sg13g2_nand2_1 _2468_ (.Y(_1549_),
    .A(_1545_),
    .B(_1548_));
 sg13g2_buf_2 _2469_ (.A(_1549_),
    .X(_1550_));
 sg13g2_nand2_1 _2470_ (.Y(_1551_),
    .A(net112),
    .B(_1550_));
 sg13g2_buf_2 _2471_ (.A(_1551_),
    .X(_1552_));
 sg13g2_nand3_1 _2472_ (.B(_1400_),
    .C(_1402_),
    .A(_1399_),
    .Y(_1553_));
 sg13g2_buf_1 _2473_ (.A(_1553_),
    .X(_1554_));
 sg13g2_xnor2_1 _2474_ (.Y(_1555_),
    .A(_1380_),
    .B(_1405_));
 sg13g2_a21o_1 _2475_ (.A2(_1413_),
    .A1(_1410_),
    .B1(_1555_),
    .X(_1556_));
 sg13g2_buf_1 _2476_ (.A(_1556_),
    .X(_1557_));
 sg13g2_nor2_1 _2477_ (.A(net154),
    .B(net144),
    .Y(_1558_));
 sg13g2_nand3_1 _2478_ (.B(_1552_),
    .C(_1558_),
    .A(_1542_),
    .Y(_1559_));
 sg13g2_buf_8 _2479_ (.A(net83),
    .X(_1560_));
 sg13g2_buf_8 _2480_ (.A(net57),
    .X(_1561_));
 sg13g2_buf_1 _2481_ (.A(net32),
    .X(_1562_));
 sg13g2_and2_1 _2482_ (.A(_1477_),
    .B(_1475_),
    .X(_1563_));
 sg13g2_o21ai_1 _2483_ (.B1(_1563_),
    .Y(_1564_),
    .A1(_1442_),
    .A2(_1448_));
 sg13g2_buf_1 _2484_ (.A(_1564_),
    .X(_1565_));
 sg13g2_or4_1 _2485_ (.A(_1442_),
    .B(_1448_),
    .C(net164),
    .D(_1547_),
    .X(_1566_));
 sg13g2_buf_1 _2486_ (.A(_1566_),
    .X(_1567_));
 sg13g2_nand4_1 _2487_ (.B(_1545_),
    .C(_1548_),
    .A(_1565_),
    .Y(_1568_),
    .D(_1567_));
 sg13g2_nor2_1 _2488_ (.A(net15),
    .B(_1568_),
    .Y(_1569_));
 sg13g2_and2_1 _2489_ (.A(_1301_),
    .B(_1302_),
    .X(_1570_));
 sg13g2_nor2b_1 _2490_ (.A(net187),
    .B_N(_1301_),
    .Y(_1571_));
 sg13g2_nand2b_1 _2491_ (.Y(_1572_),
    .B(net186),
    .A_N(_1303_));
 sg13g2_o21ai_1 _2492_ (.B1(_1572_),
    .Y(_1573_),
    .A1(_1570_),
    .A2(_1571_));
 sg13g2_inv_2 _2493_ (.Y(_1574_),
    .A(_1197_));
 sg13g2_a21oi_1 _2494_ (.A1(_1302_),
    .A2(_1571_),
    .Y(_1575_),
    .B1(_1574_));
 sg13g2_a221oi_1 _2495_ (.B2(_1575_),
    .C1(_1537_),
    .B1(_1573_),
    .A1(_1360_),
    .Y(_1576_),
    .A2(_1440_));
 sg13g2_nor3_2 _2496_ (.A(net170),
    .B(net165),
    .C(_1526_),
    .Y(_1577_));
 sg13g2_nor2_1 _2497_ (.A(_1576_),
    .B(_1577_),
    .Y(_1578_));
 sg13g2_buf_1 _2498_ (.A(_1578_),
    .X(_1579_));
 sg13g2_nand3_1 _2499_ (.B(_1513_),
    .C(net143),
    .A(net155),
    .Y(_1580_));
 sg13g2_buf_2 _2500_ (.A(_1580_),
    .X(_1581_));
 sg13g2_buf_1 _2501_ (.A(_1581_),
    .X(_1582_));
 sg13g2_buf_8 _2502_ (.A(net83),
    .X(_1583_));
 sg13g2_or2_1 _2503_ (.X(_1584_),
    .B(_1432_),
    .A(net165));
 sg13g2_nand4_1 _2504_ (.B(_1430_),
    .C(_1584_),
    .A(_1250_),
    .Y(_1585_),
    .D(net164));
 sg13g2_buf_1 _2505_ (.A(_1585_),
    .X(_1586_));
 sg13g2_nor2_1 _2506_ (.A(_1250_),
    .B(net164),
    .Y(_1587_));
 sg13g2_nor3_1 _2507_ (.A(_1250_),
    .B(_1300_),
    .C(_1461_),
    .Y(_1588_));
 sg13g2_a22oi_1 _2508_ (.Y(_1589_),
    .B1(_1588_),
    .B2(_1495_),
    .A2(_1587_),
    .A1(_1494_));
 sg13g2_buf_2 _2509_ (.A(_1589_),
    .X(_1590_));
 sg13g2_nand2_1 _2510_ (.Y(_1591_),
    .A(_1586_),
    .B(_1590_));
 sg13g2_buf_1 _2511_ (.A(_1591_),
    .X(_1592_));
 sg13g2_nand2_2 _2512_ (.Y(_1593_),
    .A(net55),
    .B(net111));
 sg13g2_buf_1 _2513_ (.A(net60),
    .X(_1594_));
 sg13g2_a21oi_1 _2514_ (.A1(net56),
    .A2(_1593_),
    .Y(_1595_),
    .B1(_1594_));
 sg13g2_nand2_1 _2515_ (.Y(_1596_),
    .A(_1410_),
    .B(_1413_));
 sg13g2_buf_1 _2516_ (.A(_1596_),
    .X(_1597_));
 sg13g2_nor2_1 _2517_ (.A(net154),
    .B(_1597_),
    .Y(_1598_));
 sg13g2_buf_1 _2518_ (.A(_1598_),
    .X(_1599_));
 sg13g2_buf_1 _2519_ (.A(net110),
    .X(_1600_));
 sg13g2_o21ai_1 _2520_ (.B1(net81),
    .Y(_1601_),
    .A1(_1569_),
    .A2(_1595_));
 sg13g2_buf_1 _2521_ (.A(_1415_),
    .X(_1602_));
 sg13g2_buf_1 _2522_ (.A(net130),
    .X(_1603_));
 sg13g2_buf_1 _2523_ (.A(net109),
    .X(_1604_));
 sg13g2_buf_1 _2524_ (.A(_1555_),
    .X(_1605_));
 sg13g2_buf_1 _2525_ (.A(net163),
    .X(_1606_));
 sg13g2_nor2_2 _2526_ (.A(net84),
    .B(_1581_),
    .Y(_1607_));
 sg13g2_buf_1 _2527_ (.A(net155),
    .X(_1608_));
 sg13g2_buf_1 _2528_ (.A(_1513_),
    .X(_1609_));
 sg13g2_nor2_1 _2529_ (.A(net166),
    .B(net131),
    .Y(_1610_));
 sg13g2_buf_1 _2530_ (.A(net113),
    .X(_1611_));
 sg13g2_a221oi_1 _2531_ (.B2(_1610_),
    .C1(net79),
    .B1(net60),
    .A1(net142),
    .Y(_1612_),
    .A2(net108));
 sg13g2_nor3_1 _2532_ (.A(net159),
    .B(_1607_),
    .C(_1612_),
    .Y(_1613_));
 sg13g2_buf_1 _2533_ (.A(net85),
    .X(_1614_));
 sg13g2_buf_1 _2534_ (.A(net54),
    .X(_1615_));
 sg13g2_o21ai_1 _2535_ (.B1(net143),
    .Y(_1616_),
    .A1(_1502_),
    .A2(_1504_));
 sg13g2_buf_2 _2536_ (.A(_1616_),
    .X(_1617_));
 sg13g2_a21oi_1 _2537_ (.A1(net160),
    .A2(_1434_),
    .Y(_1618_),
    .B1(_1461_));
 sg13g2_buf_1 _2538_ (.A(_1618_),
    .X(_1619_));
 sg13g2_nor3_1 _2539_ (.A(_1442_),
    .B(_1448_),
    .C(net164),
    .Y(_1620_));
 sg13g2_buf_1 _2540_ (.A(_1620_),
    .X(_1621_));
 sg13g2_nor2_1 _2541_ (.A(net129),
    .B(net153),
    .Y(_1622_));
 sg13g2_buf_1 _2542_ (.A(_1622_),
    .X(_1623_));
 sg13g2_nor2_1 _2543_ (.A(net113),
    .B(net78),
    .Y(_1624_));
 sg13g2_buf_2 _2544_ (.A(_1624_),
    .X(_1625_));
 sg13g2_buf_1 _2545_ (.A(net167),
    .X(_1626_));
 sg13g2_a221oi_1 _2546_ (.B2(_1625_),
    .C1(net162),
    .B1(_1617_),
    .A1(net30),
    .Y(_1627_),
    .A2(_1607_));
 sg13g2_or3_1 _2547_ (.A(net80),
    .B(_1613_),
    .C(_1627_),
    .X(_1628_));
 sg13g2_buf_1 _2548_ (.A(net130),
    .X(_1629_));
 sg13g2_buf_1 _2549_ (.A(net107),
    .X(_1630_));
 sg13g2_or2_1 _2550_ (.X(_1631_),
    .B(_1418_),
    .A(_1380_));
 sg13g2_buf_1 _2551_ (.A(_1631_),
    .X(_1632_));
 sg13g2_nor2_1 _2552_ (.A(_1555_),
    .B(_1632_),
    .Y(_1633_));
 sg13g2_buf_1 _2553_ (.A(_1633_),
    .X(_1634_));
 sg13g2_nand2_2 _2554_ (.Y(_1635_),
    .A(net131),
    .B(net152));
 sg13g2_nand2_1 _2555_ (.Y(_1636_),
    .A(_1484_),
    .B(_1635_));
 sg13g2_mux2_1 _2556_ (.A0(_1517_),
    .A1(_1625_),
    .S(_1636_),
    .X(_1637_));
 sg13g2_buf_1 _2557_ (.A(_1404_),
    .X(_1638_));
 sg13g2_buf_1 _2558_ (.A(net141),
    .X(_1639_));
 sg13g2_buf_1 _2559_ (.A(_1639_),
    .X(_1640_));
 sg13g2_a21oi_1 _2560_ (.A1(net77),
    .A2(_1637_),
    .Y(_1641_),
    .B1(net106));
 sg13g2_nand2_1 _2561_ (.Y(_1642_),
    .A(_1628_),
    .B(_1641_));
 sg13g2_nand4_1 _2562_ (.B(_1559_),
    .C(_1601_),
    .A(_1523_),
    .Y(_1643_),
    .D(_1642_));
 sg13g2_buf_1 _2563_ (.A(_1392_),
    .X(_1644_));
 sg13g2_a221oi_1 _2564_ (.B2(_1590_),
    .C1(_1504_),
    .B1(_1586_),
    .A1(net155),
    .Y(_1645_),
    .A2(_1547_));
 sg13g2_buf_2 _2565_ (.A(_1645_),
    .X(_1646_));
 sg13g2_nor2_1 _2566_ (.A(net178),
    .B(_1470_),
    .Y(_1647_));
 sg13g2_a21oi_1 _2567_ (.A1(net178),
    .A2(_1470_),
    .Y(_1648_),
    .B1(_0815_));
 sg13g2_o21ai_1 _2568_ (.B1(_1436_),
    .Y(_1649_),
    .A1(_1647_),
    .A2(_1648_));
 sg13g2_or3_1 _2569_ (.A(_1436_),
    .B(_1647_),
    .C(_1648_),
    .X(_1650_));
 sg13g2_nand4_1 _2570_ (.B(_1530_),
    .C(_1649_),
    .A(_1528_),
    .Y(_1651_),
    .D(_1650_));
 sg13g2_buf_1 _2571_ (.A(_1651_),
    .X(_1652_));
 sg13g2_nor3_2 _2572_ (.A(net129),
    .B(net153),
    .C(net127),
    .Y(_1653_));
 sg13g2_a22oi_1 _2573_ (.Y(_1654_),
    .B1(_1653_),
    .B2(net85),
    .A2(_1646_),
    .A1(net113));
 sg13g2_nor2_1 _2574_ (.A(net163),
    .B(_1415_),
    .Y(_1655_));
 sg13g2_buf_1 _2575_ (.A(_1655_),
    .X(_1656_));
 sg13g2_o21ai_1 _2576_ (.B1(net105),
    .Y(_1657_),
    .A1(net166),
    .A2(_1654_));
 sg13g2_buf_2 _2577_ (.A(_1657_),
    .X(_1658_));
 sg13g2_buf_1 _2578_ (.A(net163),
    .X(_1659_));
 sg13g2_buf_1 _2579_ (.A(_1597_),
    .X(_1660_));
 sg13g2_buf_1 _2580_ (.A(_1660_),
    .X(_1661_));
 sg13g2_nand2_2 _2581_ (.Y(_1662_),
    .A(_1565_),
    .B(_1567_));
 sg13g2_a22oi_1 _2582_ (.Y(_1663_),
    .B1(_1653_),
    .B2(net54),
    .A2(_1662_),
    .A1(net112));
 sg13g2_and4_1 _2583_ (.A(net158),
    .B(_1661_),
    .C(net161),
    .D(_1663_),
    .X(_1664_));
 sg13g2_nor2_2 _2584_ (.A(_1560_),
    .B(net54),
    .Y(_1665_));
 sg13g2_nand3_1 _2585_ (.B(_1410_),
    .C(_1413_),
    .A(net163),
    .Y(_1666_));
 sg13g2_buf_2 _2586_ (.A(_1666_),
    .X(_1667_));
 sg13g2_buf_1 _2587_ (.A(_1667_),
    .X(_1668_));
 sg13g2_buf_8 _2588_ (.A(_1506_),
    .X(_1669_));
 sg13g2_buf_1 _2589_ (.A(net53),
    .X(_1670_));
 sg13g2_buf_1 _2590_ (.A(net111),
    .X(_1671_));
 sg13g2_nor3_1 _2591_ (.A(_1611_),
    .B(_1670_),
    .C(net75),
    .Y(_1672_));
 sg13g2_nor3_1 _2592_ (.A(_1665_),
    .B(net125),
    .C(_1672_),
    .Y(_1673_));
 sg13g2_nor3_1 _2593_ (.A(net129),
    .B(net153),
    .C(_1531_),
    .Y(_1674_));
 sg13g2_buf_2 _2594_ (.A(_1674_),
    .X(_1675_));
 sg13g2_nor3_2 _2595_ (.A(net84),
    .B(net85),
    .C(_1675_),
    .Y(_1676_));
 sg13g2_nor2_1 _2596_ (.A(_1055_),
    .B(net188),
    .Y(_1677_));
 sg13g2_nand3_1 _2597_ (.B(_1408_),
    .C(_1677_),
    .A(net175),
    .Y(_1678_));
 sg13g2_o21ai_1 _2598_ (.B1(_1678_),
    .Y(_1679_),
    .A1(_1381_),
    .A2(_1408_));
 sg13g2_nand3_1 _2599_ (.B(net189),
    .C(_1107_),
    .A(net175),
    .Y(_1680_));
 sg13g2_o21ai_1 _2600_ (.B1(_1680_),
    .Y(_1681_),
    .A1(net189),
    .A2(_1394_));
 sg13g2_nor2_1 _2601_ (.A(net176),
    .B(_1408_),
    .Y(_1682_));
 sg13g2_a22oi_1 _2602_ (.Y(_1683_),
    .B1(_1681_),
    .B2(_1682_),
    .A2(_1679_),
    .A1(net176));
 sg13g2_buf_2 _2603_ (.A(_1683_),
    .X(_1684_));
 sg13g2_nand3_1 _2604_ (.B(_1513_),
    .C(_1547_),
    .A(net155),
    .Y(_1685_));
 sg13g2_buf_2 _2605_ (.A(_1685_),
    .X(_1686_));
 sg13g2_nor2_1 _2606_ (.A(net79),
    .B(_1686_),
    .Y(_1687_));
 sg13g2_nor3_1 _2607_ (.A(_1676_),
    .B(_1684_),
    .C(_1687_),
    .Y(_1688_));
 sg13g2_nor2_2 _2608_ (.A(net112),
    .B(net53),
    .Y(_1689_));
 sg13g2_buf_1 _2609_ (.A(_1515_),
    .X(_1690_));
 sg13g2_buf_1 _2610_ (.A(_1632_),
    .X(_1691_));
 sg13g2_nand2_1 _2611_ (.Y(_1692_),
    .A(_1691_),
    .B(net143));
 sg13g2_nand2_1 _2612_ (.Y(_1693_),
    .A(net52),
    .B(_1692_));
 sg13g2_nand3_1 _2613_ (.B(_1410_),
    .C(_1413_),
    .A(net167),
    .Y(_1694_));
 sg13g2_buf_1 _2614_ (.A(_1694_),
    .X(_1695_));
 sg13g2_buf_1 _2615_ (.A(_1695_),
    .X(_1696_));
 sg13g2_a221oi_1 _2616_ (.B2(_1693_),
    .C1(net124),
    .B1(_1689_),
    .A1(net56),
    .Y(_1697_),
    .A2(_1665_));
 sg13g2_nor4_1 _2617_ (.A(_1664_),
    .B(_1673_),
    .C(_1688_),
    .D(_1697_),
    .Y(_1698_));
 sg13g2_a21o_1 _2618_ (.A2(_1698_),
    .A1(_1658_),
    .B1(net106),
    .X(_1699_));
 sg13g2_buf_1 _2619_ (.A(net157),
    .X(_1700_));
 sg13g2_buf_1 _2620_ (.A(net60),
    .X(_1701_));
 sg13g2_buf_1 _2621_ (.A(_1532_),
    .X(_1702_));
 sg13g2_buf_1 _2622_ (.A(net103),
    .X(_1703_));
 sg13g2_o21ai_1 _2623_ (.B1(net74),
    .Y(_1704_),
    .A1(_1700_),
    .A2(_1701_));
 sg13g2_nand3_1 _2624_ (.B(_1480_),
    .C(net143),
    .A(_1473_),
    .Y(_1705_));
 sg13g2_buf_1 _2625_ (.A(_1705_),
    .X(_1706_));
 sg13g2_buf_1 _2626_ (.A(net162),
    .X(_1707_));
 sg13g2_a221oi_1 _2627_ (.B2(_1625_),
    .C1(net156),
    .B1(net73),
    .A1(net34),
    .Y(_1708_),
    .A2(_1704_));
 sg13g2_buf_1 _2628_ (.A(_1675_),
    .X(_1709_));
 sg13g2_o21ai_1 _2629_ (.B1(net55),
    .Y(_1710_),
    .A1(net54),
    .A2(net111));
 sg13g2_nor3_1 _2630_ (.A(net129),
    .B(net153),
    .C(_1547_),
    .Y(_1711_));
 sg13g2_buf_1 _2631_ (.A(_1711_),
    .X(_1712_));
 sg13g2_a21oi_1 _2632_ (.A1(_1611_),
    .A2(net72),
    .Y(_1713_),
    .B1(net159));
 sg13g2_o21ai_1 _2633_ (.B1(_1713_),
    .Y(_1714_),
    .A1(net51),
    .A2(_1710_));
 sg13g2_nand3b_1 _2634_ (.B(_1714_),
    .C(net77),
    .Y(_1715_),
    .A_N(_1708_));
 sg13g2_buf_8 _2635_ (.A(net84),
    .X(_1716_));
 sg13g2_buf_1 _2636_ (.A(net50),
    .X(_1717_));
 sg13g2_buf_1 _2637_ (.A(net27),
    .X(_1718_));
 sg13g2_nand2_1 _2638_ (.Y(_1719_),
    .A(_1606_),
    .B(_1671_));
 sg13g2_buf_1 _2639_ (.A(net28),
    .X(_1720_));
 sg13g2_a21oi_1 _2640_ (.A1(net14),
    .A2(_1719_),
    .Y(_1721_),
    .B1(net13));
 sg13g2_nand2_1 _2641_ (.Y(_1722_),
    .A(net83),
    .B(_1482_));
 sg13g2_buf_2 _2642_ (.A(_1722_),
    .X(_1723_));
 sg13g2_o21ai_1 _2643_ (.B1(_1531_),
    .Y(_1724_),
    .A1(net129),
    .A2(net153));
 sg13g2_buf_1 _2644_ (.A(_1724_),
    .X(_1725_));
 sg13g2_nand2_1 _2645_ (.Y(_1726_),
    .A(_1407_),
    .B(_1420_));
 sg13g2_buf_1 _2646_ (.A(_1726_),
    .X(_1727_));
 sg13g2_nor2_1 _2647_ (.A(net71),
    .B(_1727_),
    .Y(_1728_));
 sg13g2_nor2_1 _2648_ (.A(_1723_),
    .B(_1728_),
    .Y(_1729_));
 sg13g2_buf_1 _2649_ (.A(net126),
    .X(_1730_));
 sg13g2_o21ai_1 _2650_ (.B1(net102),
    .Y(_1731_),
    .A1(_1721_),
    .A2(_1729_));
 sg13g2_nand3_1 _2651_ (.B(_1715_),
    .C(_1731_),
    .A(net106),
    .Y(_1732_));
 sg13g2_nand3_1 _2652_ (.B(_1699_),
    .C(_1732_),
    .A(net76),
    .Y(_1733_));
 sg13g2_nor2_1 _2653_ (.A(_0651_),
    .B(_1001_),
    .Y(_1734_));
 sg13g2_a21oi_2 _2654_ (.B1(_1386_),
    .Y(_1735_),
    .A2(_1384_),
    .A1(_1378_));
 sg13g2_and2_1 _2655_ (.A(_0530_),
    .B(_0891_),
    .X(_1736_));
 sg13g2_o21ai_1 _2656_ (.B1(_1736_),
    .Y(_1737_),
    .A1(_1734_),
    .A2(_1735_));
 sg13g2_a21o_1 _2657_ (.A2(_1384_),
    .A1(_1378_),
    .B1(_1386_),
    .X(_1738_));
 sg13g2_nor2b_1 _2658_ (.A(_0891_),
    .B_N(_0530_),
    .Y(_1739_));
 sg13g2_nand3_1 _2659_ (.B(_1738_),
    .C(_1739_),
    .A(_1387_),
    .Y(_1740_));
 sg13g2_nor2b_1 _2660_ (.A(_0530_),
    .B_N(_0891_),
    .Y(_1741_));
 sg13g2_nand3_1 _2661_ (.B(_1738_),
    .C(_1741_),
    .A(_1387_),
    .Y(_1742_));
 sg13g2_nor2_1 _2662_ (.A(net182),
    .B(_0902_),
    .Y(_1743_));
 sg13g2_o21ai_1 _2663_ (.B1(_1743_),
    .Y(_1744_),
    .A1(_1734_),
    .A2(_1735_));
 sg13g2_nand4_1 _2664_ (.B(_1740_),
    .C(_1742_),
    .A(_1737_),
    .Y(_1745_),
    .D(_1744_));
 sg13g2_buf_1 _2665_ (.A(_1745_),
    .X(_1746_));
 sg13g2_buf_1 _2666_ (.A(_1746_),
    .X(_1747_));
 sg13g2_buf_1 _2667_ (.A(net101),
    .X(_1748_));
 sg13g2_nand3_1 _2668_ (.B(_1733_),
    .C(_1748_),
    .A(_1643_),
    .Y(_1749_));
 sg13g2_nand2b_1 _2669_ (.Y(_1750_),
    .B(_0880_),
    .A_N(net198));
 sg13g2_nand2b_1 _2670_ (.Y(_1751_),
    .B(net198),
    .A_N(_0880_));
 sg13g2_buf_1 _2671_ (.A(_1751_),
    .X(_1752_));
 sg13g2_and2_1 _2672_ (.A(_1750_),
    .B(_1752_),
    .X(_1753_));
 sg13g2_buf_1 _2673_ (.A(_1753_),
    .X(_1754_));
 sg13g2_nor3_1 _2674_ (.A(_1734_),
    .B(_1735_),
    .C(_1739_),
    .Y(_1755_));
 sg13g2_nor2_1 _2675_ (.A(_1741_),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_xor2_1 _2676_ (.B(_1756_),
    .A(_1754_),
    .X(_1757_));
 sg13g2_buf_2 _2677_ (.A(_1757_),
    .X(_1758_));
 sg13g2_buf_1 _2678_ (.A(_1758_),
    .X(_1759_));
 sg13g2_xnor2_1 _2679_ (.Y(_1760_),
    .A(net186),
    .B(_1303_));
 sg13g2_buf_1 _2680_ (.A(_1760_),
    .X(_1761_));
 sg13g2_nor2_1 _2681_ (.A(net69),
    .B(net169),
    .Y(_1762_));
 sg13g2_buf_1 _2682_ (.A(_1622_),
    .X(_1763_));
 sg13g2_buf_1 _2683_ (.A(net68),
    .X(_1764_));
 sg13g2_buf_8 _2684_ (.A(net113),
    .X(_1765_));
 sg13g2_buf_1 _2685_ (.A(net67),
    .X(_1766_));
 sg13g2_nor2_1 _2686_ (.A(_1406_),
    .B(net166),
    .Y(_1767_));
 sg13g2_buf_1 _2687_ (.A(_1767_),
    .X(_1768_));
 sg13g2_buf_1 _2688_ (.A(net149),
    .X(_1769_));
 sg13g2_buf_1 _2689_ (.A(_1579_),
    .X(_1770_));
 sg13g2_buf_1 _2690_ (.A(net123),
    .X(_1771_));
 sg13g2_buf_1 _2691_ (.A(net100),
    .X(_1772_));
 sg13g2_a21oi_1 _2692_ (.A1(_1766_),
    .A2(net140),
    .Y(_1773_),
    .B1(net66));
 sg13g2_buf_1 _2693_ (.A(net57),
    .X(_1774_));
 sg13g2_buf_1 _2694_ (.A(net78),
    .X(_1775_));
 sg13g2_nand2_1 _2695_ (.Y(_1776_),
    .A(_1774_),
    .B(net47));
 sg13g2_o21ai_1 _2696_ (.B1(_1776_),
    .Y(_1777_),
    .A1(net49),
    .A2(_1773_));
 sg13g2_buf_1 _2697_ (.A(net112),
    .X(_1778_));
 sg13g2_buf_1 _2698_ (.A(net65),
    .X(_1779_));
 sg13g2_buf_1 _2699_ (.A(net29),
    .X(_1780_));
 sg13g2_and2_1 _2700_ (.A(_1649_),
    .B(_1650_),
    .X(_1781_));
 sg13g2_buf_1 _2701_ (.A(_1781_),
    .X(_1782_));
 sg13g2_nand3_1 _2702_ (.B(_1782_),
    .C(net140),
    .A(net12),
    .Y(_1783_));
 sg13g2_o21ai_1 _2703_ (.B1(_1783_),
    .Y(_1784_),
    .A1(net46),
    .A2(net140));
 sg13g2_a22oi_1 _2704_ (.Y(_1785_),
    .B1(_1784_),
    .B2(net51),
    .A2(_1777_),
    .A1(net13));
 sg13g2_nor2_2 _2705_ (.A(net58),
    .B(net111),
    .Y(_1786_));
 sg13g2_o21ai_1 _2706_ (.B1(net14),
    .Y(_1787_),
    .A1(_1709_),
    .A2(_1786_));
 sg13g2_buf_1 _2707_ (.A(_1473_),
    .X(_1788_));
 sg13g2_buf_1 _2708_ (.A(_1480_),
    .X(_1789_));
 sg13g2_a21oi_1 _2709_ (.A1(net139),
    .A2(net99),
    .Y(_1790_),
    .B1(net145));
 sg13g2_buf_1 _2710_ (.A(_1790_),
    .X(_1791_));
 sg13g2_a21oi_1 _2711_ (.A1(net158),
    .A2(net45),
    .Y(_1792_),
    .B1(net77));
 sg13g2_xnor2_1 _2712_ (.Y(_1793_),
    .A(_1385_),
    .B(_1388_));
 sg13g2_buf_2 _2713_ (.A(_1793_),
    .X(_1794_));
 sg13g2_buf_1 _2714_ (.A(net154),
    .X(_1795_));
 sg13g2_nand2_2 _2715_ (.Y(_1796_),
    .A(_1794_),
    .B(net138));
 sg13g2_a221oi_1 _2716_ (.B2(_1792_),
    .C1(_1796_),
    .B1(_1787_),
    .A1(net77),
    .Y(_1797_),
    .A2(_1785_));
 sg13g2_buf_1 _2717_ (.A(net48),
    .X(_1798_));
 sg13g2_nand3_1 _2718_ (.B(_1434_),
    .C(_1544_),
    .A(net160),
    .Y(_1799_));
 sg13g2_a21oi_2 _2719_ (.B1(net143),
    .Y(_1800_),
    .A2(_1799_),
    .A1(net99));
 sg13g2_buf_1 _2720_ (.A(_1800_),
    .X(_1801_));
 sg13g2_and2_1 _2721_ (.A(_1456_),
    .B(_1506_),
    .X(_1802_));
 sg13g2_buf_1 _2722_ (.A(_1802_),
    .X(_1803_));
 sg13g2_nor2_1 _2723_ (.A(net167),
    .B(_1597_),
    .Y(_1804_));
 sg13g2_buf_1 _2724_ (.A(_1804_),
    .X(_1805_));
 sg13g2_nor2_1 _2725_ (.A(net113),
    .B(_1515_),
    .Y(_1806_));
 sg13g2_buf_1 _2726_ (.A(_1806_),
    .X(_1807_));
 sg13g2_o21ai_1 _2727_ (.B1(net24),
    .Y(_1808_),
    .A1(net74),
    .A2(_1805_));
 sg13g2_nand2_1 _2728_ (.Y(_1809_),
    .A(_1390_),
    .B(net154));
 sg13g2_buf_2 _2729_ (.A(_1809_),
    .X(_1810_));
 sg13g2_a221oi_1 _2730_ (.B2(_1808_),
    .C1(_1810_),
    .B1(_1803_),
    .A1(net25),
    .Y(_1811_),
    .A2(net44));
 sg13g2_nand2_1 _2731_ (.Y(_1812_),
    .A(net113),
    .B(net78));
 sg13g2_buf_1 _2732_ (.A(_1812_),
    .X(_1813_));
 sg13g2_nand2_1 _2733_ (.Y(_1814_),
    .A(net84),
    .B(_1515_));
 sg13g2_buf_2 _2734_ (.A(_1814_),
    .X(_1815_));
 sg13g2_nand2_1 _2735_ (.Y(_1816_),
    .A(net23),
    .B(_1815_));
 sg13g2_buf_1 _2736_ (.A(net58),
    .X(_1817_));
 sg13g2_buf_1 _2737_ (.A(net22),
    .X(_1818_));
 sg13g2_a22oi_1 _2738_ (.Y(_1819_),
    .B1(_1816_),
    .B2(net11),
    .A2(net44),
    .A1(net25));
 sg13g2_nor2_2 _2739_ (.A(_1794_),
    .B(_1795_),
    .Y(_1820_));
 sg13g2_nand2_2 _2740_ (.Y(_1821_),
    .A(_1716_),
    .B(net71));
 sg13g2_o21ai_1 _2741_ (.B1(_1632_),
    .Y(_1822_),
    .A1(_1576_),
    .A2(_1577_));
 sg13g2_buf_1 _2742_ (.A(_1822_),
    .X(_1823_));
 sg13g2_nor3_1 _2743_ (.A(net31),
    .B(_1668_),
    .C(net137),
    .Y(_1824_));
 sg13g2_nand2_1 _2744_ (.Y(_1825_),
    .A(net175),
    .B(_1677_));
 sg13g2_o21ai_1 _2745_ (.B1(net176),
    .Y(_1826_),
    .A1(_1393_),
    .A2(_1418_));
 sg13g2_nand3_1 _2746_ (.B(_1825_),
    .C(_1826_),
    .A(_1411_),
    .Y(_1827_));
 sg13g2_nand2_1 _2747_ (.Y(_1828_),
    .A(_1410_),
    .B(_1827_));
 sg13g2_inv_1 _2748_ (.Y(_1829_),
    .A(_1828_));
 sg13g2_o21ai_1 _2749_ (.B1(_1829_),
    .Y(_1830_),
    .A1(_1821_),
    .A2(_1824_));
 sg13g2_nand3_1 _2750_ (.B(_1820_),
    .C(_1830_),
    .A(_1819_),
    .Y(_1831_));
 sg13g2_nor2_1 _2751_ (.A(_1390_),
    .B(net138),
    .Y(_1832_));
 sg13g2_buf_1 _2752_ (.A(net105),
    .X(_1833_));
 sg13g2_nand3b_1 _2753_ (.B(net11),
    .C(net64),
    .Y(_1834_),
    .A_N(_1653_));
 sg13g2_nand3_1 _2754_ (.B(net74),
    .C(net144),
    .A(net47),
    .Y(_1835_));
 sg13g2_a21oi_1 _2755_ (.A1(net145),
    .A2(_1835_),
    .Y(_1836_),
    .B1(net31));
 sg13g2_o21ai_1 _2756_ (.B1(net14),
    .Y(_1837_),
    .A1(net44),
    .A2(_1836_));
 sg13g2_nand4_1 _2757_ (.B(_1832_),
    .C(_1834_),
    .A(_1552_),
    .Y(_1838_),
    .D(_1837_));
 sg13g2_nand2_1 _2758_ (.Y(_1839_),
    .A(_1831_),
    .B(_1838_));
 sg13g2_or4_1 _2759_ (.A(net70),
    .B(_1797_),
    .C(_1811_),
    .D(_1839_),
    .X(_1840_));
 sg13g2_nand3_1 _2760_ (.B(_1762_),
    .C(_1840_),
    .A(_1749_),
    .Y(_1841_));
 sg13g2_nor2_1 _2761_ (.A(_1519_),
    .B(net111),
    .Y(_1842_));
 sg13g2_buf_2 _2762_ (.A(_1842_),
    .X(_1843_));
 sg13g2_nand2_2 _2763_ (.Y(_1844_),
    .A(_1605_),
    .B(net131));
 sg13g2_a21o_1 _2764_ (.A2(_1844_),
    .A1(net68),
    .B1(net58),
    .X(_1845_));
 sg13g2_buf_1 _2765_ (.A(_1498_),
    .X(_1846_));
 sg13g2_nor2_1 _2766_ (.A(net58),
    .B(net56),
    .Y(_1847_));
 sg13g2_a221oi_1 _2767_ (.B2(net156),
    .C1(net14),
    .B1(_1847_),
    .A1(net11),
    .Y(_1848_),
    .A2(net97));
 sg13g2_a21oi_1 _2768_ (.A1(_1843_),
    .A2(_1845_),
    .Y(_1849_),
    .B1(_1848_));
 sg13g2_nand2_1 _2769_ (.Y(_1850_),
    .A(net75),
    .B(_1634_));
 sg13g2_a21oi_1 _2770_ (.A1(_1676_),
    .A2(_1850_),
    .Y(_1851_),
    .B1(net104));
 sg13g2_a21o_1 _2771_ (.A2(_1590_),
    .A1(_1586_),
    .B1(net163),
    .X(_1852_));
 sg13g2_nand2_1 _2772_ (.Y(_1853_),
    .A(net131),
    .B(_1767_));
 sg13g2_o21ai_1 _2773_ (.B1(_1483_),
    .Y(_1854_),
    .A1(net68),
    .A2(_1853_));
 sg13g2_a21o_1 _2774_ (.A2(_1854_),
    .A1(_1852_),
    .B1(net48),
    .X(_1855_));
 sg13g2_buf_1 _2775_ (.A(net141),
    .X(_1856_));
 sg13g2_a21oi_1 _2776_ (.A1(_1851_),
    .A2(_1855_),
    .Y(_1857_),
    .B1(net122));
 sg13g2_o21ai_1 _2777_ (.B1(_1857_),
    .Y(_1858_),
    .A1(net77),
    .A2(_1849_));
 sg13g2_buf_1 _2778_ (.A(net152),
    .X(_1859_));
 sg13g2_buf_8 _2779_ (.A(net131),
    .X(_1860_));
 sg13g2_nor2_2 _2780_ (.A(net96),
    .B(net149),
    .Y(_1861_));
 sg13g2_o21ai_1 _2781_ (.B1(_1687_),
    .Y(_1862_),
    .A1(net136),
    .A2(_1861_));
 sg13g2_a21oi_2 _2782_ (.B1(net157),
    .Y(_1863_),
    .A2(_1530_),
    .A1(_1528_));
 sg13g2_buf_1 _2783_ (.A(net52),
    .X(_1864_));
 sg13g2_o21ai_1 _2784_ (.B1(net21),
    .Y(_1865_),
    .A1(net162),
    .A2(_1863_));
 sg13g2_nand2_1 _2785_ (.Y(_1866_),
    .A(net113),
    .B(net53));
 sg13g2_a21o_1 _2786_ (.A2(_1865_),
    .A1(_1635_),
    .B1(_1866_),
    .X(_1867_));
 sg13g2_nand3_1 _2787_ (.B(_1862_),
    .C(_1867_),
    .A(_1600_),
    .Y(_1868_));
 sg13g2_buf_1 _2788_ (.A(net78),
    .X(_1869_));
 sg13g2_o21ai_1 _2789_ (.B1(_1689_),
    .Y(_1870_),
    .A1(net43),
    .A2(_1861_));
 sg13g2_nor2_1 _2790_ (.A(net109),
    .B(_1676_),
    .Y(_1871_));
 sg13g2_buf_1 _2791_ (.A(net138),
    .X(_1872_));
 sg13g2_a21oi_1 _2792_ (.A1(_1870_),
    .A2(_1871_),
    .Y(_1873_),
    .B1(net121));
 sg13g2_a21oi_1 _2793_ (.A1(_1868_),
    .A2(_1873_),
    .Y(_1874_),
    .B1(_1644_));
 sg13g2_buf_1 _2794_ (.A(_1416_),
    .X(_1875_));
 sg13g2_nand2_1 _2795_ (.Y(_1876_),
    .A(_1391_),
    .B(net95));
 sg13g2_o21ai_1 _2796_ (.B1(net13),
    .Y(_1877_),
    .A1(_1700_),
    .A2(_1876_));
 sg13g2_a21oi_1 _2797_ (.A1(net66),
    .A2(_1877_),
    .Y(_1878_),
    .B1(net23));
 sg13g2_and2_1 _2798_ (.A(_1506_),
    .B(_1498_),
    .X(_1879_));
 sg13g2_buf_1 _2799_ (.A(_1879_),
    .X(_1880_));
 sg13g2_nor2_1 _2800_ (.A(_1880_),
    .B(_1876_),
    .Y(_1881_));
 sg13g2_buf_1 _2801_ (.A(_1794_),
    .X(_1882_));
 sg13g2_nor2_1 _2802_ (.A(net176),
    .B(_1411_),
    .Y(_1883_));
 sg13g2_nand3_1 _2803_ (.B(_1380_),
    .C(_1408_),
    .A(net189),
    .Y(_1884_));
 sg13g2_o21ai_1 _2804_ (.B1(_1884_),
    .Y(_1885_),
    .A1(_1408_),
    .A2(_1825_));
 sg13g2_a22oi_1 _2805_ (.Y(_1886_),
    .B1(_1885_),
    .B2(net176),
    .A2(_1883_),
    .A1(_1681_));
 sg13g2_buf_1 _2806_ (.A(_1886_),
    .X(_1887_));
 sg13g2_nor3_2 _2807_ (.A(_1502_),
    .B(_1504_),
    .C(net145),
    .Y(_1888_));
 sg13g2_nor3_1 _2808_ (.A(net120),
    .B(net148),
    .C(_1888_),
    .Y(_1889_));
 sg13g2_nor2_1 _2809_ (.A(_1881_),
    .B(_1889_),
    .Y(_1890_));
 sg13g2_o21ai_1 _2810_ (.B1(net66),
    .Y(_1891_),
    .A1(net104),
    .A2(net35));
 sg13g2_a21o_1 _2811_ (.A2(_1413_),
    .A1(_1410_),
    .B1(net167),
    .X(_1892_));
 sg13g2_buf_1 _2812_ (.A(_1892_),
    .X(_1893_));
 sg13g2_nand2_1 _2813_ (.Y(_1894_),
    .A(net135),
    .B(net148));
 sg13g2_a221oi_1 _2814_ (.B2(_1891_),
    .C1(_1894_),
    .B1(net34),
    .A1(net11),
    .Y(_1895_),
    .A2(net97));
 sg13g2_o21ai_1 _2815_ (.B1(_1644_),
    .Y(_1896_),
    .A1(net106),
    .A2(_1895_));
 sg13g2_o21ai_1 _2816_ (.B1(_1896_),
    .Y(_1897_),
    .A1(_1878_),
    .A2(_1890_));
 sg13g2_nand2_1 _2817_ (.Y(_1898_),
    .A(_1480_),
    .B(_1799_));
 sg13g2_buf_2 _2818_ (.A(_1898_),
    .X(_1899_));
 sg13g2_buf_1 _2819_ (.A(_1899_),
    .X(_1900_));
 sg13g2_nand2_1 _2820_ (.Y(_1901_),
    .A(_1779_),
    .B(net73));
 sg13g2_a22oi_1 _2821_ (.Y(_1902_),
    .B1(_1901_),
    .B2(net49),
    .A2(net137),
    .A1(net42));
 sg13g2_o21ai_1 _2822_ (.B1(_1456_),
    .Y(_1903_),
    .A1(net161),
    .A2(_1686_));
 sg13g2_nand2_1 _2823_ (.Y(_1904_),
    .A(net74),
    .B(_1903_));
 sg13g2_a21oi_1 _2824_ (.A1(_1902_),
    .A2(_1904_),
    .Y(_1905_),
    .B1(net135));
 sg13g2_buf_1 _2825_ (.A(net85),
    .X(_1906_));
 sg13g2_nand2_1 _2826_ (.Y(_1907_),
    .A(net41),
    .B(_1607_));
 sg13g2_nand2_2 _2827_ (.Y(_1908_),
    .A(_1536_),
    .B(_1538_));
 sg13g2_nor3_1 _2828_ (.A(_1491_),
    .B(_1515_),
    .C(_1579_),
    .Y(_1909_));
 sg13g2_buf_1 _2829_ (.A(_1909_),
    .X(_1910_));
 sg13g2_o21ai_1 _2830_ (.B1(net29),
    .Y(_1911_),
    .A1(_1908_),
    .A2(net20));
 sg13g2_nand2b_1 _2831_ (.Y(_1912_),
    .B(_1625_),
    .A_N(_1861_));
 sg13g2_nand4_1 _2832_ (.B(_1907_),
    .C(_1911_),
    .A(net107),
    .Y(_1913_),
    .D(_1912_));
 sg13g2_buf_1 _2833_ (.A(net121),
    .X(_1914_));
 sg13g2_nand2_1 _2834_ (.Y(_1915_),
    .A(_1765_),
    .B(net103));
 sg13g2_buf_1 _2835_ (.A(_1662_),
    .X(_1916_));
 sg13g2_buf_1 _2836_ (.A(net144),
    .X(_1917_));
 sg13g2_a221oi_1 _2837_ (.B2(net93),
    .C1(net119),
    .B1(_1915_),
    .A1(net34),
    .Y(_1918_),
    .A2(net73));
 sg13g2_nor2_1 _2838_ (.A(net94),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_nand3b_1 _2839_ (.B(_1913_),
    .C(_1919_),
    .Y(_1920_),
    .A_N(_1905_));
 sg13g2_nor2_1 _2840_ (.A(net101),
    .B(net169),
    .Y(_1921_));
 sg13g2_nand2_1 _2841_ (.Y(_1922_),
    .A(net69),
    .B(_1921_));
 sg13g2_a221oi_1 _2842_ (.B2(_1920_),
    .C1(_1922_),
    .B1(_1897_),
    .A1(_1858_),
    .Y(_1923_),
    .A2(_1874_));
 sg13g2_buf_1 _2843_ (.A(_1882_),
    .X(_1924_));
 sg13g2_nor2_2 _2844_ (.A(net123),
    .B(net152),
    .Y(_1925_));
 sg13g2_buf_1 _2845_ (.A(_1515_),
    .X(_1926_));
 sg13g2_buf_1 _2846_ (.A(net40),
    .X(_1927_));
 sg13g2_o21ai_1 _2847_ (.B1(net19),
    .Y(_1928_),
    .A1(net33),
    .A2(_1925_));
 sg13g2_o21ai_1 _2848_ (.B1(net25),
    .Y(_1929_),
    .A1(net150),
    .A2(net44));
 sg13g2_nand2_1 _2849_ (.Y(_1930_),
    .A(net21),
    .B(_1859_));
 sg13g2_o21ai_1 _2850_ (.B1(net66),
    .Y(_1931_),
    .A1(_1782_),
    .A2(_1727_));
 sg13g2_nand3_1 _2851_ (.B(_1930_),
    .C(_1931_),
    .A(net12),
    .Y(_1932_));
 sg13g2_and4_1 _2852_ (.A(net81),
    .B(_1928_),
    .C(_1929_),
    .D(_1932_),
    .X(_1933_));
 sg13g2_nor3_1 _2853_ (.A(net92),
    .B(_1748_),
    .C(_1933_),
    .Y(_1934_));
 sg13g2_nand2_2 _2854_ (.Y(_1935_),
    .A(_1404_),
    .B(_1602_));
 sg13g2_nor2_2 _2855_ (.A(net54),
    .B(net127),
    .Y(_1936_));
 sg13g2_nand2_1 _2856_ (.Y(_1937_),
    .A(net67),
    .B(net54));
 sg13g2_buf_2 _2857_ (.A(_1937_),
    .X(_1938_));
 sg13g2_nor3_1 _2858_ (.A(net158),
    .B(net49),
    .C(_1938_),
    .Y(_1939_));
 sg13g2_nor2_1 _2859_ (.A(net128),
    .B(_1629_),
    .Y(_1940_));
 sg13g2_o21ai_1 _2860_ (.B1(_1940_),
    .Y(_1941_),
    .A1(_1936_),
    .A2(_1939_));
 sg13g2_nand3_1 _2861_ (.B(_1819_),
    .C(_1941_),
    .A(_1935_),
    .Y(_1942_));
 sg13g2_and4_1 _2862_ (.A(_1737_),
    .B(_1740_),
    .C(_1742_),
    .D(_1744_),
    .X(_1943_));
 sg13g2_buf_1 _2863_ (.A(_1943_),
    .X(_1944_));
 sg13g2_buf_1 _2864_ (.A(net118),
    .X(_1945_));
 sg13g2_nand2_1 _2865_ (.Y(_1946_),
    .A(_1555_),
    .B(net157));
 sg13g2_buf_1 _2866_ (.A(_1946_),
    .X(_1947_));
 sg13g2_nand2_1 _2867_ (.Y(_1948_),
    .A(net150),
    .B(net134));
 sg13g2_o21ai_1 _2868_ (.B1(net104),
    .Y(_1949_),
    .A1(_1663_),
    .A2(_1948_));
 sg13g2_o21ai_1 _2869_ (.B1(_1769_),
    .Y(_1950_),
    .A1(_1676_),
    .A2(_1687_));
 sg13g2_nor2b_1 _2870_ (.A(_1949_),
    .B_N(_1950_),
    .Y(_1951_));
 sg13g2_nor4_1 _2871_ (.A(_1673_),
    .B(_1697_),
    .C(_1810_),
    .D(_1951_),
    .Y(_1952_));
 sg13g2_a21oi_2 _2872_ (.B1(net157),
    .Y(_1953_),
    .A2(_1789_),
    .A1(net139));
 sg13g2_or2_1 _2873_ (.X(_1954_),
    .B(_1953_),
    .A(_1582_));
 sg13g2_a22oi_1 _2874_ (.Y(_1955_),
    .B1(_1954_),
    .B2(net46),
    .A2(_1936_),
    .A1(net161));
 sg13g2_a21oi_1 _2875_ (.A1(_1776_),
    .A2(_1955_),
    .Y(_1956_),
    .B1(net156));
 sg13g2_nand2_1 _2876_ (.Y(_1957_),
    .A(net132),
    .B(net110));
 sg13g2_nor2b_1 _2877_ (.A(_1957_),
    .B_N(_1714_),
    .Y(_1958_));
 sg13g2_nor2b_1 _2878_ (.A(_1956_),
    .B_N(_1958_),
    .Y(_1959_));
 sg13g2_o21ai_1 _2879_ (.B1(_1719_),
    .Y(_1960_),
    .A1(net35),
    .A2(_1728_));
 sg13g2_nor2_1 _2880_ (.A(net123),
    .B(net134),
    .Y(_1961_));
 sg13g2_a21oi_1 _2881_ (.A1(_1927_),
    .A2(_1961_),
    .Y(_1962_),
    .B1(net15));
 sg13g2_a22oi_1 _2882_ (.Y(_1963_),
    .B1(_1962_),
    .B2(_1818_),
    .A2(_1960_),
    .A1(_1718_));
 sg13g2_nand2_1 _2883_ (.Y(_1964_),
    .A(_1404_),
    .B(_1597_));
 sg13g2_buf_1 _2884_ (.A(_1964_),
    .X(_1965_));
 sg13g2_nor3_1 _2885_ (.A(_1924_),
    .B(_1963_),
    .C(_1965_),
    .Y(_1966_));
 sg13g2_nor4_1 _2886_ (.A(_1945_),
    .B(_1952_),
    .C(_1959_),
    .D(_1966_),
    .Y(_1967_));
 sg13g2_buf_1 _2887_ (.A(net53),
    .X(_1968_));
 sg13g2_nand3_1 _2888_ (.B(net18),
    .C(_1961_),
    .A(net32),
    .Y(_1969_));
 sg13g2_nand2_1 _2889_ (.Y(_1970_),
    .A(net167),
    .B(net96));
 sg13g2_nand3_1 _2890_ (.B(net41),
    .C(_1970_),
    .A(net65),
    .Y(_1971_));
 sg13g2_a21oi_1 _2891_ (.A1(_1969_),
    .A2(_1971_),
    .Y(_1972_),
    .B1(net21));
 sg13g2_nand2_1 _2892_ (.Y(_1973_),
    .A(_1817_),
    .B(_1823_));
 sg13g2_a21oi_1 _2893_ (.A1(_1970_),
    .A2(_1973_),
    .Y(_1974_),
    .B1(_1815_));
 sg13g2_buf_1 _2894_ (.A(net109),
    .X(_1975_));
 sg13g2_o21ai_1 _2895_ (.B1(net63),
    .Y(_1976_),
    .A1(_1972_),
    .A2(_1974_));
 sg13g2_nand3_1 _2896_ (.B(_1628_),
    .C(_1976_),
    .A(net94),
    .Y(_1977_));
 sg13g2_buf_1 _2897_ (.A(net134),
    .X(_1978_));
 sg13g2_nor3_1 _2898_ (.A(_1764_),
    .B(_1594_),
    .C(net117),
    .Y(_1979_));
 sg13g2_nor3_1 _2899_ (.A(net15),
    .B(_1550_),
    .C(_1979_),
    .Y(_1980_));
 sg13g2_buf_1 _2900_ (.A(_1582_),
    .X(_1981_));
 sg13g2_nor2_2 _2901_ (.A(_1614_),
    .B(net111),
    .Y(_1982_));
 sg13g2_a221oi_1 _2902_ (.B2(net13),
    .C1(_1798_),
    .B1(net140),
    .A1(net17),
    .Y(_1983_),
    .A2(_1982_));
 sg13g2_nor2_1 _2903_ (.A(net154),
    .B(_1415_),
    .Y(_1984_));
 sg13g2_buf_2 _2904_ (.A(_1984_),
    .X(_0078_));
 sg13g2_o21ai_1 _2905_ (.B1(_0078_),
    .Y(_0079_),
    .A1(_1980_),
    .A2(_1983_));
 sg13g2_o21ai_1 _2906_ (.B1(net21),
    .Y(_0080_),
    .A1(_1766_),
    .A2(_1861_));
 sg13g2_and3_1 _2907_ (.X(_0081_),
    .A(_1818_),
    .B(_1534_),
    .C(_0080_));
 sg13g2_o21ai_1 _2908_ (.B1(net81),
    .Y(_0082_),
    .A1(_1569_),
    .A2(_0081_));
 sg13g2_nand4_1 _2909_ (.B(_1977_),
    .C(_0079_),
    .A(_1924_),
    .Y(_0083_),
    .D(_0082_));
 sg13g2_nand3_1 _2910_ (.B(net99),
    .C(net144),
    .A(net139),
    .Y(_0084_));
 sg13g2_nor2_1 _2911_ (.A(net24),
    .B(_0084_),
    .Y(_0085_));
 sg13g2_nand3_1 _2912_ (.B(_1480_),
    .C(net131),
    .A(net139),
    .Y(_0086_));
 sg13g2_buf_2 _2913_ (.A(_0086_),
    .X(_0087_));
 sg13g2_a21oi_1 _2914_ (.A1(net24),
    .A2(_0087_),
    .Y(_0088_),
    .B1(net45));
 sg13g2_nor2b_1 _2915_ (.A(_0085_),
    .B_N(_0088_),
    .Y(_0089_));
 sg13g2_buf_1 _2916_ (.A(net144),
    .X(_0090_));
 sg13g2_a21oi_1 _2917_ (.A1(net116),
    .A2(net45),
    .Y(_0091_),
    .B1(_1796_));
 sg13g2_a22oi_1 _2918_ (.Y(_0092_),
    .B1(_0091_),
    .B2(_1787_),
    .A2(_0089_),
    .A1(_1832_));
 sg13g2_xor2_1 _2919_ (.B(_1303_),
    .A(_1215_),
    .X(_0093_));
 sg13g2_buf_1 _2920_ (.A(_0093_),
    .X(_0094_));
 sg13g2_nor2_1 _2921_ (.A(_1758_),
    .B(net168),
    .Y(_0095_));
 sg13g2_o21ai_1 _2922_ (.B1(_0095_),
    .Y(_0096_),
    .A1(net70),
    .A2(_0092_));
 sg13g2_a221oi_1 _2923_ (.B2(_0083_),
    .C1(_0096_),
    .B1(_1967_),
    .A1(_1934_),
    .Y(_0097_),
    .A2(_1942_));
 sg13g2_nand2_1 _2924_ (.Y(_0098_),
    .A(net69),
    .B(net169));
 sg13g2_buf_1 _2925_ (.A(net71),
    .X(_0099_));
 sg13g2_nand2_2 _2926_ (.Y(_0100_),
    .A(net67),
    .B(_1675_));
 sg13g2_a21oi_1 _2927_ (.A1(net30),
    .A2(net148),
    .Y(_0101_),
    .B1(_1712_));
 sg13g2_nand2_1 _2928_ (.Y(_0102_),
    .A(net15),
    .B(_0101_));
 sg13g2_nand3_1 _2929_ (.B(_0100_),
    .C(_0102_),
    .A(net39),
    .Y(_0103_));
 sg13g2_nand3_1 _2930_ (.B(net78),
    .C(_0087_),
    .A(net112),
    .Y(_0104_));
 sg13g2_buf_2 _2931_ (.A(_0104_),
    .X(_0105_));
 sg13g2_and2_1 _2932_ (.A(net39),
    .B(_0105_),
    .X(_0106_));
 sg13g2_nand2_1 _2933_ (.Y(_0107_),
    .A(net17),
    .B(net33));
 sg13g2_a21oi_1 _2934_ (.A1(_0106_),
    .A2(_0107_),
    .Y(_0108_),
    .B1(_1975_));
 sg13g2_a21oi_1 _2935_ (.A1(net98),
    .A2(_0103_),
    .Y(_0109_),
    .B1(_0108_));
 sg13g2_nor2_1 _2936_ (.A(_1605_),
    .B(_1597_),
    .Y(_0110_));
 sg13g2_buf_1 _2937_ (.A(_0110_),
    .X(_0111_));
 sg13g2_o21ai_1 _2938_ (.B1(net19),
    .Y(_0112_),
    .A1(net74),
    .A2(_1525_));
 sg13g2_nand2_1 _2939_ (.Y(_0113_),
    .A(_0105_),
    .B(_0112_));
 sg13g2_a21oi_1 _2940_ (.A1(net89),
    .A2(_0113_),
    .Y(_0114_),
    .B1(_1640_));
 sg13g2_nor2_1 _2941_ (.A(net50),
    .B(net145),
    .Y(_0115_));
 sg13g2_inv_1 _2942_ (.Y(_0116_),
    .A(_1547_));
 sg13g2_nand3_1 _2943_ (.B(_1513_),
    .C(_0116_),
    .A(net155),
    .Y(_0117_));
 sg13g2_buf_1 _2944_ (.A(_0117_),
    .X(_0118_));
 sg13g2_nor2_1 _2945_ (.A(net46),
    .B(_0118_),
    .Y(_0119_));
 sg13g2_o21ai_1 _2946_ (.B1(net102),
    .Y(_0120_),
    .A1(_0115_),
    .A2(_0119_));
 sg13g2_nor3_1 _2947_ (.A(net129),
    .B(net153),
    .C(net143),
    .Y(_0121_));
 sg13g2_buf_1 _2948_ (.A(_0121_),
    .X(_0122_));
 sg13g2_o21ai_1 _2949_ (.B1(net11),
    .Y(_0123_),
    .A1(net62),
    .A2(_0115_));
 sg13g2_nor2_1 _2950_ (.A(net89),
    .B(net20),
    .Y(_0124_));
 sg13g2_nand3_1 _2951_ (.B(_0123_),
    .C(_0124_),
    .A(_0120_),
    .Y(_0125_));
 sg13g2_nor4_1 _2952_ (.A(net129),
    .B(net153),
    .C(_1547_),
    .D(net143),
    .Y(_0126_));
 sg13g2_buf_2 _2953_ (.A(_0126_),
    .X(_0127_));
 sg13g2_o21ai_1 _2954_ (.B1(_1846_),
    .Y(_0128_),
    .A1(net25),
    .A2(_0127_));
 sg13g2_a21oi_1 _2955_ (.A1(_0111_),
    .A2(_0128_),
    .Y(_0129_),
    .B1(_1914_));
 sg13g2_a221oi_1 _2956_ (.B2(_0129_),
    .C1(net76),
    .B1(_0125_),
    .A1(_0109_),
    .Y(_0130_),
    .A2(_0114_));
 sg13g2_nand2_2 _2957_ (.Y(_0131_),
    .A(_1583_),
    .B(_1662_));
 sg13g2_nand3_1 _2958_ (.B(_0100_),
    .C(_0131_),
    .A(net39),
    .Y(_0132_));
 sg13g2_nand2_1 _2959_ (.Y(_0133_),
    .A(net15),
    .B(net62));
 sg13g2_a22oi_1 _2960_ (.Y(_0134_),
    .B1(_0133_),
    .B2(net11),
    .A2(_1786_),
    .A1(net23));
 sg13g2_a21oi_1 _2961_ (.A1(_1600_),
    .A2(_0132_),
    .Y(_0135_),
    .B1(_0134_));
 sg13g2_nor2_1 _2962_ (.A(net92),
    .B(_0135_),
    .Y(_0136_));
 sg13g2_nor4_1 _2963_ (.A(net91),
    .B(_0098_),
    .C(_0130_),
    .D(_0136_),
    .Y(_0137_));
 sg13g2_nor2_1 _2964_ (.A(net39),
    .B(_1521_),
    .Y(_0138_));
 sg13g2_o21ai_1 _2965_ (.B1(net166),
    .Y(_0139_),
    .A1(_1576_),
    .A2(_1577_));
 sg13g2_nand3_1 _2966_ (.B(net108),
    .C(_0139_),
    .A(net142),
    .Y(_0140_));
 sg13g2_nand2_1 _2967_ (.Y(_0141_),
    .A(net35),
    .B(_0140_));
 sg13g2_a21oi_1 _2968_ (.A1(net34),
    .A2(net73),
    .Y(_0142_),
    .B1(net119));
 sg13g2_o21ai_1 _2969_ (.B1(_0142_),
    .Y(_0143_),
    .A1(_0138_),
    .A2(_0141_));
 sg13g2_nand4_1 _2970_ (.B(_1593_),
    .C(_1907_),
    .A(_1875_),
    .Y(_0144_),
    .D(_1911_));
 sg13g2_nand4_1 _2971_ (.B(_1913_),
    .C(_0143_),
    .A(_1640_),
    .Y(_0145_),
    .D(_0144_));
 sg13g2_a21oi_1 _2972_ (.A1(net161),
    .A2(net59),
    .Y(_0146_),
    .B1(net145));
 sg13g2_o21ai_1 _2973_ (.B1(net22),
    .Y(_0147_),
    .A1(_0122_),
    .A2(_0146_));
 sg13g2_nor2_1 _2974_ (.A(_1917_),
    .B(net20),
    .Y(_0148_));
 sg13g2_buf_1 _2975_ (.A(net79),
    .X(_0149_));
 sg13g2_a21oi_1 _2976_ (.A1(net38),
    .A2(_1550_),
    .Y(_0150_),
    .B1(net64));
 sg13g2_nand2_1 _2977_ (.Y(_0151_),
    .A(_1507_),
    .B(_1498_));
 sg13g2_a221oi_1 _2978_ (.B2(_0151_),
    .C1(net122),
    .B1(_0150_),
    .A1(_0147_),
    .Y(_0152_),
    .A2(_0148_));
 sg13g2_nor2_1 _2979_ (.A(net92),
    .B(_0152_),
    .Y(_0153_));
 sg13g2_a21oi_1 _2980_ (.A1(_1815_),
    .A2(_1907_),
    .Y(_0154_),
    .B1(net150));
 sg13g2_a22oi_1 _2981_ (.Y(_0155_),
    .B1(_0151_),
    .B2(net38),
    .A2(_1845_),
    .A1(_1843_));
 sg13g2_or2_1 _2982_ (.X(_0156_),
    .B(_0155_),
    .A(net80));
 sg13g2_o21ai_1 _2983_ (.B1(_1857_),
    .Y(_0157_),
    .A1(_0154_),
    .A2(_0156_));
 sg13g2_o21ai_1 _2984_ (.B1(_1629_),
    .Y(_0158_),
    .A1(_1663_),
    .A2(_1769_));
 sg13g2_nor2_1 _2985_ (.A(net32),
    .B(_0087_),
    .Y(_0159_));
 sg13g2_o21ai_1 _2986_ (.B1(_1859_),
    .Y(_0160_),
    .A1(_1687_),
    .A2(_0159_));
 sg13g2_nand2b_1 _2987_ (.Y(_0161_),
    .B(_0160_),
    .A_N(_0158_));
 sg13g2_buf_1 _2988_ (.A(net132),
    .X(_0162_));
 sg13g2_a21oi_1 _2989_ (.A1(_1873_),
    .A2(_0161_),
    .Y(_0163_),
    .B1(_0162_));
 sg13g2_nand3_1 _2990_ (.B(_1759_),
    .C(net169),
    .A(net91),
    .Y(_0164_));
 sg13g2_a221oi_1 _2991_ (.B2(_0163_),
    .C1(_0164_),
    .B1(_0157_),
    .A1(_0145_),
    .Y(_0165_),
    .A2(_0153_));
 sg13g2_nand3_1 _2992_ (.B(_1758_),
    .C(net168),
    .A(_1746_),
    .Y(_0166_));
 sg13g2_and2_1 _2993_ (.A(net68),
    .B(_1635_),
    .X(_0167_));
 sg13g2_nand2b_1 _2994_ (.Y(_0168_),
    .B(_1525_),
    .A_N(_0167_));
 sg13g2_nor3_2 _2995_ (.A(_1502_),
    .B(_1504_),
    .C(net123),
    .Y(_0169_));
 sg13g2_nor2_1 _2996_ (.A(net32),
    .B(_0169_),
    .Y(_0170_));
 sg13g2_o21ai_1 _2997_ (.B1(net156),
    .Y(_0171_),
    .A1(_1927_),
    .A2(_0170_));
 sg13g2_a22oi_1 _2998_ (.Y(_0172_),
    .B1(_0171_),
    .B2(net77),
    .A2(_0106_),
    .A1(_0168_));
 sg13g2_nor2_1 _2999_ (.A(_1421_),
    .B(_1780_),
    .Y(_0173_));
 sg13g2_o21ai_1 _3000_ (.B1(net14),
    .Y(_0174_),
    .A1(net93),
    .A2(_0173_));
 sg13g2_a21oi_1 _3001_ (.A1(_0106_),
    .A2(_0174_),
    .Y(_0175_),
    .B1(net125));
 sg13g2_nor4_1 _3002_ (.A(_1796_),
    .B(_0166_),
    .C(_0172_),
    .D(_0175_),
    .Y(_0176_));
 sg13g2_nand2_1 _3003_ (.Y(_0177_),
    .A(_1794_),
    .B(_1638_));
 sg13g2_o21ai_1 _3004_ (.B1(net66),
    .Y(_0178_),
    .A1(net48),
    .A2(_1557_));
 sg13g2_a22oi_1 _3005_ (.Y(_0179_),
    .B1(net72),
    .B2(_0178_),
    .A2(_1846_),
    .A1(net46));
 sg13g2_nor3_1 _3006_ (.A(_0177_),
    .B(_0166_),
    .C(_0179_),
    .Y(_0180_));
 sg13g2_nand2b_1 _3007_ (.Y(_0181_),
    .B(_1425_),
    .A_N(_1426_));
 sg13g2_xnor2_1 _3008_ (.Y(_0182_),
    .A(_1572_),
    .B(_0181_));
 sg13g2_buf_2 _3009_ (.A(_0182_),
    .X(_0183_));
 sg13g2_xnor2_1 _3010_ (.Y(_0184_),
    .A(_1301_),
    .B(_1440_));
 sg13g2_buf_2 _3011_ (.A(_0184_),
    .X(_0185_));
 sg13g2_xnor2_1 _3012_ (.Y(_0186_),
    .A(_1197_),
    .B(_0185_));
 sg13g2_o21ai_1 _3013_ (.B1(net26),
    .Y(_0187_),
    .A1(net44),
    .A2(_1880_));
 sg13g2_nor2_1 _3014_ (.A(net90),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_buf_1 _3015_ (.A(net123),
    .X(_0189_));
 sg13g2_nor2_2 _3016_ (.A(_1492_),
    .B(net78),
    .Y(_0190_));
 sg13g2_o21ai_1 _3017_ (.B1(_0190_),
    .Y(_0191_),
    .A1(net154),
    .A2(net87));
 sg13g2_nor2_1 _3018_ (.A(_1404_),
    .B(_1498_),
    .Y(_0192_));
 sg13g2_o21ai_1 _3019_ (.B1(net18),
    .Y(_0193_),
    .A1(net20),
    .A2(_0192_));
 sg13g2_and4_1 _3020_ (.A(_0088_),
    .B(net90),
    .C(_0191_),
    .D(_0193_),
    .X(_0194_));
 sg13g2_o21ai_1 _3021_ (.B1(_0078_),
    .Y(_0195_),
    .A1(net47),
    .A2(_1925_));
 sg13g2_o21ai_1 _3022_ (.B1(_1391_),
    .Y(_0196_),
    .A1(_1938_),
    .A2(_0195_));
 sg13g2_nor4_1 _3023_ (.A(_0166_),
    .B(_0188_),
    .C(_0194_),
    .D(_0196_),
    .Y(_0197_));
 sg13g2_or4_1 _3024_ (.A(_0180_),
    .B(_0183_),
    .C(_0186_),
    .D(_0197_),
    .X(_0198_));
 sg13g2_or3_1 _3025_ (.A(_0165_),
    .B(_0176_),
    .C(_0198_),
    .X(_0199_));
 sg13g2_nor4_1 _3026_ (.A(_1923_),
    .B(_0097_),
    .C(_0137_),
    .D(_0199_),
    .Y(_0200_));
 sg13g2_and2_1 _3027_ (.A(_1480_),
    .B(_1799_),
    .X(_0201_));
 sg13g2_buf_2 _3028_ (.A(_0201_),
    .X(_0202_));
 sg13g2_nor2_1 _3029_ (.A(net60),
    .B(_1768_),
    .Y(_0203_));
 sg13g2_nand2_1 _3030_ (.Y(_0204_),
    .A(net51),
    .B(_0203_));
 sg13g2_nand3_1 _3031_ (.B(_0202_),
    .C(_0204_),
    .A(_1776_),
    .Y(_0205_));
 sg13g2_nor2_1 _3032_ (.A(net96),
    .B(net144),
    .Y(_0206_));
 sg13g2_buf_1 _3033_ (.A(net112),
    .X(_0207_));
 sg13g2_a21oi_1 _3034_ (.A1(_0207_),
    .A2(net73),
    .Y(_0208_),
    .B1(net148));
 sg13g2_o21ai_1 _3035_ (.B1(net49),
    .Y(_0209_),
    .A1(_0206_),
    .A2(_0208_));
 sg13g2_o21ai_1 _3036_ (.B1(_0209_),
    .Y(_0210_),
    .A1(_0202_),
    .A2(net148));
 sg13g2_a21oi_1 _3037_ (.A1(net155),
    .A2(_1513_),
    .Y(_0211_),
    .B1(_1863_));
 sg13g2_o21ai_1 _3038_ (.B1(_1581_),
    .Y(_0212_),
    .A1(net112),
    .A2(_0211_));
 sg13g2_nor3_1 _3039_ (.A(net109),
    .B(net61),
    .C(net39),
    .Y(_0213_));
 sg13g2_a21o_1 _3040_ (.A2(_0212_),
    .A1(net107),
    .B1(_0213_),
    .X(_0214_));
 sg13g2_o21ai_1 _3041_ (.B1(net85),
    .Y(_0215_),
    .A1(net83),
    .A2(_1591_));
 sg13g2_buf_1 _3042_ (.A(_0215_),
    .X(_0216_));
 sg13g2_nand2_1 _3043_ (.Y(_0217_),
    .A(net156),
    .B(_0216_));
 sg13g2_o21ai_1 _3044_ (.B1(net100),
    .Y(_0218_),
    .A1(net157),
    .A2(_1667_));
 sg13g2_buf_1 _3045_ (.A(net55),
    .X(_0219_));
 sg13g2_a221oi_1 _3046_ (.B2(_0218_),
    .C1(net16),
    .B1(net42),
    .A1(net43),
    .Y(_0220_),
    .A2(net87));
 sg13g2_nand3_1 _3047_ (.B(_1565_),
    .C(_1567_),
    .A(net166),
    .Y(_0221_));
 sg13g2_a21o_1 _3048_ (.A2(_0221_),
    .A1(net109),
    .B1(_1888_),
    .X(_0222_));
 sg13g2_o21ai_1 _3049_ (.B1(net158),
    .Y(_0223_),
    .A1(_0220_),
    .A2(_0222_));
 sg13g2_o21ai_1 _3050_ (.B1(_0223_),
    .Y(_0224_),
    .A1(_0214_),
    .A2(_0217_));
 sg13g2_nand2b_1 _3051_ (.Y(_0225_),
    .B(_0224_),
    .A_N(_0210_));
 sg13g2_nor2_1 _3052_ (.A(_1509_),
    .B(net53),
    .Y(_0226_));
 sg13g2_buf_2 _3053_ (.A(_0226_),
    .X(_0227_));
 sg13g2_nand2_1 _3054_ (.Y(_0228_),
    .A(net49),
    .B(_1853_));
 sg13g2_a221oi_1 _3055_ (.B2(_0228_),
    .C1(_1843_),
    .B1(_0227_),
    .A1(net136),
    .Y(_0229_),
    .A2(_1900_));
 sg13g2_o21ai_1 _3056_ (.B1(net76),
    .Y(_0230_),
    .A1(_1935_),
    .A2(_0229_));
 sg13g2_a221oi_1 _3057_ (.B2(net94),
    .C1(_0230_),
    .B1(_0225_),
    .A1(_0078_),
    .Y(_0231_),
    .A2(_0205_));
 sg13g2_nor3_2 _3058_ (.A(net167),
    .B(net151),
    .C(_1654_),
    .Y(_0232_));
 sg13g2_nor2_1 _3059_ (.A(_1390_),
    .B(net159),
    .Y(_0233_));
 sg13g2_a21oi_2 _3060_ (.B1(net53),
    .Y(_0234_),
    .A2(net78),
    .A1(net83));
 sg13g2_nor2_1 _3061_ (.A(_1803_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_nor2_1 _3062_ (.A(_1390_),
    .B(net110),
    .Y(_0236_));
 sg13g2_a221oi_1 _3063_ (.B2(_0235_),
    .C1(_0236_),
    .B1(_0233_),
    .A1(_1882_),
    .Y(_0237_),
    .A2(_0232_));
 sg13g2_a21oi_1 _3064_ (.A1(net151),
    .A2(net75),
    .Y(_0238_),
    .B1(_1723_));
 sg13g2_nand3_1 _3065_ (.B(net53),
    .C(_1581_),
    .A(net112),
    .Y(_0239_));
 sg13g2_buf_1 _3066_ (.A(_0239_),
    .X(_0240_));
 sg13g2_nand2_1 _3067_ (.Y(_0241_),
    .A(_1558_),
    .B(_0240_));
 sg13g2_nand3_1 _3068_ (.B(net85),
    .C(_1725_),
    .A(net84),
    .Y(_0242_));
 sg13g2_nand3_1 _3069_ (.B(net58),
    .C(_0140_),
    .A(net67),
    .Y(_0243_));
 sg13g2_nand4_1 _3070_ (.B(net95),
    .C(_0242_),
    .A(_1638_),
    .Y(_0244_),
    .D(_0243_));
 sg13g2_o21ai_1 _3071_ (.B1(_0244_),
    .Y(_0245_),
    .A1(_0238_),
    .A2(_0241_));
 sg13g2_o21ai_1 _3072_ (.B1(_1863_),
    .Y(_0246_),
    .A1(_1619_),
    .A2(_1621_));
 sg13g2_nand2_1 _3073_ (.Y(_0247_),
    .A(net80),
    .B(net15));
 sg13g2_a22oi_1 _3074_ (.Y(_0248_),
    .B1(_0247_),
    .B2(net13),
    .A2(_0246_),
    .A1(net33));
 sg13g2_buf_1 _3075_ (.A(net138),
    .X(_0249_));
 sg13g2_nand3_1 _3076_ (.B(_1513_),
    .C(net137),
    .A(net155),
    .Y(_0250_));
 sg13g2_nand3_1 _3077_ (.B(net54),
    .C(_0250_),
    .A(net55),
    .Y(_0251_));
 sg13g2_nand2_1 _3078_ (.Y(_0252_),
    .A(net115),
    .B(_0251_));
 sg13g2_nor4_1 _3079_ (.A(net156),
    .B(_1607_),
    .C(_0248_),
    .D(_0252_),
    .Y(_0253_));
 sg13g2_nor3_2 _3080_ (.A(net83),
    .B(_1506_),
    .C(_1675_),
    .Y(_0254_));
 sg13g2_a21oi_1 _3081_ (.A1(_1515_),
    .A2(net73),
    .Y(_0255_),
    .B1(_1543_));
 sg13g2_nor2_2 _3082_ (.A(net163),
    .B(net166),
    .Y(_0256_));
 sg13g2_o21ai_1 _3083_ (.B1(_0256_),
    .Y(_0257_),
    .A1(_0254_),
    .A2(_0255_));
 sg13g2_nor2_1 _3084_ (.A(_1591_),
    .B(net150),
    .Y(_0258_));
 sg13g2_a221oi_1 _3085_ (.B2(net57),
    .C1(net130),
    .B1(_0258_),
    .A1(net152),
    .Y(_0259_),
    .A2(_0254_));
 sg13g2_nor2_1 _3086_ (.A(_1660_),
    .B(net33),
    .Y(_0260_));
 sg13g2_nand2_1 _3087_ (.Y(_0261_),
    .A(net100),
    .B(net152));
 sg13g2_o21ai_1 _3088_ (.B1(_0227_),
    .Y(_0262_),
    .A1(net19),
    .A2(_0261_));
 sg13g2_a221oi_1 _3089_ (.B2(_0262_),
    .C1(net106),
    .B1(_0260_),
    .A1(_0257_),
    .Y(_0263_),
    .A2(_0259_));
 sg13g2_nor4_1 _3090_ (.A(_0237_),
    .B(_0245_),
    .C(_0253_),
    .D(_0263_),
    .Y(_0264_));
 sg13g2_o21ai_1 _3091_ (.B1(_1921_),
    .Y(_0265_),
    .A1(_0231_),
    .A2(_0264_));
 sg13g2_nor2_1 _3092_ (.A(net127),
    .B(_1899_),
    .Y(_0266_));
 sg13g2_nand2_1 _3093_ (.Y(_0267_),
    .A(net166),
    .B(net143));
 sg13g2_a21oi_1 _3094_ (.A1(_1899_),
    .A2(_0267_),
    .Y(_0268_),
    .B1(net59));
 sg13g2_o21ai_1 _3095_ (.B1(net89),
    .Y(_0269_),
    .A1(_0266_),
    .A2(_0268_));
 sg13g2_nor2_1 _3096_ (.A(_1583_),
    .B(_1800_),
    .Y(_0270_));
 sg13g2_nor2_2 _3097_ (.A(_1415_),
    .B(_1768_),
    .Y(_0271_));
 sg13g2_o21ai_1 _3098_ (.B1(_0271_),
    .Y(_0272_),
    .A1(_1982_),
    .A2(_0270_));
 sg13g2_a21o_1 _3099_ (.A2(_0272_),
    .A1(_0269_),
    .B1(net51),
    .X(_0273_));
 sg13g2_nor2_1 _3100_ (.A(net59),
    .B(_1667_),
    .Y(_0274_));
 sg13g2_o21ai_1 _3101_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_1550_),
    .A2(_0169_));
 sg13g2_nor2_1 _3102_ (.A(_1509_),
    .B(_1675_),
    .Y(_0276_));
 sg13g2_buf_2 _3103_ (.A(_0276_),
    .X(_0277_));
 sg13g2_nor2_1 _3104_ (.A(_1684_),
    .B(_1800_),
    .Y(_0278_));
 sg13g2_o21ai_1 _3105_ (.B1(_1667_),
    .Y(_0279_),
    .A1(net103),
    .A2(_1684_));
 sg13g2_a221oi_1 _3106_ (.B2(net93),
    .C1(net141),
    .B1(_0279_),
    .A1(_0277_),
    .Y(_0280_),
    .A2(_0278_));
 sg13g2_and2_1 _3107_ (.A(_0275_),
    .B(_0280_),
    .X(_0281_));
 sg13g2_nor2_1 _3108_ (.A(net41),
    .B(net56),
    .Y(_0282_));
 sg13g2_nor3_1 _3109_ (.A(_0282_),
    .B(net24),
    .C(net42),
    .Y(_0283_));
 sg13g2_nor2_1 _3110_ (.A(net120),
    .B(net110),
    .Y(_0284_));
 sg13g2_o21ai_1 _3111_ (.B1(_0284_),
    .Y(_0285_),
    .A1(net121),
    .A2(_0283_));
 sg13g2_o21ai_1 _3112_ (.B1(net136),
    .Y(_0286_),
    .A1(net24),
    .A2(net42));
 sg13g2_and2_1 _3113_ (.A(_1899_),
    .B(_0256_),
    .X(_0287_));
 sg13g2_nor3_1 _3114_ (.A(_1626_),
    .B(net29),
    .C(_1675_),
    .Y(_0288_));
 sg13g2_o21ai_1 _3115_ (.B1(net38),
    .Y(_0289_),
    .A1(_0287_),
    .A2(_0288_));
 sg13g2_nand2_1 _3116_ (.Y(_0290_),
    .A(_1390_),
    .B(net109));
 sg13g2_a21oi_1 _3117_ (.A1(net150),
    .A2(_1843_),
    .Y(_0291_),
    .B1(_0290_));
 sg13g2_nand3_1 _3118_ (.B(_0289_),
    .C(_0291_),
    .A(_0286_),
    .Y(_0292_));
 sg13g2_a22oi_1 _3119_ (.Y(_0293_),
    .B1(_0285_),
    .B2(_0292_),
    .A2(_0281_),
    .A1(_0273_));
 sg13g2_nor2_1 _3120_ (.A(_1676_),
    .B(net90),
    .Y(_0294_));
 sg13g2_o21ai_1 _3121_ (.B1(_1689_),
    .Y(_0295_),
    .A1(net39),
    .A2(net136));
 sg13g2_o21ai_1 _3122_ (.B1(net29),
    .Y(_0296_),
    .A1(net79),
    .A2(net111));
 sg13g2_nand4_1 _3123_ (.B(_0100_),
    .C(_0251_),
    .A(net159),
    .Y(_0297_),
    .D(_0296_));
 sg13g2_nand3_1 _3124_ (.B(_0259_),
    .C(_0297_),
    .A(_0257_),
    .Y(_0298_));
 sg13g2_nor2_1 _3125_ (.A(_1524_),
    .B(_0227_),
    .Y(_0299_));
 sg13g2_a21oi_1 _3126_ (.A1(net80),
    .A2(_0299_),
    .Y(_0300_),
    .B1(_1856_));
 sg13g2_a221oi_1 _3127_ (.B2(_0300_),
    .C1(_0237_),
    .B1(_0298_),
    .A1(_0294_),
    .Y(_0301_),
    .A2(_0295_));
 sg13g2_or3_1 _3128_ (.A(net101),
    .B(_0293_),
    .C(_0301_),
    .X(_0302_));
 sg13g2_nand3_1 _3129_ (.B(net33),
    .C(net64),
    .A(net62),
    .Y(_0303_));
 sg13g2_nor3_1 _3130_ (.A(_1492_),
    .B(net53),
    .C(_1592_),
    .Y(_0304_));
 sg13g2_o21ai_1 _3131_ (.B1(net55),
    .Y(_0305_),
    .A1(_1800_),
    .A2(_1888_));
 sg13g2_nand2b_1 _3132_ (.Y(_0306_),
    .B(_0305_),
    .A_N(_0304_));
 sg13g2_nor2_1 _3133_ (.A(_1810_),
    .B(_0306_),
    .Y(_0307_));
 sg13g2_nand3_1 _3134_ (.B(_1515_),
    .C(_1617_),
    .A(net57),
    .Y(_0308_));
 sg13g2_buf_1 _3135_ (.A(_0308_),
    .X(_0309_));
 sg13g2_a21oi_1 _3136_ (.A1(net104),
    .A2(_0169_),
    .Y(_0310_),
    .B1(_0309_));
 sg13g2_a21oi_1 _3137_ (.A1(net51),
    .A2(_0260_),
    .Y(_0311_),
    .B1(_0310_));
 sg13g2_o21ai_1 _3138_ (.B1(_0227_),
    .Y(_0312_),
    .A1(net43),
    .A2(_0206_));
 sg13g2_and2_1 _3139_ (.A(_1820_),
    .B(_0312_),
    .X(_0313_));
 sg13g2_a221oi_1 _3140_ (.B2(_0313_),
    .C1(net118),
    .B1(_0311_),
    .A1(_0303_),
    .Y(_0314_),
    .A2(_0307_));
 sg13g2_a21oi_1 _3141_ (.A1(net54),
    .A2(_1860_),
    .Y(_0315_),
    .B1(_1675_));
 sg13g2_a21oi_1 _3142_ (.A1(net84),
    .A2(_1617_),
    .Y(_0316_),
    .B1(net78));
 sg13g2_nand3_1 _3143_ (.B(_1590_),
    .C(_1863_),
    .A(_1586_),
    .Y(_0317_));
 sg13g2_o21ai_1 _3144_ (.B1(_1948_),
    .Y(_0318_),
    .A1(net65),
    .A2(_0317_));
 sg13g2_a221oi_1 _3145_ (.B2(net117),
    .C1(_0318_),
    .B1(_0316_),
    .A1(_1815_),
    .Y(_0319_),
    .A2(_0315_));
 sg13g2_nand2_1 _3146_ (.Y(_0320_),
    .A(_1493_),
    .B(net29));
 sg13g2_a221oi_1 _3147_ (.B2(_0315_),
    .C1(_1948_),
    .B1(_0320_),
    .A1(net27),
    .Y(_0321_),
    .A2(net62));
 sg13g2_nor4_1 _3148_ (.A(net102),
    .B(_1796_),
    .C(_0319_),
    .D(_0321_),
    .Y(_0322_));
 sg13g2_a21oi_2 _3149_ (.B1(_1560_),
    .Y(_0323_),
    .A2(net103),
    .A1(_1614_));
 sg13g2_o21ai_1 _3150_ (.B1(_1864_),
    .Y(_0324_),
    .A1(_1936_),
    .A2(_0323_));
 sg13g2_buf_1 _3151_ (.A(net84),
    .X(_0325_));
 sg13g2_o21ai_1 _3152_ (.B1(net30),
    .Y(_0326_),
    .A1(_0325_),
    .A2(net136));
 sg13g2_a21oi_1 _3153_ (.A1(net62),
    .A2(_0326_),
    .Y(_0327_),
    .B1(net102));
 sg13g2_a21oi_1 _3154_ (.A1(_1815_),
    .A2(_0315_),
    .Y(_0328_),
    .B1(net90));
 sg13g2_a221oi_1 _3155_ (.B2(_0327_),
    .C1(_0328_),
    .B1(_0324_),
    .A1(net121),
    .Y(_0329_),
    .A2(net63));
 sg13g2_nor2_1 _3156_ (.A(net82),
    .B(_0121_),
    .Y(_0330_));
 sg13g2_nand2_1 _3157_ (.Y(_0331_),
    .A(net105),
    .B(net72));
 sg13g2_a21o_1 _3158_ (.A2(_0331_),
    .A1(_0330_),
    .B1(_0170_),
    .X(_0332_));
 sg13g2_nor2_1 _3159_ (.A(net122),
    .B(_0316_),
    .Y(_0333_));
 sg13g2_nand2_1 _3160_ (.Y(_0334_),
    .A(net120),
    .B(_1760_));
 sg13g2_a21oi_1 _3161_ (.A1(_0332_),
    .A2(_0333_),
    .Y(_0335_),
    .B1(_0334_));
 sg13g2_a22oi_1 _3162_ (.Y(_0336_),
    .B1(_0329_),
    .B2(_0335_),
    .A2(_0322_),
    .A1(net169));
 sg13g2_o21ai_1 _3163_ (.B1(_0336_),
    .Y(_0337_),
    .A1(net168),
    .A2(_0314_));
 sg13g2_o21ai_1 _3164_ (.B1(_1981_),
    .Y(_0338_),
    .A1(_1562_),
    .A2(_1671_));
 sg13g2_nand2_1 _3165_ (.Y(_0339_),
    .A(net13),
    .B(_0338_));
 sg13g2_nand4_1 _3166_ (.B(_0100_),
    .C(_0309_),
    .A(_1707_),
    .Y(_0340_),
    .D(_0339_));
 sg13g2_a21oi_1 _3167_ (.A1(net72),
    .A2(_1978_),
    .Y(_0341_),
    .B1(_1791_));
 sg13g2_a21oi_1 _3168_ (.A1(_0330_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(_1707_));
 sg13g2_a21oi_1 _3169_ (.A1(_0105_),
    .A2(_0342_),
    .Y(_0343_),
    .B1(_1957_));
 sg13g2_a22oi_1 _3170_ (.Y(_0344_),
    .B1(_0340_),
    .B2(_0343_),
    .A2(_0306_),
    .A1(_0284_));
 sg13g2_nand2_1 _3171_ (.Y(_0345_),
    .A(_1746_),
    .B(net168));
 sg13g2_and4_1 _3172_ (.A(net142),
    .B(net108),
    .C(net96),
    .D(net148),
    .X(_0346_));
 sg13g2_a22oi_1 _3173_ (.Y(_0347_),
    .B1(_0346_),
    .B2(net50),
    .A2(net148),
    .A1(net45));
 sg13g2_nor2b_1 _3174_ (.A(_0127_),
    .B_N(_1456_),
    .Y(_0348_));
 sg13g2_and2_1 _3175_ (.A(_0347_),
    .B(_0348_),
    .X(_0349_));
 sg13g2_nor2_1 _3176_ (.A(net106),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_nor2_1 _3177_ (.A(net76),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nor3_2 _3178_ (.A(net157),
    .B(_1619_),
    .C(_1621_),
    .Y(_0352_));
 sg13g2_o21ai_1 _3179_ (.B1(net36),
    .Y(_0353_),
    .A1(net75),
    .A2(_0352_));
 sg13g2_nand2_1 _3180_ (.Y(_0354_),
    .A(_0277_),
    .B(_0353_));
 sg13g2_nand3_1 _3181_ (.B(_0151_),
    .C(_0354_),
    .A(net98),
    .Y(_0355_));
 sg13g2_o21ai_1 _3182_ (.B1(_1981_),
    .Y(_0356_),
    .A1(_1982_),
    .A2(_0323_));
 sg13g2_nand2_1 _3183_ (.Y(_0357_),
    .A(_0111_),
    .B(_0356_));
 sg13g2_nor2_1 _3184_ (.A(net167),
    .B(net96),
    .Y(_0358_));
 sg13g2_a221oi_1 _3185_ (.B2(_0358_),
    .C1(net80),
    .B1(net12),
    .A1(net142),
    .Y(_0359_),
    .A2(net108));
 sg13g2_nand2b_1 _3186_ (.Y(_0360_),
    .B(_0359_),
    .A_N(_0323_));
 sg13g2_a21oi_1 _3187_ (.A1(net17),
    .A2(_1686_),
    .Y(_0361_),
    .B1(net80));
 sg13g2_nor3_1 _3188_ (.A(net115),
    .B(_0345_),
    .C(_0361_),
    .Y(_0362_));
 sg13g2_nand4_1 _3189_ (.B(_0357_),
    .C(_0360_),
    .A(_0355_),
    .Y(_0363_),
    .D(_0362_));
 sg13g2_o21ai_1 _3190_ (.B1(_0363_),
    .Y(_0364_),
    .A1(_0345_),
    .A2(_0351_));
 sg13g2_nand2_1 _3191_ (.Y(_0365_),
    .A(net69),
    .B(_0186_));
 sg13g2_a221oi_1 _3192_ (.B2(_0364_),
    .C1(_0365_),
    .B1(_0344_),
    .A1(_0302_),
    .Y(_0366_),
    .A2(_0337_));
 sg13g2_nor3_1 _3193_ (.A(_1676_),
    .B(_1696_),
    .C(_1672_),
    .Y(_0367_));
 sg13g2_o21ai_1 _3194_ (.B1(_1875_),
    .Y(_0368_),
    .A1(_1803_),
    .A2(_0234_));
 sg13g2_nand3_1 _3195_ (.B(net41),
    .C(_0246_),
    .A(net37),
    .Y(_0369_));
 sg13g2_nand3_1 _3196_ (.B(net98),
    .C(_0369_),
    .A(_0240_),
    .Y(_0370_));
 sg13g2_nand3_1 _3197_ (.B(_0368_),
    .C(_0370_),
    .A(_1658_),
    .Y(_0371_));
 sg13g2_or3_1 _3198_ (.A(_1810_),
    .B(_0367_),
    .C(_0371_),
    .X(_0372_));
 sg13g2_o21ai_1 _3199_ (.B1(net127),
    .Y(_0373_),
    .A1(net57),
    .A2(_0087_));
 sg13g2_a21oi_1 _3200_ (.A1(net43),
    .A2(_1925_),
    .Y(_0374_),
    .B1(_1615_));
 sg13g2_a21oi_1 _3201_ (.A1(_1615_),
    .A2(_0099_),
    .Y(_0375_),
    .B1(_1935_));
 sg13g2_o21ai_1 _3202_ (.B1(_0375_),
    .Y(_0376_),
    .A1(net38),
    .A2(_0374_));
 sg13g2_nor2_1 _3203_ (.A(net55),
    .B(net71),
    .Y(_0377_));
 sg13g2_nor2_1 _3204_ (.A(net117),
    .B(_1964_),
    .Y(_0378_));
 sg13g2_o21ai_1 _3205_ (.B1(_0378_),
    .Y(_0379_),
    .A1(net35),
    .A2(_0377_));
 sg13g2_a22oi_1 _3206_ (.Y(_0380_),
    .B1(_0376_),
    .B2(_0379_),
    .A2(_0373_),
    .A1(net19));
 sg13g2_and2_1 _3207_ (.A(net83),
    .B(_1662_),
    .X(_0381_));
 sg13g2_buf_2 _3208_ (.A(_0381_),
    .X(_0382_));
 sg13g2_and2_1 _3209_ (.A(_1844_),
    .B(_0382_),
    .X(_0383_));
 sg13g2_nor3_1 _3210_ (.A(net35),
    .B(net23),
    .C(_0358_),
    .Y(_0384_));
 sg13g2_nor4_1 _3211_ (.A(net140),
    .B(net90),
    .C(_0383_),
    .D(_0384_),
    .Y(_0385_));
 sg13g2_a21oi_1 _3212_ (.A1(_1716_),
    .A2(net93),
    .Y(_0386_),
    .B1(net117));
 sg13g2_a21oi_1 _3213_ (.A1(_0105_),
    .A2(_0386_),
    .Y(_0387_),
    .B1(net107));
 sg13g2_a21oi_1 _3214_ (.A1(net159),
    .A2(_1483_),
    .Y(_0388_),
    .B1(net87));
 sg13g2_a21oi_1 _3215_ (.A1(_0325_),
    .A2(net75),
    .Y(_0389_),
    .B1(net149));
 sg13g2_o21ai_1 _3216_ (.B1(_0389_),
    .Y(_0390_),
    .A1(net23),
    .A2(_0388_));
 sg13g2_nand2_1 _3217_ (.Y(_0391_),
    .A(_1552_),
    .B(_0131_));
 sg13g2_buf_1 _3218_ (.A(net128),
    .X(_0392_));
 sg13g2_a221oi_1 _3219_ (.B2(net63),
    .C1(net86),
    .B1(_0391_),
    .A1(_0387_),
    .Y(_0393_),
    .A2(_0390_));
 sg13g2_or4_1 _3220_ (.A(net88),
    .B(_0380_),
    .C(_0385_),
    .D(_0393_),
    .X(_0394_));
 sg13g2_nand2_1 _3221_ (.Y(_0395_),
    .A(net40),
    .B(net134));
 sg13g2_a21oi_1 _3222_ (.A1(_1635_),
    .A2(_0395_),
    .Y(_0396_),
    .B1(_1508_));
 sg13g2_nor2_2 _3223_ (.A(net96),
    .B(net150),
    .Y(_0397_));
 sg13g2_o21ai_1 _3224_ (.B1(_1817_),
    .Y(_0398_),
    .A1(net47),
    .A2(_0397_));
 sg13g2_nand2_1 _3225_ (.Y(_0399_),
    .A(_0277_),
    .B(_0398_));
 sg13g2_o21ai_1 _3226_ (.B1(_0399_),
    .Y(_0400_),
    .A1(_1821_),
    .A2(_0396_));
 sg13g2_o21ai_1 _3227_ (.B1(_1820_),
    .Y(_0401_),
    .A1(net80),
    .A2(_0299_));
 sg13g2_a21o_1 _3228_ (.A2(_0400_),
    .A1(_1630_),
    .B1(_0401_),
    .X(_0402_));
 sg13g2_xnor2_1 _3229_ (.Y(_0403_),
    .A(_1574_),
    .B(_0185_));
 sg13g2_nand3_1 _3230_ (.B(_1740_),
    .C(_1744_),
    .A(_1737_),
    .Y(_0404_));
 sg13g2_nor2_1 _3231_ (.A(_1742_),
    .B(_1754_),
    .Y(_0405_));
 sg13g2_a21oi_1 _3232_ (.A1(_1754_),
    .A2(_0404_),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_nor2_1 _3233_ (.A(_0403_),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_nand4_1 _3234_ (.B(_0394_),
    .C(_0402_),
    .A(_0372_),
    .Y(_0408_),
    .D(_0407_));
 sg13g2_nor2_1 _3235_ (.A(net46),
    .B(net148),
    .Y(_0409_));
 sg13g2_a21oi_1 _3236_ (.A1(_0219_),
    .A2(_1908_),
    .Y(_0410_),
    .B1(net36));
 sg13g2_o21ai_1 _3237_ (.B1(_0410_),
    .Y(_0411_),
    .A1(net119),
    .A2(_1843_));
 sg13g2_o21ai_1 _3238_ (.B1(_1720_),
    .Y(_0412_),
    .A1(_0377_),
    .A2(_1843_));
 sg13g2_nand2_1 _3239_ (.Y(_0413_),
    .A(_1550_),
    .B(_0206_));
 sg13g2_nand3_1 _3240_ (.B(_1832_),
    .C(_0413_),
    .A(net169),
    .Y(_0414_));
 sg13g2_a221oi_1 _3241_ (.B2(_0412_),
    .C1(_0414_),
    .B1(_0411_),
    .A1(_0127_),
    .Y(_0415_),
    .A2(_0409_));
 sg13g2_o21ai_1 _3242_ (.B1(_0186_),
    .Y(_0416_),
    .A1(net118),
    .A2(net168));
 sg13g2_nor3_1 _3243_ (.A(net69),
    .B(_0415_),
    .C(_0416_),
    .Y(_0417_));
 sg13g2_nand2_1 _3244_ (.Y(_0418_),
    .A(net74),
    .B(_1978_));
 sg13g2_o21ai_1 _3245_ (.B1(_1507_),
    .Y(_0419_),
    .A1(net57),
    .A2(net71));
 sg13g2_o21ai_1 _3246_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_1938_),
    .A2(_0418_));
 sg13g2_nand4_1 _3247_ (.B(_0078_),
    .C(_0133_),
    .A(_1686_),
    .Y(_0421_),
    .D(_0420_));
 sg13g2_nor2_1 _3248_ (.A(net120),
    .B(net168),
    .Y(_0422_));
 sg13g2_a21oi_1 _3249_ (.A1(net139),
    .A2(net99),
    .Y(_0423_),
    .B1(net131));
 sg13g2_xnor2_1 _3250_ (.Y(_0424_),
    .A(net52),
    .B(_0423_));
 sg13g2_nand2_1 _3251_ (.Y(_0425_),
    .A(net141),
    .B(net98));
 sg13g2_a21o_1 _3252_ (.A2(_0424_),
    .A1(net27),
    .B1(_0425_),
    .X(_0426_));
 sg13g2_nand2_1 _3253_ (.Y(_0427_),
    .A(net48),
    .B(_1646_));
 sg13g2_nor2_1 _3254_ (.A(net130),
    .B(net145),
    .Y(_0428_));
 sg13g2_and4_1 _3255_ (.A(_1528_),
    .B(_1530_),
    .C(_1649_),
    .D(_1650_),
    .X(_0429_));
 sg13g2_buf_2 _3256_ (.A(_0429_),
    .X(_0430_));
 sg13g2_nor3_1 _3257_ (.A(net129),
    .B(net153),
    .C(_0430_),
    .Y(_0431_));
 sg13g2_o21ai_1 _3258_ (.B1(net26),
    .Y(_0432_),
    .A1(_0428_),
    .A2(_0431_));
 sg13g2_o21ai_1 _3259_ (.B1(net41),
    .Y(_0433_),
    .A1(net59),
    .A2(net100));
 sg13g2_nor2_1 _3260_ (.A(net141),
    .B(_1550_),
    .Y(_0434_));
 sg13g2_nand4_1 _3261_ (.B(_0432_),
    .C(_0433_),
    .A(_0427_),
    .Y(_0435_),
    .D(_0434_));
 sg13g2_o21ai_1 _3262_ (.B1(net32),
    .Y(_0436_),
    .A1(_0121_),
    .A2(net45));
 sg13g2_or2_1 _3263_ (.X(_0437_),
    .B(_0246_),
    .A(net50));
 sg13g2_nor2_1 _3264_ (.A(net124),
    .B(_1953_),
    .Y(_0438_));
 sg13g2_nand4_1 _3265_ (.B(_0436_),
    .C(_0437_),
    .A(net128),
    .Y(_0439_),
    .D(_0438_));
 sg13g2_and4_1 _3266_ (.A(_0422_),
    .B(_0426_),
    .C(_0435_),
    .D(_0439_),
    .X(_0440_));
 sg13g2_nand2_1 _3267_ (.Y(_0441_),
    .A(_1892_),
    .B(_1695_));
 sg13g2_a21oi_1 _3268_ (.A1(net135),
    .A2(_1695_),
    .Y(_0442_),
    .B1(_0430_));
 sg13g2_a22oi_1 _3269_ (.Y(_0443_),
    .B1(_0442_),
    .B2(net16),
    .A2(_0441_),
    .A1(_0202_));
 sg13g2_a22oi_1 _3270_ (.Y(_0444_),
    .B1(_0443_),
    .B2(net119),
    .A2(_0424_),
    .A1(net27));
 sg13g2_nand2_1 _3271_ (.Y(_0445_),
    .A(net100),
    .B(_1652_));
 sg13g2_a21oi_2 _3272_ (.B1(_0202_),
    .Y(_0446_),
    .A2(_1652_),
    .A1(net57));
 sg13g2_nor2_1 _3273_ (.A(_0149_),
    .B(_0423_),
    .Y(_0447_));
 sg13g2_a221oi_1 _3274_ (.B2(net49),
    .C1(net125),
    .B1(_0447_),
    .A1(_0445_),
    .Y(_0448_),
    .A2(_0446_));
 sg13g2_nor4_1 _3275_ (.A(net106),
    .B(_0444_),
    .C(_0334_),
    .D(_0448_),
    .Y(_0449_));
 sg13g2_a21oi_1 _3276_ (.A1(_0421_),
    .A2(_0440_),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_a22oi_1 _3277_ (.Y(_0451_),
    .B1(_0417_),
    .B2(_0450_),
    .A2(_0186_),
    .A1(_0183_));
 sg13g2_nor2_1 _3278_ (.A(net41),
    .B(_0397_),
    .Y(_0452_));
 sg13g2_a21oi_1 _3279_ (.A1(net26),
    .A2(net93),
    .Y(_0453_),
    .B1(net126));
 sg13g2_o21ai_1 _3280_ (.B1(_0453_),
    .Y(_0454_),
    .A1(net23),
    .A2(_0452_));
 sg13g2_nand2_1 _3281_ (.Y(_0455_),
    .A(net151),
    .B(_1782_));
 sg13g2_a22oi_1 _3282_ (.Y(_0456_),
    .B1(net87),
    .B2(_0455_),
    .A2(net41),
    .A1(net151));
 sg13g2_a21oi_1 _3283_ (.A1(net50),
    .A2(net111),
    .Y(_0457_),
    .B1(net144));
 sg13g2_o21ai_1 _3284_ (.B1(_0457_),
    .Y(_0458_),
    .A1(net23),
    .A2(_0456_));
 sg13g2_nand2_1 _3285_ (.Y(_0459_),
    .A(net37),
    .B(_1646_));
 sg13g2_nand3_1 _3286_ (.B(net40),
    .C(_1863_),
    .A(net37),
    .Y(_0460_));
 sg13g2_nand4_1 _3287_ (.B(_0459_),
    .C(_0105_),
    .A(net95),
    .Y(_0461_),
    .D(_0460_));
 sg13g2_nand3_1 _3288_ (.B(_0458_),
    .C(_0461_),
    .A(_0454_),
    .Y(_0462_));
 sg13g2_nand2b_1 _3289_ (.Y(_0463_),
    .B(net37),
    .A_N(net137));
 sg13g2_a21oi_1 _3290_ (.A1(_1543_),
    .A2(net137),
    .Y(_0464_),
    .B1(net68));
 sg13g2_a21o_1 _3291_ (.A2(_0464_),
    .A1(_0463_),
    .B1(net36),
    .X(_0465_));
 sg13g2_nand2_1 _3292_ (.Y(_0466_),
    .A(net67),
    .B(_1800_));
 sg13g2_nor2_2 _3293_ (.A(_1691_),
    .B(_1532_),
    .Y(_0467_));
 sg13g2_a22oi_1 _3294_ (.Y(_0468_),
    .B1(_0467_),
    .B2(_1623_),
    .A2(_1953_),
    .A1(net57));
 sg13g2_and3_1 _3295_ (.X(_0469_),
    .A(net158),
    .B(_0466_),
    .C(_0468_));
 sg13g2_a221oi_1 _3296_ (.B2(_0469_),
    .C1(net90),
    .B1(_0465_),
    .A1(net136),
    .Y(_0470_),
    .A2(_0391_));
 sg13g2_a21oi_1 _3297_ (.A1(net31),
    .A2(net20),
    .Y(_0471_),
    .B1(_0382_));
 sg13g2_nand2b_1 _3298_ (.Y(_0472_),
    .B(_0256_),
    .A_N(_0471_));
 sg13g2_o21ai_1 _3299_ (.B1(net29),
    .Y(_0473_),
    .A1(net52),
    .A2(_1844_));
 sg13g2_o21ai_1 _3300_ (.B1(net79),
    .Y(_0474_),
    .A1(net58),
    .A2(_1592_));
 sg13g2_a22oi_1 _3301_ (.Y(_0475_),
    .B1(_0473_),
    .B2(_0474_),
    .A2(_0373_),
    .A1(net21));
 sg13g2_a21o_1 _3302_ (.A2(_0475_),
    .A1(net110),
    .B1(net114),
    .X(_0476_));
 sg13g2_a221oi_1 _3303_ (.B2(_0472_),
    .C1(_0476_),
    .B1(_0470_),
    .A1(net94),
    .Y(_0477_),
    .A2(_0462_));
 sg13g2_o21ai_1 _3304_ (.B1(_1562_),
    .Y(_0478_),
    .A1(net39),
    .A2(net136));
 sg13g2_o21ai_1 _3305_ (.B1(_0399_),
    .Y(_0479_),
    .A1(_0396_),
    .A2(_0478_));
 sg13g2_a221oi_1 _3306_ (.B2(net149),
    .C1(net16),
    .B1(_1675_),
    .A1(_1788_),
    .Y(_0480_),
    .A2(net99));
 sg13g2_o21ai_1 _3307_ (.B1(_0078_),
    .Y(_0481_),
    .A1(net33),
    .A2(_0480_));
 sg13g2_nand3_1 _3308_ (.B(net22),
    .C(_0250_),
    .A(net48),
    .Y(_0482_));
 sg13g2_nand4_1 _3309_ (.B(net89),
    .C(_0242_),
    .A(net121),
    .Y(_0483_),
    .D(_0482_));
 sg13g2_nand3_1 _3310_ (.B(_0481_),
    .C(_0483_),
    .A(net88),
    .Y(_0484_));
 sg13g2_a221oi_1 _3311_ (.B2(net81),
    .C1(_0484_),
    .B1(_0479_),
    .A1(_1914_),
    .Y(_0485_),
    .A2(_0371_));
 sg13g2_or3_1 _3312_ (.A(_1945_),
    .B(_0477_),
    .C(_0485_),
    .X(_0486_));
 sg13g2_o21ai_1 _3313_ (.B1(net116),
    .Y(_0487_),
    .A1(net24),
    .A2(_1665_));
 sg13g2_o21ai_1 _3314_ (.B1(_0084_),
    .Y(_0488_),
    .A1(net82),
    .A2(net52));
 sg13g2_o21ai_1 _3315_ (.B1(net141),
    .Y(_0489_),
    .A1(net65),
    .A2(_0118_));
 sg13g2_a221oi_1 _3316_ (.B2(net74),
    .C1(_0489_),
    .B1(_0488_),
    .A1(_0445_),
    .Y(_0490_),
    .A2(_0446_));
 sg13g2_a21oi_1 _3317_ (.A1(_0487_),
    .A2(_0490_),
    .Y(_0491_),
    .B1(net114));
 sg13g2_nand3_1 _3318_ (.B(net139),
    .C(net99),
    .A(net157),
    .Y(_0492_));
 sg13g2_buf_1 _3319_ (.A(_0492_),
    .X(_0493_));
 sg13g2_a21oi_1 _3320_ (.A1(net87),
    .A2(_0493_),
    .Y(_0494_),
    .B1(net21));
 sg13g2_nor2_1 _3321_ (.A(net38),
    .B(net119),
    .Y(_0495_));
 sg13g2_o21ai_1 _3322_ (.B1(_0495_),
    .Y(_0496_),
    .A1(net45),
    .A2(_0494_));
 sg13g2_a221oi_1 _3323_ (.B2(_0430_),
    .C1(net65),
    .B1(_1899_),
    .A1(net68),
    .Y(_0497_),
    .A2(_1617_));
 sg13g2_or3_1 _3324_ (.A(net64),
    .B(_0497_),
    .C(_0270_),
    .X(_0498_));
 sg13g2_nand3_1 _3325_ (.B(_0496_),
    .C(_0498_),
    .A(net94),
    .Y(_0499_));
 sg13g2_a21oi_1 _3326_ (.A1(_1828_),
    .A2(_0419_),
    .Y(_0500_),
    .B1(_1872_));
 sg13g2_a21oi_1 _3327_ (.A1(_0436_),
    .A2(_0500_),
    .Y(_0501_),
    .B1(net120));
 sg13g2_nand2_1 _3328_ (.Y(_0502_),
    .A(net59),
    .B(net127));
 sg13g2_a221oi_1 _3329_ (.B2(net61),
    .C1(net47),
    .B1(_0169_),
    .A1(_0430_),
    .Y(_0503_),
    .A2(_1667_));
 sg13g2_a22oi_1 _3330_ (.Y(_0504_),
    .B1(_0433_),
    .B2(_0503_),
    .A2(net72),
    .A1(_0502_));
 sg13g2_or2_1 _3331_ (.X(_0505_),
    .B(_0504_),
    .A(net86));
 sg13g2_a221oi_1 _3332_ (.B2(_0505_),
    .C1(net70),
    .B1(_0501_),
    .A1(_0491_),
    .Y(_0506_),
    .A2(_0499_));
 sg13g2_nor3_1 _3333_ (.A(net169),
    .B(_0183_),
    .C(_0506_),
    .Y(_0507_));
 sg13g2_a22oi_1 _3334_ (.Y(_0509_),
    .B1(_0486_),
    .B2(_0507_),
    .A2(_0451_),
    .A1(_0408_));
 sg13g2_a21o_1 _3335_ (.A2(_0366_),
    .A1(_0265_),
    .B1(_0509_),
    .X(_0510_));
 sg13g2_inv_1 _3336_ (.Y(_0511_),
    .A(_0183_));
 sg13g2_nor3_1 _3337_ (.A(net37),
    .B(net62),
    .C(net42),
    .Y(_0512_));
 sg13g2_a21oi_1 _3338_ (.A1(net27),
    .A2(net44),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_o21ai_1 _3339_ (.B1(_1626_),
    .Y(_0514_),
    .A1(net151),
    .A2(net34));
 sg13g2_nand2_1 _3340_ (.Y(_0515_),
    .A(net163),
    .B(net55));
 sg13g2_a21oi_1 _3341_ (.A1(net162),
    .A2(net100),
    .Y(_0516_),
    .B1(net68));
 sg13g2_a221oi_1 _3342_ (.B2(_1689_),
    .C1(_1607_),
    .B1(_0516_),
    .A1(net22),
    .Y(_0517_),
    .A2(_0515_));
 sg13g2_a21oi_1 _3343_ (.A1(net162),
    .A2(_0430_),
    .Y(_0518_),
    .B1(net62));
 sg13g2_nand2b_1 _3344_ (.Y(_0520_),
    .B(net22),
    .A_N(_0256_));
 sg13g2_o21ai_1 _3345_ (.B1(net102),
    .Y(_0521_),
    .A1(_0518_),
    .A2(_0520_));
 sg13g2_a221oi_1 _3346_ (.B2(_0517_),
    .C1(_0521_),
    .B1(_0514_),
    .A1(_0256_),
    .Y(_0522_),
    .A2(_0513_));
 sg13g2_o21ai_1 _3347_ (.B1(_1968_),
    .Y(_0523_),
    .A1(net50),
    .A2(net62));
 sg13g2_o21ai_1 _3348_ (.B1(net107),
    .Y(_0524_),
    .A1(net140),
    .A2(_0523_));
 sg13g2_o21ai_1 _3349_ (.B1(_1938_),
    .Y(_0525_),
    .A1(_0190_),
    .A2(_0493_));
 sg13g2_nor2_1 _3350_ (.A(net128),
    .B(net162),
    .Y(_0526_));
 sg13g2_a22oi_1 _3351_ (.Y(_0527_),
    .B1(_0430_),
    .B2(_0352_),
    .A2(net56),
    .A1(net61));
 sg13g2_nor4_1 _3352_ (.A(net128),
    .B(net158),
    .C(net12),
    .D(_0527_),
    .Y(_0528_));
 sg13g2_a221oi_1 _3353_ (.B2(_0526_),
    .C1(_0528_),
    .B1(_0525_),
    .A1(net121),
    .Y(_0529_),
    .A2(_0524_));
 sg13g2_a221oi_1 _3354_ (.B2(net159),
    .C1(net48),
    .B1(net75),
    .A1(_1788_),
    .Y(_0531_),
    .A2(_1789_));
 sg13g2_o21ai_1 _3355_ (.B1(net141),
    .Y(_0532_),
    .A1(_1456_),
    .A2(net28));
 sg13g2_o21ai_1 _3356_ (.B1(_1935_),
    .Y(_0533_),
    .A1(_0531_),
    .A2(_0532_));
 sg13g2_nor2_1 _3357_ (.A(net151),
    .B(net125),
    .Y(_0534_));
 sg13g2_mux2_1 _3358_ (.A0(_1550_),
    .A1(_1646_),
    .S(net79),
    .X(_0535_));
 sg13g2_a21oi_1 _3359_ (.A1(net40),
    .A2(_0267_),
    .Y(_0536_),
    .B1(net61));
 sg13g2_nor2_1 _3360_ (.A(net22),
    .B(net124),
    .Y(_0537_));
 sg13g2_nor4_1 _3361_ (.A(_1456_),
    .B(net30),
    .C(_1610_),
    .D(net124),
    .Y(_0538_));
 sg13g2_a221oi_1 _3362_ (.B2(_0537_),
    .C1(_0538_),
    .B1(_0536_),
    .A1(_0534_),
    .Y(_0539_),
    .A2(_0535_));
 sg13g2_a21oi_1 _3363_ (.A1(_0533_),
    .A2(_0539_),
    .Y(_0540_),
    .B1(net88));
 sg13g2_o21ai_1 _3364_ (.B1(_0540_),
    .Y(_0542_),
    .A1(_0522_),
    .A2(_0529_));
 sg13g2_nand3_1 _3365_ (.B(net40),
    .C(_0467_),
    .A(net65),
    .Y(_0543_));
 sg13g2_o21ai_1 _3366_ (.B1(_0543_),
    .Y(_0544_),
    .A1(_1552_),
    .A2(_0467_));
 sg13g2_or4_1 _3367_ (.A(net121),
    .B(net116),
    .C(net93),
    .D(_0544_),
    .X(_0545_));
 sg13g2_a21oi_1 _3368_ (.A1(net26),
    .A2(net127),
    .Y(_0546_),
    .B1(_0352_));
 sg13g2_nor2_1 _3369_ (.A(net119),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_nor2_1 _3370_ (.A(_1669_),
    .B(net123),
    .Y(_0548_));
 sg13g2_o21ai_1 _3371_ (.B1(_0216_),
    .Y(_0549_),
    .A1(net21),
    .A2(_0548_));
 sg13g2_o21ai_1 _3372_ (.B1(net115),
    .Y(_0550_),
    .A1(_0547_),
    .A2(_0549_));
 sg13g2_nor3_1 _3373_ (.A(net65),
    .B(net71),
    .C(_1667_),
    .Y(_0551_));
 sg13g2_o21ai_1 _3374_ (.B1(net31),
    .Y(_0553_),
    .A1(net34),
    .A2(_0551_));
 sg13g2_nand3_1 _3375_ (.B(_1534_),
    .C(net127),
    .A(net12),
    .Y(_0554_));
 sg13g2_nand4_1 _3376_ (.B(net116),
    .C(_0553_),
    .A(net86),
    .Y(_0555_),
    .D(_0554_));
 sg13g2_nand4_1 _3377_ (.B(_0545_),
    .C(_0550_),
    .A(net76),
    .Y(_0556_),
    .D(_0555_));
 sg13g2_nand3_1 _3378_ (.B(_0542_),
    .C(_0556_),
    .A(_1921_),
    .Y(_0557_));
 sg13g2_nor4_1 _3379_ (.A(net120),
    .B(_1599_),
    .C(_1936_),
    .D(_0304_),
    .Y(_0558_));
 sg13g2_nor2_1 _3380_ (.A(net67),
    .B(_1534_),
    .Y(_0559_));
 sg13g2_o21ai_1 _3381_ (.B1(net35),
    .Y(_0560_),
    .A1(_1908_),
    .A2(_0559_));
 sg13g2_nor2_1 _3382_ (.A(_0190_),
    .B(net90),
    .Y(_0561_));
 sg13g2_a21oi_1 _3383_ (.A1(net37),
    .A2(_0127_),
    .Y(_0562_),
    .B1(_1695_));
 sg13g2_nand2b_1 _3384_ (.Y(_0564_),
    .B(net125),
    .A_N(_0562_));
 sg13g2_a221oi_1 _3385_ (.B2(_0324_),
    .C1(_0177_),
    .B1(_0564_),
    .A1(_0560_),
    .Y(_0565_),
    .A2(_0561_));
 sg13g2_a21oi_1 _3386_ (.A1(_1690_),
    .A2(_1617_),
    .Y(_0566_),
    .B1(net37));
 sg13g2_nor3_1 _3387_ (.A(net51),
    .B(_0382_),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_nor2b_1 _3388_ (.A(_1957_),
    .B_N(_0567_),
    .Y(_0568_));
 sg13g2_nor4_1 _3389_ (.A(_0345_),
    .B(_0558_),
    .C(_0565_),
    .D(_0568_),
    .Y(_0569_));
 sg13g2_o21ai_1 _3390_ (.B1(_1869_),
    .Y(_0570_),
    .A1(net79),
    .A2(_0430_));
 sg13g2_a21oi_1 _3391_ (.A1(_0131_),
    .A2(_0570_),
    .Y(_0571_),
    .B1(net124));
 sg13g2_a21oi_1 _3392_ (.A1(_1475_),
    .A2(net103),
    .Y(_0572_),
    .B1(net142));
 sg13g2_a21oi_1 _3393_ (.A1(_0116_),
    .A2(net103),
    .Y(_0573_),
    .B1(net108));
 sg13g2_nand2_1 _3394_ (.Y(_0575_),
    .A(_1456_),
    .B(_1804_));
 sg13g2_nor4_1 _3395_ (.A(_0559_),
    .B(_0572_),
    .C(_0573_),
    .D(_0575_),
    .Y(_0576_));
 sg13g2_nor3_1 _3396_ (.A(net161),
    .B(net12),
    .C(_0575_),
    .Y(_0577_));
 sg13g2_nor4_1 _3397_ (.A(_1796_),
    .B(_0571_),
    .C(_0576_),
    .D(_0577_),
    .Y(_0578_));
 sg13g2_o21ai_1 _3398_ (.B1(_0578_),
    .Y(_0579_),
    .A1(net77),
    .A2(_0567_));
 sg13g2_a21oi_1 _3399_ (.A1(_0569_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(_1762_));
 sg13g2_nor2_1 _3400_ (.A(net152),
    .B(net149),
    .Y(_0581_));
 sg13g2_a22oi_1 _3401_ (.Y(_0582_),
    .B1(_0581_),
    .B2(_1869_),
    .A2(net149),
    .A1(net71));
 sg13g2_nor2_1 _3402_ (.A(net128),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_nand2_1 _3403_ (.Y(_0584_),
    .A(net154),
    .B(_1968_));
 sg13g2_nor2_1 _3404_ (.A(net27),
    .B(_0584_),
    .Y(_0586_));
 sg13g2_nand2_1 _3405_ (.Y(_0587_),
    .A(net75),
    .B(_0581_));
 sg13g2_o21ai_1 _3406_ (.B1(_0587_),
    .Y(_0588_),
    .A1(net47),
    .A2(net117));
 sg13g2_a221oi_1 _3407_ (.B2(_0588_),
    .C1(net63),
    .B1(_0586_),
    .A1(_1689_),
    .Y(_0589_),
    .A2(_0583_));
 sg13g2_o21ai_1 _3408_ (.B1(_1906_),
    .Y(_0590_),
    .A1(net56),
    .A2(net134));
 sg13g2_a221oi_1 _3409_ (.B2(net16),
    .C1(net138),
    .B1(_0590_),
    .A1(net28),
    .Y(_0591_),
    .A2(_0277_));
 sg13g2_nor2_1 _3410_ (.A(_0118_),
    .B(_0267_),
    .Y(_0592_));
 sg13g2_o21ai_1 _3411_ (.B1(net162),
    .Y(_0593_),
    .A1(_0227_),
    .A2(_0592_));
 sg13g2_a21oi_1 _3412_ (.A1(_0591_),
    .A2(_0593_),
    .Y(_0594_),
    .B1(net118));
 sg13g2_o21ai_1 _3413_ (.B1(_1813_),
    .Y(_0595_),
    .A1(_1593_),
    .A2(_0203_));
 sg13g2_nor3_1 _3414_ (.A(net18),
    .B(net87),
    .C(net149),
    .Y(_0597_));
 sg13g2_a21oi_1 _3415_ (.A1(_1593_),
    .A2(_0597_),
    .Y(_0598_),
    .B1(net120));
 sg13g2_nor2_1 _3416_ (.A(_1702_),
    .B(_0430_),
    .Y(_0599_));
 sg13g2_a22oi_1 _3417_ (.Y(_0600_),
    .B1(_1900_),
    .B2(_1774_),
    .A2(_0599_),
    .A1(net18));
 sg13g2_o21ai_1 _3418_ (.B1(net110),
    .Y(_0601_),
    .A1(_1659_),
    .A2(_0600_));
 sg13g2_a22oi_1 _3419_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net114),
    .A2(_0598_),
    .A1(_0595_));
 sg13g2_nand4_1 _3420_ (.B(net142),
    .C(net108),
    .A(net163),
    .Y(_0603_),
    .D(net123));
 sg13g2_nand4_1 _3421_ (.B(net142),
    .C(net108),
    .A(net167),
    .Y(_0604_),
    .D(net137));
 sg13g2_nand4_1 _3422_ (.B(net29),
    .C(_0603_),
    .A(net65),
    .Y(_0605_),
    .D(_0604_));
 sg13g2_nand3_1 _3423_ (.B(net41),
    .C(_1852_),
    .A(net32),
    .Y(_0606_));
 sg13g2_nand3_1 _3424_ (.B(_0605_),
    .C(_0606_),
    .A(net107),
    .Y(_0608_));
 sg13g2_nor3_1 _3425_ (.A(_0392_),
    .B(_1944_),
    .C(_0608_),
    .Y(_0609_));
 sg13g2_a221oi_1 _3426_ (.B2(net101),
    .C1(_0609_),
    .B1(_0602_),
    .A1(_0589_),
    .Y(_0610_),
    .A2(_0594_));
 sg13g2_nand2_1 _3427_ (.Y(_0611_),
    .A(_0466_),
    .B(_0468_));
 sg13g2_nor2_1 _3428_ (.A(net13),
    .B(_0464_),
    .Y(_0612_));
 sg13g2_o21ai_1 _3429_ (.B1(net95),
    .Y(_0613_),
    .A1(_0611_),
    .A2(_0612_));
 sg13g2_nand4_1 _3430_ (.B(net30),
    .C(net75),
    .A(net61),
    .Y(_0614_),
    .D(net98));
 sg13g2_o21ai_1 _3431_ (.B1(_0614_),
    .Y(_0615_),
    .A1(net95),
    .A2(_0118_));
 sg13g2_nor3_1 _3432_ (.A(net32),
    .B(net87),
    .C(net105),
    .Y(_0616_));
 sg13g2_a21oi_1 _3433_ (.A1(net103),
    .A2(net98),
    .Y(_0617_),
    .B1(net48));
 sg13g2_nor4_1 _3434_ (.A(net31),
    .B(_0441_),
    .C(_0616_),
    .D(_0617_),
    .Y(_0619_));
 sg13g2_nand2_1 _3435_ (.Y(_0620_),
    .A(net36),
    .B(net105));
 sg13g2_nand3_1 _3436_ (.B(net89),
    .C(_0087_),
    .A(net48),
    .Y(_0621_));
 sg13g2_o21ai_1 _3437_ (.B1(net105),
    .Y(_0622_),
    .A1(net26),
    .A2(net51));
 sg13g2_a22oi_1 _3438_ (.Y(_0623_),
    .B1(_0622_),
    .B2(_1786_),
    .A2(_0621_),
    .A1(_0620_));
 sg13g2_nor4_1 _3439_ (.A(_0177_),
    .B(_0615_),
    .C(_0619_),
    .D(_0623_),
    .Y(_0624_));
 sg13g2_and2_1 _3440_ (.A(_0459_),
    .B(_0105_),
    .X(_0625_));
 sg13g2_nand2_1 _3441_ (.Y(_0626_),
    .A(_0441_),
    .B(_0625_));
 sg13g2_nand4_1 _3442_ (.B(net139),
    .C(net99),
    .A(net157),
    .Y(_0627_),
    .D(net96));
 sg13g2_nand3_1 _3443_ (.B(net43),
    .C(_0627_),
    .A(net61),
    .Y(_0628_));
 sg13g2_a21o_1 _3444_ (.A2(_0628_),
    .A1(_0457_),
    .B1(net128),
    .X(_0630_));
 sg13g2_xnor2_1 _3445_ (.Y(_0631_),
    .A(net40),
    .B(_1610_));
 sg13g2_a221oi_1 _3446_ (.B2(_0631_),
    .C1(net125),
    .B1(_0227_),
    .A1(net12),
    .Y(_0632_),
    .A2(_1625_));
 sg13g2_nor3_1 _3447_ (.A(net88),
    .B(_0630_),
    .C(_0632_),
    .Y(_0633_));
 sg13g2_a22oi_1 _3448_ (.Y(_0634_),
    .B1(_0626_),
    .B2(_0633_),
    .A2(_0624_),
    .A1(_0613_));
 sg13g2_nand2b_1 _3449_ (.Y(_0635_),
    .B(_0634_),
    .A_N(_0610_));
 sg13g2_nand2_1 _3450_ (.Y(_0636_),
    .A(net138),
    .B(net130));
 sg13g2_nor4_1 _3451_ (.A(net36),
    .B(_1499_),
    .C(_0377_),
    .D(_0636_),
    .Y(_0637_));
 sg13g2_a21oi_1 _3452_ (.A1(_1940_),
    .A2(_0475_),
    .Y(_0638_),
    .B1(_0637_));
 sg13g2_nand2_1 _3453_ (.Y(_0639_),
    .A(_1534_),
    .B(_0202_));
 sg13g2_a221oi_1 _3454_ (.B2(_1717_),
    .C1(net104),
    .B1(_0639_),
    .A1(net136),
    .Y(_0641_),
    .A2(_0419_));
 sg13g2_a21oi_1 _3455_ (.A1(_1520_),
    .A2(_1763_),
    .Y(_0642_),
    .B1(net87));
 sg13g2_o21ai_1 _3456_ (.B1(net105),
    .Y(_0643_),
    .A1(net82),
    .A2(_1540_));
 sg13g2_a221oi_1 _3457_ (.B2(net135),
    .C1(net31),
    .B1(_0643_),
    .A1(_1815_),
    .Y(_0644_),
    .A2(_0642_));
 sg13g2_o21ai_1 _3458_ (.B1(_1820_),
    .Y(_0645_),
    .A1(_0641_),
    .A2(_0644_));
 sg13g2_o21ai_1 _3459_ (.B1(_0645_),
    .Y(_0646_),
    .A1(net92),
    .A2(_0638_));
 sg13g2_nor2_1 _3460_ (.A(net76),
    .B(_1747_),
    .Y(_0647_));
 sg13g2_xnor2_1 _3461_ (.Y(_0648_),
    .A(net138),
    .B(_1557_));
 sg13g2_a21o_1 _3462_ (.A2(_0648_),
    .A1(net44),
    .B1(net14),
    .X(_0649_));
 sg13g2_nand2_1 _3463_ (.Y(_0650_),
    .A(_1717_),
    .B(_1917_));
 sg13g2_nand2_1 _3464_ (.Y(_0652_),
    .A(net119),
    .B(net127));
 sg13g2_a221oi_1 _3465_ (.B2(net11),
    .C1(net115),
    .B1(_0652_),
    .A1(_1786_),
    .Y(_0653_),
    .A2(_0650_));
 sg13g2_a21oi_1 _3466_ (.A1(_0639_),
    .A2(_0649_),
    .Y(_0654_),
    .B1(_0653_));
 sg13g2_a221oi_1 _3467_ (.B2(_0654_),
    .C1(net69),
    .B1(_0647_),
    .A1(net91),
    .Y(_0655_),
    .A2(_0646_));
 sg13g2_a22oi_1 _3468_ (.Y(_0656_),
    .B1(_0635_),
    .B2(_0655_),
    .A2(_0580_),
    .A1(_0557_));
 sg13g2_nor2_1 _3469_ (.A(net166),
    .B(_1581_),
    .Y(_0657_));
 sg13g2_o21ai_1 _3470_ (.B1(_1723_),
    .Y(_0658_),
    .A1(_1866_),
    .A2(_0657_));
 sg13g2_nor2_1 _3471_ (.A(_1524_),
    .B(_0254_),
    .Y(_0659_));
 sg13g2_a221oi_1 _3472_ (.B2(net89),
    .C1(net128),
    .B1(_0659_),
    .A1(net98),
    .Y(_0660_),
    .A2(_0658_));
 sg13g2_nor2_1 _3473_ (.A(net67),
    .B(_1899_),
    .Y(_0661_));
 sg13g2_o21ai_1 _3474_ (.B1(net159),
    .Y(_0663_),
    .A1(_0661_),
    .A2(_0254_));
 sg13g2_nand3_1 _3475_ (.B(_0259_),
    .C(_0663_),
    .A(_0257_),
    .Y(_0664_));
 sg13g2_nor2_1 _3476_ (.A(_1623_),
    .B(_0467_),
    .Y(_0665_));
 sg13g2_nand3_1 _3477_ (.B(net93),
    .C(_1692_),
    .A(net82),
    .Y(_0666_));
 sg13g2_o21ai_1 _3478_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_1723_),
    .A2(_0665_));
 sg13g2_nand2_1 _3479_ (.Y(_0668_),
    .A(net156),
    .B(_0667_));
 sg13g2_nor2_1 _3480_ (.A(_1935_),
    .B(_0232_),
    .Y(_0669_));
 sg13g2_nand3_1 _3481_ (.B(_0240_),
    .C(_1723_),
    .A(_1558_),
    .Y(_0670_));
 sg13g2_nand3_1 _3482_ (.B(_0244_),
    .C(_0670_),
    .A(net120),
    .Y(_0671_));
 sg13g2_a221oi_1 _3483_ (.B2(_0669_),
    .C1(_0671_),
    .B1(_0668_),
    .A1(_0660_),
    .Y(_0672_),
    .A2(_0664_));
 sg13g2_nor3_1 _3484_ (.A(_1916_),
    .B(_1887_),
    .C(net20),
    .Y(_0673_));
 sg13g2_nand2b_1 _3485_ (.Y(_0674_),
    .B(_0216_),
    .A_N(_0212_));
 sg13g2_and2_1 _3486_ (.A(net95),
    .B(_0674_),
    .X(_0675_));
 sg13g2_o21ai_1 _3487_ (.B1(net52),
    .Y(_0676_),
    .A1(_1771_),
    .A2(net144));
 sg13g2_a21oi_1 _3488_ (.A1(net16),
    .A2(_0676_),
    .Y(_0677_),
    .B1(_1709_));
 sg13g2_a21oi_1 _3489_ (.A1(_0216_),
    .A2(_0677_),
    .Y(_0678_),
    .B1(_1894_));
 sg13g2_nor4_1 _3490_ (.A(_1810_),
    .B(_0673_),
    .C(_0675_),
    .D(_0678_),
    .Y(_0679_));
 sg13g2_o21ai_1 _3491_ (.B1(net19),
    .Y(_0680_),
    .A1(_1703_),
    .A2(net117));
 sg13g2_nand4_1 _3492_ (.B(_0202_),
    .C(_0078_),
    .A(net114),
    .Y(_0681_),
    .D(_0204_));
 sg13g2_a21oi_1 _3493_ (.A1(net14),
    .A2(_0680_),
    .Y(_0682_),
    .B1(_0681_));
 sg13g2_nand2_1 _3494_ (.Y(_0684_),
    .A(net42),
    .B(_0515_));
 sg13g2_nand4_1 _3495_ (.B(net110),
    .C(_1821_),
    .A(net114),
    .Y(_0685_),
    .D(_0684_));
 sg13g2_nand3_1 _3496_ (.B(net169),
    .C(_0685_),
    .A(_1944_),
    .Y(_0686_));
 sg13g2_or4_1 _3497_ (.A(_0672_),
    .B(_0679_),
    .C(_0682_),
    .D(_0686_),
    .X(_0687_));
 sg13g2_nor2_1 _3498_ (.A(net17),
    .B(net64),
    .Y(_0688_));
 sg13g2_nor3_1 _3499_ (.A(_0190_),
    .B(net119),
    .C(_1880_),
    .Y(_0689_));
 sg13g2_o21ai_1 _3500_ (.B1(net86),
    .Y(_0690_),
    .A1(_0688_),
    .A2(_0689_));
 sg13g2_o21ai_1 _3501_ (.B1(net117),
    .Y(_0691_),
    .A1(net45),
    .A2(_0559_));
 sg13g2_nand4_1 _3502_ (.B(net63),
    .C(_0348_),
    .A(net115),
    .Y(_0692_),
    .D(_0691_));
 sg13g2_nand2_1 _3503_ (.Y(_0693_),
    .A(_1554_),
    .B(_1656_));
 sg13g2_nor3_1 _3504_ (.A(_1938_),
    .B(_0693_),
    .C(_0665_),
    .Y(_0695_));
 sg13g2_nor4_1 _3505_ (.A(_1795_),
    .B(_1833_),
    .C(_1982_),
    .D(_0323_),
    .Y(_0696_));
 sg13g2_nor3_1 _3506_ (.A(net114),
    .B(_0695_),
    .C(_0696_),
    .Y(_0697_));
 sg13g2_nor2_1 _3507_ (.A(_1639_),
    .B(_1893_),
    .Y(_0698_));
 sg13g2_a21oi_1 _3508_ (.A1(net17),
    .A2(_0309_),
    .Y(_0699_),
    .B1(_0693_));
 sg13g2_a21oi_1 _3509_ (.A1(_0349_),
    .A2(_0698_),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_nand4_1 _3510_ (.B(_0692_),
    .C(_0697_),
    .A(_0690_),
    .Y(_0701_),
    .D(_0700_));
 sg13g2_nand3_1 _3511_ (.B(net17),
    .C(_0309_),
    .A(_1604_),
    .Y(_0702_));
 sg13g2_nor3_2 _3512_ (.A(_1502_),
    .B(_1504_),
    .C(net96),
    .Y(_0703_));
 sg13g2_o21ai_1 _3513_ (.B1(_0703_),
    .Y(_0704_),
    .A1(net40),
    .A2(net150));
 sg13g2_nor2_1 _3514_ (.A(net109),
    .B(_1801_),
    .Y(_0706_));
 sg13g2_a22oi_1 _3515_ (.Y(_0707_),
    .B1(_0704_),
    .B2(_0706_),
    .A2(_0149_),
    .A1(_1661_));
 sg13g2_nand2b_1 _3516_ (.Y(_0708_),
    .B(_1820_),
    .A_N(_0304_));
 sg13g2_a21oi_1 _3517_ (.A1(_0702_),
    .A2(_0707_),
    .Y(_0709_),
    .B1(_0708_));
 sg13g2_nor4_1 _3518_ (.A(net118),
    .B(net168),
    .C(_0307_),
    .D(_0709_),
    .Y(_0710_));
 sg13g2_a21oi_1 _3519_ (.A1(_0701_),
    .A2(_0710_),
    .Y(_0711_),
    .B1(_0095_));
 sg13g2_o21ai_1 _3520_ (.B1(net66),
    .Y(_0712_),
    .A1(_1701_),
    .A2(net117));
 sg13g2_nand3_1 _3521_ (.B(net24),
    .C(_0712_),
    .A(net63),
    .Y(_0713_));
 sg13g2_nand2_1 _3522_ (.Y(_0714_),
    .A(net94),
    .B(_0713_));
 sg13g2_nand2_1 _3523_ (.Y(_0715_),
    .A(net116),
    .B(_0446_));
 sg13g2_a22oi_1 _3524_ (.Y(_0717_),
    .B1(net64),
    .B2(_1791_),
    .A2(_0122_),
    .A1(net102));
 sg13g2_nand3_1 _3525_ (.B(_0090_),
    .C(net42),
    .A(net74),
    .Y(_0718_));
 sg13g2_a22oi_1 _3526_ (.Y(_0719_),
    .B1(_0718_),
    .B2(_1798_),
    .A2(_0717_),
    .A1(_0715_));
 sg13g2_o21ai_1 _3527_ (.B1(_0491_),
    .Y(_0720_),
    .A1(_0714_),
    .A2(_0719_));
 sg13g2_nand2_1 _3528_ (.Y(_0721_),
    .A(net18),
    .B(_0099_));
 sg13g2_nand2_1 _3529_ (.Y(_0722_),
    .A(_1668_),
    .B(_1801_));
 sg13g2_a21oi_1 _3530_ (.A1(_0721_),
    .A2(_0722_),
    .Y(_0723_),
    .B1(net15));
 sg13g2_o21ai_1 _3531_ (.B1(net94),
    .Y(_0724_),
    .A1(_1595_),
    .A2(_0723_));
 sg13g2_a21oi_1 _3532_ (.A1(_0501_),
    .A2(_0724_),
    .Y(_0725_),
    .B1(net101));
 sg13g2_a21oi_1 _3533_ (.A1(_0720_),
    .A2(_0725_),
    .Y(_0726_),
    .B1(net69));
 sg13g2_o21ai_1 _3534_ (.B1(net89),
    .Y(_0728_),
    .A1(net61),
    .A2(net42));
 sg13g2_a21o_1 _3535_ (.A2(_0721_),
    .A1(_0277_),
    .B1(_0728_),
    .X(_0729_));
 sg13g2_o21ai_1 _3536_ (.B1(net98),
    .Y(_0730_),
    .A1(net103),
    .A2(_1953_));
 sg13g2_or2_1 _3537_ (.X(_0731_),
    .B(_0730_),
    .A(_1815_));
 sg13g2_a21oi_1 _3538_ (.A1(_1775_),
    .A2(_0397_),
    .Y(_0732_),
    .B1(_1603_));
 sg13g2_a221oi_1 _3539_ (.B2(net61),
    .C1(net107),
    .B1(_0603_),
    .A1(net139),
    .Y(_0733_),
    .A2(net99));
 sg13g2_a21oi_1 _3540_ (.A1(_1665_),
    .A2(_0732_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_a21oi_1 _3541_ (.A1(net28),
    .A2(_1703_),
    .Y(_0735_),
    .B1(_1864_));
 sg13g2_a21oi_1 _3542_ (.A1(_0274_),
    .A2(_0735_),
    .Y(_0736_),
    .B1(_1872_));
 sg13g2_nand4_1 _3543_ (.B(_0731_),
    .C(_0734_),
    .A(_0729_),
    .Y(_0737_),
    .D(_0736_));
 sg13g2_a22oi_1 _3544_ (.Y(_0739_),
    .B1(_0665_),
    .B2(_1665_),
    .A2(_1693_),
    .A1(_1689_));
 sg13g2_nand2_1 _3545_ (.Y(_0740_),
    .A(_0698_),
    .B(_0739_));
 sg13g2_a21o_1 _3546_ (.A2(_0608_),
    .A1(_1658_),
    .B1(_0392_),
    .X(_0741_));
 sg13g2_nand4_1 _3547_ (.B(_0737_),
    .C(_0740_),
    .A(net76),
    .Y(_0742_),
    .D(_0741_));
 sg13g2_and2_1 _3548_ (.A(_1552_),
    .B(_0131_),
    .X(_0743_));
 sg13g2_o21ai_1 _3549_ (.B1(net135),
    .Y(_0744_),
    .A1(net151),
    .A2(net124));
 sg13g2_a221oi_1 _3550_ (.B2(_0744_),
    .C1(_0630_),
    .B1(_0625_),
    .A1(_1829_),
    .Y(_0745_),
    .A2(_0743_));
 sg13g2_a21oi_1 _3551_ (.A1(_0466_),
    .A2(_0468_),
    .Y(_0746_),
    .B1(net135));
 sg13g2_nor3_1 _3552_ (.A(net135),
    .B(net31),
    .C(_0464_),
    .Y(_0747_));
 sg13g2_o21ai_1 _3553_ (.B1(_1534_),
    .Y(_0748_),
    .A1(net43),
    .A2(_1692_));
 sg13g2_a221oi_1 _3554_ (.B2(_0748_),
    .C1(net116),
    .B1(_0227_),
    .A1(net12),
    .Y(_0750_),
    .A2(_1625_));
 sg13g2_nor4_1 _3555_ (.A(net115),
    .B(_0746_),
    .C(_0747_),
    .D(_0750_),
    .Y(_0751_));
 sg13g2_a21oi_1 _3556_ (.A1(net16),
    .A2(_1925_),
    .Y(_0752_),
    .B1(net49));
 sg13g2_o21ai_1 _3557_ (.B1(net38),
    .Y(_0753_),
    .A1(_0703_),
    .A2(net44));
 sg13g2_o21ai_1 _3558_ (.B1(_0753_),
    .Y(_0754_),
    .A1(net13),
    .A2(_0752_));
 sg13g2_a21oi_1 _3559_ (.A1(net81),
    .A2(_0754_),
    .Y(_0755_),
    .B1(net88));
 sg13g2_o21ai_1 _3560_ (.B1(_0755_),
    .Y(_0756_),
    .A1(_0745_),
    .A2(_0751_));
 sg13g2_nand3_1 _3561_ (.B(_0742_),
    .C(_0756_),
    .A(net70),
    .Y(_0757_));
 sg13g2_a22oi_1 _3562_ (.Y(_0758_),
    .B1(_0726_),
    .B2(_0757_),
    .A2(_0711_),
    .A1(_0687_));
 sg13g2_or3_1 _3563_ (.A(_0511_),
    .B(_0656_),
    .C(_0758_),
    .X(_0759_));
 sg13g2_o21ai_1 _3564_ (.B1(net140),
    .Y(_0761_),
    .A1(net27),
    .A2(_1916_));
 sg13g2_a21oi_1 _3565_ (.A1(net37),
    .A2(net134),
    .Y(_0762_),
    .B1(net18));
 sg13g2_a221oi_1 _3566_ (.B2(_1456_),
    .C1(net90),
    .B1(_0762_),
    .A1(_1844_),
    .Y(_0763_),
    .A2(_0382_));
 sg13g2_o21ai_1 _3567_ (.B1(_0763_),
    .Y(_0764_),
    .A1(_0330_),
    .A2(_0761_));
 sg13g2_a21oi_1 _3568_ (.A1(_1593_),
    .A2(_0570_),
    .Y(_0765_),
    .B1(net31));
 sg13g2_a221oi_1 _3569_ (.B2(net150),
    .C1(_1938_),
    .B1(net66),
    .A1(net142),
    .Y(_0766_),
    .A2(net108));
 sg13g2_o21ai_1 _3570_ (.B1(net81),
    .Y(_0767_),
    .A1(_0765_),
    .A2(_0766_));
 sg13g2_nand3_1 _3571_ (.B(_1770_),
    .C(net134),
    .A(net126),
    .Y(_0768_));
 sg13g2_a21oi_1 _3572_ (.A1(_1606_),
    .A2(net18),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_mux2_1 _3573_ (.A0(_1686_),
    .A1(net56),
    .S(_0271_),
    .X(_0770_));
 sg13g2_a22oi_1 _3574_ (.Y(_0772_),
    .B1(_0770_),
    .B2(_1779_),
    .A2(_0769_),
    .A1(_0100_));
 sg13g2_a21oi_1 _3575_ (.A1(_1778_),
    .A2(net43),
    .Y(_0773_),
    .B1(net18));
 sg13g2_o21ai_1 _3576_ (.B1(net126),
    .Y(_0774_),
    .A1(_1702_),
    .A2(net134));
 sg13g2_a21oi_1 _3577_ (.A1(_0773_),
    .A2(_0774_),
    .Y(_0775_),
    .B1(net24));
 sg13g2_a21o_1 _3578_ (.A2(_0775_),
    .A1(_0772_),
    .B1(net122),
    .X(_0776_));
 sg13g2_nand4_1 _3579_ (.B(_0764_),
    .C(_0767_),
    .A(net92),
    .Y(_0777_),
    .D(_0776_));
 sg13g2_nand2_1 _3580_ (.Y(_0778_),
    .A(_1658_),
    .B(_0368_));
 sg13g2_nand2_1 _3581_ (.Y(_0779_),
    .A(net47),
    .B(_0467_));
 sg13g2_a221oi_1 _3582_ (.B2(_1665_),
    .C1(net125),
    .B1(_0779_),
    .A1(_1484_),
    .Y(_0780_),
    .A2(_1843_));
 sg13g2_or4_1 _3583_ (.A(_1810_),
    .B(_0778_),
    .C(_0780_),
    .D(_0367_),
    .X(_0781_));
 sg13g2_nand2_2 _3584_ (.Y(_0783_),
    .A(_0183_),
    .B(_0403_));
 sg13g2_nor2_1 _3585_ (.A(_0783_),
    .B(_0345_),
    .Y(_0784_));
 sg13g2_o21ai_1 _3586_ (.B1(_0219_),
    .Y(_0785_),
    .A1(_1982_),
    .A2(_0167_));
 sg13g2_a21oi_1 _3587_ (.A1(_1763_),
    .A2(_1947_),
    .Y(_0786_),
    .B1(_0397_));
 sg13g2_o21ai_1 _3588_ (.B1(_0277_),
    .Y(_0787_),
    .A1(net36),
    .A2(_0786_));
 sg13g2_a21oi_1 _3589_ (.A1(_0785_),
    .A2(_0787_),
    .Y(_0788_),
    .B1(_1730_));
 sg13g2_or2_1 _3590_ (.X(_0789_),
    .B(_0788_),
    .A(_0401_));
 sg13g2_nand4_1 _3591_ (.B(_0781_),
    .C(_0784_),
    .A(_0777_),
    .Y(_0790_),
    .D(_0789_));
 sg13g2_nor2_1 _3592_ (.A(_1761_),
    .B(_0783_),
    .Y(_0791_));
 sg13g2_nand3_1 _3593_ (.B(net152),
    .C(_0118_),
    .A(net79),
    .Y(_0792_));
 sg13g2_nand2b_1 _3594_ (.Y(_0794_),
    .B(net59),
    .A_N(_1662_));
 sg13g2_nand4_1 _3595_ (.B(_1609_),
    .C(_1770_),
    .A(_1608_),
    .Y(_0795_),
    .D(_1726_));
 sg13g2_o21ai_1 _3596_ (.B1(_0795_),
    .Y(_0796_),
    .A1(net55),
    .A2(_1725_));
 sg13g2_o21ai_1 _3597_ (.B1(net110),
    .Y(_0797_),
    .A1(net71),
    .A2(net152));
 sg13g2_a221oi_1 _3598_ (.B2(net28),
    .C1(_0797_),
    .B1(_0796_),
    .A1(_0792_),
    .Y(_0798_),
    .A2(_0794_));
 sg13g2_nand3b_1 _3599_ (.B(net118),
    .C(net132),
    .Y(_0799_),
    .A_N(_0798_));
 sg13g2_nor2_1 _3600_ (.A(_1602_),
    .B(_1861_),
    .Y(_0800_));
 sg13g2_a221oi_1 _3601_ (.B2(net49),
    .C1(net138),
    .B1(_0800_),
    .A1(net104),
    .Y(_0801_),
    .A2(_0320_));
 sg13g2_nand3_1 _3602_ (.B(_1926_),
    .C(_0768_),
    .A(net26),
    .Y(_0802_));
 sg13g2_a21oi_1 _3603_ (.A1(net17),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0584_));
 sg13g2_nor3_1 _3604_ (.A(net26),
    .B(net93),
    .C(_1786_),
    .Y(_0805_));
 sg13g2_nor3_1 _3605_ (.A(_0801_),
    .B(_0803_),
    .C(_0805_),
    .Y(_0806_));
 sg13g2_inv_1 _3606_ (.Y(_0807_),
    .A(_1758_));
 sg13g2_o21ai_1 _3607_ (.B1(_0807_),
    .Y(_0808_),
    .A1(_0799_),
    .A2(_0806_));
 sg13g2_nor4_1 _3608_ (.A(net88),
    .B(_1747_),
    .C(_1761_),
    .D(_0783_),
    .Y(_0809_));
 sg13g2_a221oi_1 _3609_ (.B2(_1860_),
    .C1(_1765_),
    .B1(_1899_),
    .A1(_1669_),
    .Y(_0810_),
    .A2(_1498_));
 sg13g2_nand3b_1 _3610_ (.B(_0474_),
    .C(_1829_),
    .Y(_0811_),
    .A_N(_0810_));
 sg13g2_and2_1 _3611_ (.A(net86),
    .B(_0811_),
    .X(_0812_));
 sg13g2_a221oi_1 _3612_ (.B2(_1686_),
    .C1(net82),
    .B1(net56),
    .A1(net60),
    .Y(_0813_),
    .A2(net123));
 sg13g2_nor2_1 _3613_ (.A(_0446_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_a21oi_2 _3614_ (.B1(_0810_),
    .Y(_0816_),
    .A2(_1686_),
    .A1(_0207_));
 sg13g2_a22oi_1 _3615_ (.Y(_0817_),
    .B1(_0744_),
    .B2(_0816_),
    .A2(_0814_),
    .A1(net64));
 sg13g2_nor3_1 _3616_ (.A(net125),
    .B(_0446_),
    .C(_0813_),
    .Y(_0818_));
 sg13g2_nor3_1 _3617_ (.A(net86),
    .B(_0444_),
    .C(_0818_),
    .Y(_0819_));
 sg13g2_a21oi_1 _3618_ (.A1(_0812_),
    .A2(_0817_),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_a22oi_1 _3619_ (.Y(_0821_),
    .B1(_0809_),
    .B2(_0820_),
    .A2(_0808_),
    .A1(_0791_));
 sg13g2_a21oi_1 _3620_ (.A1(_1771_),
    .A2(_0202_),
    .Y(_0822_),
    .B1(net59));
 sg13g2_nor4_1 _3621_ (.A(_1684_),
    .B(net72),
    .C(_0822_),
    .D(_0266_),
    .Y(_0823_));
 sg13g2_nor3_1 _3622_ (.A(_1534_),
    .B(_1866_),
    .C(_1684_),
    .Y(_0824_));
 sg13g2_a21oi_1 _3623_ (.A1(_0240_),
    .A2(_1723_),
    .Y(_0825_),
    .B1(net104));
 sg13g2_nor4_1 _3624_ (.A(net122),
    .B(_0823_),
    .C(_0824_),
    .D(_0825_),
    .Y(_0827_));
 sg13g2_nor3_1 _3625_ (.A(net23),
    .B(_0703_),
    .C(_0548_),
    .Y(_0828_));
 sg13g2_nor2_1 _3626_ (.A(net32),
    .B(_0703_),
    .Y(_0829_));
 sg13g2_nor3_1 _3627_ (.A(_1764_),
    .B(_0829_),
    .C(_1936_),
    .Y(_0830_));
 sg13g2_o21ai_1 _3628_ (.B1(_0271_),
    .Y(_0831_),
    .A1(_0828_),
    .A2(_0830_));
 sg13g2_nand2_1 _3629_ (.Y(_0832_),
    .A(net92),
    .B(_0232_));
 sg13g2_a21oi_1 _3630_ (.A1(_0235_),
    .A2(_0233_),
    .Y(_0833_),
    .B1(_0236_));
 sg13g2_nand3_1 _3631_ (.B(_0242_),
    .C(_0078_),
    .A(_0240_),
    .Y(_0834_));
 sg13g2_nand2_1 _3632_ (.Y(_0835_),
    .A(_1758_),
    .B(_0834_));
 sg13g2_a221oi_1 _3633_ (.B2(_0833_),
    .C1(_0835_),
    .B1(_0832_),
    .A1(_0827_),
    .Y(_0836_),
    .A2(_0831_));
 sg13g2_nand2_1 _3634_ (.Y(_0837_),
    .A(net70),
    .B(_1759_));
 sg13g2_a21o_1 _3635_ (.A2(_1568_),
    .A1(net100),
    .B1(_0127_),
    .X(_0838_));
 sg13g2_nand3_1 _3636_ (.B(_1586_),
    .C(_1590_),
    .A(net130),
    .Y(_0839_));
 sg13g2_nand3_1 _3637_ (.B(_1565_),
    .C(_1567_),
    .A(net126),
    .Y(_0840_));
 sg13g2_and3_1 _3638_ (.X(_0841_),
    .A(net50),
    .B(_0839_),
    .C(_0840_));
 sg13g2_a221oi_1 _3639_ (.B2(_0838_),
    .C1(_0841_),
    .B1(net38),
    .A1(net162),
    .Y(_0842_),
    .A2(net109));
 sg13g2_nand2_1 _3640_ (.Y(_0843_),
    .A(net104),
    .B(net20));
 sg13g2_nand4_1 _3641_ (.B(net68),
    .C(net60),
    .A(_1778_),
    .Y(_0844_),
    .D(net137));
 sg13g2_and3_1 _3642_ (.X(_0845_),
    .A(_1593_),
    .B(net89),
    .C(_0844_));
 sg13g2_a221oi_1 _3643_ (.B2(_1911_),
    .C1(net115),
    .B1(_0845_),
    .A1(_0842_),
    .Y(_0846_),
    .A2(_0843_));
 sg13g2_a21oi_1 _3644_ (.A1(net145),
    .A2(_0317_),
    .Y(_0848_),
    .B1(net30));
 sg13g2_nor3_1 _3645_ (.A(net124),
    .B(net20),
    .C(_0848_),
    .Y(_0849_));
 sg13g2_or2_1 _3646_ (.X(_0850_),
    .B(_1888_),
    .A(_1667_));
 sg13g2_a221oi_1 _3647_ (.B2(net151),
    .C1(_0850_),
    .B1(_0382_),
    .A1(_1516_),
    .Y(_0851_),
    .A2(net73));
 sg13g2_a21oi_1 _3648_ (.A1(_1608_),
    .A2(_1609_),
    .Y(_0852_),
    .B1(_1684_));
 sg13g2_o21ai_1 _3649_ (.B1(net28),
    .Y(_0853_),
    .A1(_1561_),
    .A2(_0852_));
 sg13g2_a21oi_1 _3650_ (.A1(net97),
    .A2(_0853_),
    .Y(_0854_),
    .B1(net80));
 sg13g2_nor4_1 _3651_ (.A(net122),
    .B(_0849_),
    .C(_0851_),
    .D(_0854_),
    .Y(_0855_));
 sg13g2_o21ai_1 _3652_ (.B1(net76),
    .Y(_0856_),
    .A1(_0846_),
    .A2(_0855_));
 sg13g2_nand3b_1 _3653_ (.B(_0837_),
    .C(_0856_),
    .Y(_0857_),
    .A_N(_0836_));
 sg13g2_a21oi_1 _3654_ (.A1(net67),
    .A2(_0087_),
    .Y(_0859_),
    .B1(_0423_));
 sg13g2_xnor2_1 _3655_ (.Y(_0860_),
    .A(net21),
    .B(_0859_));
 sg13g2_nand2_1 _3656_ (.Y(_0861_),
    .A(net64),
    .B(_0860_));
 sg13g2_o21ai_1 _3657_ (.B1(net16),
    .Y(_0862_),
    .A1(net22),
    .A2(net140));
 sg13g2_a21oi_1 _3658_ (.A1(_1908_),
    .A2(_0862_),
    .Y(_0863_),
    .B1(_1828_));
 sg13g2_o21ai_1 _3659_ (.B1(_0863_),
    .Y(_0864_),
    .A1(_1534_),
    .A2(_0762_));
 sg13g2_nand2_1 _3660_ (.Y(_0865_),
    .A(net28),
    .B(net51));
 sg13g2_nand4_1 _3661_ (.B(_0865_),
    .C(_0105_),
    .A(net39),
    .Y(_0866_),
    .D(_0131_));
 sg13g2_a21oi_1 _3662_ (.A1(_0744_),
    .A2(_0866_),
    .Y(_0867_),
    .B1(net86));
 sg13g2_nand3_1 _3663_ (.B(_0864_),
    .C(_0867_),
    .A(_0861_),
    .Y(_0868_));
 sg13g2_o21ai_1 _3664_ (.B1(net97),
    .Y(_0870_),
    .A1(net38),
    .A2(_0452_));
 sg13g2_or2_1 _3665_ (.X(_0871_),
    .B(_0127_),
    .A(net130));
 sg13g2_o21ai_1 _3666_ (.B1(net122),
    .Y(_0872_),
    .A1(_0115_),
    .A2(_0871_));
 sg13g2_a21oi_1 _3667_ (.A1(net63),
    .A2(_0870_),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_nor3_1 _3668_ (.A(net88),
    .B(net118),
    .C(_0873_),
    .Y(_0874_));
 sg13g2_a21oi_1 _3669_ (.A1(_1833_),
    .A2(_0816_),
    .Y(_0875_),
    .B1(net115));
 sg13g2_nand2_1 _3670_ (.Y(_0876_),
    .A(_1552_),
    .B(_0305_));
 sg13g2_a22oi_1 _3671_ (.Y(_0877_),
    .B1(_0860_),
    .B2(net63),
    .A2(_0876_),
    .A1(net95));
 sg13g2_and2_1 _3672_ (.A(net121),
    .B(_0312_),
    .X(_0878_));
 sg13g2_nand2_1 _3673_ (.Y(_0879_),
    .A(net88),
    .B(net101));
 sg13g2_a221oi_1 _3674_ (.B2(_0187_),
    .C1(_0879_),
    .B1(_0878_),
    .A1(_0875_),
    .Y(_0881_),
    .A2(_0877_));
 sg13g2_a221oi_1 _3675_ (.B2(_0874_),
    .C1(_0881_),
    .B1(_0868_),
    .A1(_0807_),
    .Y(_0882_),
    .A2(net168));
 sg13g2_a22oi_1 _3676_ (.Y(_0883_),
    .B1(_0857_),
    .B2(_0882_),
    .A2(_0821_),
    .A1(_0790_));
 sg13g2_xnor2_1 _3677_ (.Y(_0884_),
    .A(_0607_),
    .B(_0957_));
 sg13g2_or3_1 _3678_ (.A(net197),
    .B(_0979_),
    .C(_0884_),
    .X(_0885_));
 sg13g2_nand3_1 _3679_ (.B(_0979_),
    .C(_0884_),
    .A(net197),
    .Y(_0886_));
 sg13g2_nand2_1 _3680_ (.Y(_0887_),
    .A(_1750_),
    .B(_1756_));
 sg13g2_inv_2 _3681_ (.Y(_0888_),
    .A(_0990_));
 sg13g2_nor2_1 _3682_ (.A(net199),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_nand3_1 _3683_ (.B(_0887_),
    .C(_0889_),
    .A(_1752_),
    .Y(_0890_));
 sg13g2_a21oi_1 _3684_ (.A1(_0885_),
    .A2(_0886_),
    .Y(_0892_),
    .B1(_0890_));
 sg13g2_nand3_1 _3685_ (.B(_0968_),
    .C(_0884_),
    .A(net197),
    .Y(_0893_));
 sg13g2_nand3b_1 _3686_ (.B(_0979_),
    .C(_0884_),
    .Y(_0894_),
    .A_N(net197));
 sg13g2_nor2_1 _3687_ (.A(_1734_),
    .B(_1735_),
    .Y(_0895_));
 sg13g2_nand2_1 _3688_ (.Y(_0896_),
    .A(_0902_),
    .B(_0895_));
 sg13g2_nand2_1 _3689_ (.Y(_0897_),
    .A(_0990_),
    .B(_1752_));
 sg13g2_inv_1 _3690_ (.Y(_0898_),
    .A(net199));
 sg13g2_nand2_1 _3691_ (.Y(_0899_),
    .A(_0898_),
    .B(_1752_));
 sg13g2_nor2_1 _3692_ (.A(net180),
    .B(_0895_),
    .Y(_0900_));
 sg13g2_a221oi_1 _3693_ (.B2(_0899_),
    .C1(_0900_),
    .B1(_0897_),
    .A1(net182),
    .Y(_0901_),
    .A2(_0896_));
 sg13g2_nand3_1 _3694_ (.B(_0888_),
    .C(_1750_),
    .A(net199),
    .Y(_0903_));
 sg13g2_inv_1 _3695_ (.Y(_0904_),
    .A(_0903_));
 sg13g2_nand3_1 _3696_ (.B(_0896_),
    .C(_0904_),
    .A(net182),
    .Y(_0905_));
 sg13g2_nor3_1 _3697_ (.A(net180),
    .B(_0895_),
    .C(_0903_),
    .Y(_0906_));
 sg13g2_a21oi_1 _3698_ (.A1(net199),
    .A2(_0888_),
    .Y(_0907_),
    .B1(_1750_));
 sg13g2_nor3_1 _3699_ (.A(_0898_),
    .B(_0990_),
    .C(_1752_),
    .Y(_0908_));
 sg13g2_nor4_1 _3700_ (.A(_0889_),
    .B(_0906_),
    .C(_0907_),
    .D(_0908_),
    .Y(_0909_));
 sg13g2_nand3b_1 _3701_ (.B(_0905_),
    .C(_0909_),
    .Y(_0910_),
    .A_N(_0901_));
 sg13g2_a21oi_1 _3702_ (.A1(_0893_),
    .A2(_0894_),
    .Y(_0911_),
    .B1(_0910_));
 sg13g2_or2_1 _3703_ (.X(_0912_),
    .B(_0911_),
    .A(_0892_));
 sg13g2_nand2_1 _3704_ (.Y(_0914_),
    .A(_1241_),
    .B(_0793_));
 sg13g2_nor2_1 _3705_ (.A(_1241_),
    .B(_0793_),
    .Y(_0915_));
 sg13g2_nor2_1 _3706_ (.A(_0760_),
    .B(_1489_),
    .Y(_0916_));
 sg13g2_nand2_1 _3707_ (.Y(_0917_),
    .A(net181),
    .B(_1489_));
 sg13g2_o21ai_1 _3708_ (.B1(_0917_),
    .Y(_0918_),
    .A1(_1242_),
    .A2(_0916_));
 sg13g2_or2_1 _3709_ (.X(_0919_),
    .B(_0918_),
    .A(_0915_));
 sg13g2_buf_1 _3710_ (.A(_0919_),
    .X(_0920_));
 sg13g2_xnor2_1 _3711_ (.Y(_0921_),
    .A(_1236_),
    .B(_0683_));
 sg13g2_buf_2 _3712_ (.A(_0921_),
    .X(_0922_));
 sg13g2_nor2_1 _3713_ (.A(net193),
    .B(_0705_),
    .Y(_0923_));
 sg13g2_nand3b_1 _3714_ (.B(_0923_),
    .C(_1246_),
    .Y(_0925_),
    .A_N(_0922_));
 sg13g2_nor2b_1 _3715_ (.A(_0705_),
    .B_N(net193),
    .Y(_0926_));
 sg13g2_inv_1 _3716_ (.Y(_0927_),
    .A(_1245_));
 sg13g2_nor2_1 _3717_ (.A(_1244_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nand3_1 _3718_ (.B(_0926_),
    .C(_0928_),
    .A(_0922_),
    .Y(_0929_));
 sg13g2_a22oi_1 _3719_ (.Y(_0930_),
    .B1(_0925_),
    .B2(_0929_),
    .A2(_0920_),
    .A1(_0914_));
 sg13g2_nand3_1 _3720_ (.B(_1253_),
    .C(_0922_),
    .A(_0727_),
    .Y(_0931_));
 sg13g2_nor2b_1 _3721_ (.A(_1245_),
    .B_N(_1244_),
    .Y(_0932_));
 sg13g2_nand4_1 _3722_ (.B(_0705_),
    .C(_0922_),
    .A(net193),
    .Y(_0933_),
    .D(_0932_));
 sg13g2_a22oi_1 _3723_ (.Y(_0934_),
    .B1(_0931_),
    .B2(_0933_),
    .A2(_0920_),
    .A1(_0914_));
 sg13g2_nand3_1 _3724_ (.B(_0922_),
    .C(_0923_),
    .A(_1253_),
    .Y(_0936_));
 sg13g2_nand3_1 _3725_ (.B(_0926_),
    .C(_0932_),
    .A(_0922_),
    .Y(_0937_));
 sg13g2_nand2_1 _3726_ (.Y(_0938_),
    .A(_0914_),
    .B(_0920_));
 sg13g2_a21oi_1 _3727_ (.A1(_0936_),
    .A2(_0937_),
    .Y(_0939_),
    .B1(_0938_));
 sg13g2_nand3_1 _3728_ (.B(_0922_),
    .C(_0928_),
    .A(_0727_),
    .Y(_0940_));
 sg13g2_nand4_1 _3729_ (.B(_0705_),
    .C(_1246_),
    .A(net193),
    .Y(_0941_),
    .D(_0922_));
 sg13g2_a21oi_1 _3730_ (.A1(_0940_),
    .A2(_0941_),
    .Y(_0942_),
    .B1(_0938_));
 sg13g2_or4_1 _3731_ (.A(_0930_),
    .B(_0934_),
    .C(_0939_),
    .D(_0942_),
    .X(_0943_));
 sg13g2_a21oi_1 _3732_ (.A1(_0912_),
    .A2(_0943_),
    .Y(_0944_),
    .B1(net1));
 sg13g2_o21ai_1 _3733_ (.B1(_1780_),
    .Y(_0945_),
    .A1(_0277_),
    .A2(_1728_));
 sg13g2_a21oi_1 _3734_ (.A1(_1723_),
    .A2(_0945_),
    .Y(_0947_),
    .B1(_0636_));
 sg13g2_nand2_1 _3735_ (.Y(_0948_),
    .A(_1794_),
    .B(_0271_));
 sg13g2_a221oi_1 _3736_ (.B2(_0948_),
    .C1(_1821_),
    .B1(_0548_),
    .A1(net40),
    .Y(_0949_),
    .A2(net28));
 sg13g2_a221oi_1 _3737_ (.B2(_1847_),
    .C1(net27),
    .B1(_1684_),
    .A1(net22),
    .Y(_0950_),
    .A2(net97));
 sg13g2_nor4_1 _3738_ (.A(_1856_),
    .B(_1975_),
    .C(_0949_),
    .D(_0950_),
    .Y(_0951_));
 sg13g2_nor3_1 _3739_ (.A(_0162_),
    .B(_0947_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_nor3_1 _3740_ (.A(net158),
    .B(_1803_),
    .C(_0234_),
    .Y(_0953_));
 sg13g2_nor3_1 _3741_ (.A(_1730_),
    .B(_0953_),
    .C(_0232_),
    .Y(_0954_));
 sg13g2_nand2b_1 _3742_ (.Y(_0955_),
    .B(_1873_),
    .A_N(_0954_));
 sg13g2_nand3_1 _3743_ (.B(_0189_),
    .C(net149),
    .A(net26),
    .Y(_0956_));
 sg13g2_nand4_1 _3744_ (.B(_1617_),
    .C(_1915_),
    .A(net19),
    .Y(_0958_),
    .D(_0956_));
 sg13g2_nand3b_1 _3745_ (.B(_0958_),
    .C(_1630_),
    .Y(_0959_),
    .A_N(_0828_));
 sg13g2_a21oi_1 _3746_ (.A1(_1906_),
    .A2(_1823_),
    .Y(_0960_),
    .B1(_1775_));
 sg13g2_a221oi_1 _3747_ (.B2(_0960_),
    .C1(_1893_),
    .B1(_1915_),
    .A1(_1517_),
    .Y(_0961_),
    .A2(_1706_));
 sg13g2_nor3_1 _3748_ (.A(_0249_),
    .B(_1918_),
    .C(_0961_),
    .Y(_0962_));
 sg13g2_nand2_1 _3749_ (.Y(_0963_),
    .A(_0959_),
    .B(_0962_));
 sg13g2_nor2_1 _3750_ (.A(net86),
    .B(_0851_),
    .Y(_0964_));
 sg13g2_a21oi_1 _3751_ (.A1(net159),
    .A2(_1690_),
    .Y(_0965_),
    .B1(_1561_));
 sg13g2_o21ai_1 _3752_ (.B1(net97),
    .Y(_0966_),
    .A1(net35),
    .A2(_0965_));
 sg13g2_o21ai_1 _3753_ (.B1(_0189_),
    .Y(_0967_),
    .A1(net161),
    .A2(_1670_));
 sg13g2_a221oi_1 _3754_ (.B2(_0967_),
    .C1(_1696_),
    .B1(net34),
    .A1(net35),
    .Y(_0969_),
    .A2(net97));
 sg13g2_a21oi_1 _3755_ (.A1(net102),
    .A2(_0966_),
    .Y(_0970_),
    .B1(_0969_));
 sg13g2_a21oi_1 _3756_ (.A1(_0964_),
    .A2(_0970_),
    .Y(_0971_),
    .B1(net92));
 sg13g2_a221oi_1 _3757_ (.B2(_0971_),
    .C1(net70),
    .B1(_0963_),
    .A1(_0952_),
    .Y(_0972_),
    .A2(_0955_));
 sg13g2_nor3_1 _3758_ (.A(_0127_),
    .B(_0572_),
    .C(_0573_),
    .Y(_0973_));
 sg13g2_nor3_1 _3759_ (.A(net124),
    .B(net45),
    .C(_0813_),
    .Y(_0974_));
 sg13g2_o21ai_1 _3760_ (.B1(_0974_),
    .Y(_0975_),
    .A1(_1718_),
    .A2(_0973_));
 sg13g2_o21ai_1 _3761_ (.B1(net46),
    .Y(_0976_),
    .A1(_1772_),
    .A2(_1953_));
 sg13g2_nand4_1 _3762_ (.B(net19),
    .C(_1617_),
    .A(_1659_),
    .Y(_0977_),
    .D(_0976_));
 sg13g2_or3_1 _3763_ (.A(net156),
    .B(net19),
    .C(_0859_),
    .X(_0978_));
 sg13g2_nand4_1 _3764_ (.B(_0975_),
    .C(_0977_),
    .A(net81),
    .Y(_0980_),
    .D(_0978_));
 sg13g2_nor2_1 _3765_ (.A(net81),
    .B(_0816_),
    .Y(_0981_));
 sg13g2_nor2_1 _3766_ (.A(net92),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_o21ai_1 _3767_ (.B1(net16),
    .Y(_0983_),
    .A1(net30),
    .A2(_0467_));
 sg13g2_nand2_1 _3768_ (.Y(_0984_),
    .A(net97),
    .B(_0983_));
 sg13g2_o21ai_1 _3769_ (.B1(_1540_),
    .Y(_0985_),
    .A1(_1926_),
    .A2(_1844_));
 sg13g2_a21oi_1 _3770_ (.A1(net46),
    .A2(_0985_),
    .Y(_0986_),
    .B1(_0127_));
 sg13g2_o21ai_1 _3771_ (.B1(_1604_),
    .Y(_0987_),
    .A1(net158),
    .A2(_1910_));
 sg13g2_a221oi_1 _3772_ (.B2(_0987_),
    .C1(_0249_),
    .B1(_0986_),
    .A1(_1805_),
    .Y(_0988_),
    .A2(_0984_));
 sg13g2_a221oi_1 _3773_ (.B2(net72),
    .C1(net132),
    .B1(_0445_),
    .A1(net46),
    .Y(_0989_),
    .A2(_1908_));
 sg13g2_a21oi_1 _3774_ (.A1(_0347_),
    .A2(_0989_),
    .Y(_0991_),
    .B1(_1832_));
 sg13g2_o21ai_1 _3775_ (.B1(net101),
    .Y(_0992_),
    .A1(_0988_),
    .A2(_0991_));
 sg13g2_a21oi_1 _3776_ (.A1(_0980_),
    .A2(_0982_),
    .Y(_0993_),
    .B1(_0992_));
 sg13g2_nor4_1 _3777_ (.A(_0098_),
    .B(_0783_),
    .C(_0972_),
    .D(_0993_),
    .Y(_0994_));
 sg13g2_nor2_1 _3778_ (.A(_1697_),
    .B(_1810_),
    .Y(_0995_));
 sg13g2_nor2_1 _3779_ (.A(_0778_),
    .B(_0780_),
    .Y(_0996_));
 sg13g2_a21oi_1 _3780_ (.A1(net66),
    .A2(_0493_),
    .Y(_0997_),
    .B1(_1815_));
 sg13g2_nor3_1 _3781_ (.A(net116),
    .B(_1607_),
    .C(_0997_),
    .Y(_0998_));
 sg13g2_o21ai_1 _3782_ (.B1(net60),
    .Y(_0999_),
    .A1(_0139_),
    .A2(_1804_));
 sg13g2_a221oi_1 _3783_ (.B2(_0999_),
    .C1(net126),
    .B1(_1625_),
    .A1(net30),
    .Y(_1000_),
    .A2(_1516_));
 sg13g2_nand3_1 _3784_ (.B(net100),
    .C(_0493_),
    .A(net82),
    .Y(_1002_));
 sg13g2_nor2_1 _3785_ (.A(net135),
    .B(net52),
    .Y(_1003_));
 sg13g2_a221oi_1 _3786_ (.B2(_1003_),
    .C1(net141),
    .B1(_1002_),
    .A1(net95),
    .Y(_1004_),
    .A2(_0316_));
 sg13g2_nand2b_1 _3787_ (.Y(_1005_),
    .B(_1004_),
    .A_N(_1000_));
 sg13g2_nor2_1 _3788_ (.A(net82),
    .B(_0087_),
    .Y(_1006_));
 sg13g2_nor3_1 _3789_ (.A(net59),
    .B(net29),
    .C(_0358_),
    .Y(_1007_));
 sg13g2_nor2_1 _3790_ (.A(net126),
    .B(net43),
    .Y(_1008_));
 sg13g2_o21ai_1 _3791_ (.B1(_1008_),
    .Y(_1009_),
    .A1(_1006_),
    .A2(_1007_));
 sg13g2_nand4_1 _3792_ (.B(net52),
    .C(net58),
    .A(net50),
    .Y(_1010_),
    .D(net137));
 sg13g2_nand3_1 _3793_ (.B(net105),
    .C(_1010_),
    .A(_1552_),
    .Y(_1011_));
 sg13g2_nand3_1 _3794_ (.B(_0502_),
    .C(net72),
    .A(net107),
    .Y(_1013_));
 sg13g2_nand4_1 _3795_ (.B(_1009_),
    .C(_1011_),
    .A(net122),
    .Y(_1014_),
    .D(_1013_));
 sg13g2_o21ai_1 _3796_ (.B1(_1014_),
    .Y(_1015_),
    .A1(_0998_),
    .A2(_1005_));
 sg13g2_and2_1 _3797_ (.A(_1520_),
    .B(_0795_),
    .X(_1016_));
 sg13g2_o21ai_1 _3798_ (.B1(_1016_),
    .Y(_1017_),
    .A1(net36),
    .A2(_0786_));
 sg13g2_nand4_1 _3799_ (.B(_1599_),
    .C(_0785_),
    .A(_1392_),
    .Y(_1018_),
    .D(_1017_));
 sg13g2_nor4_1 _3800_ (.A(net118),
    .B(_1758_),
    .C(_0094_),
    .D(_0783_),
    .Y(_1019_));
 sg13g2_o21ai_1 _3801_ (.B1(net33),
    .Y(_1020_),
    .A1(net47),
    .A2(_1853_));
 sg13g2_nand4_1 _3802_ (.B(_1938_),
    .C(_0078_),
    .A(net132),
    .Y(_1021_),
    .D(_1020_));
 sg13g2_nand3_1 _3803_ (.B(_1019_),
    .C(_1021_),
    .A(_1018_),
    .Y(_1022_));
 sg13g2_a221oi_1 _3804_ (.B2(_1523_),
    .C1(_1022_),
    .B1(_1015_),
    .A1(_0995_),
    .Y(_1024_),
    .A2(_0996_));
 sg13g2_nand3_1 _3805_ (.B(_0183_),
    .C(_0403_),
    .A(_0095_),
    .Y(_1025_));
 sg13g2_o21ai_1 _3806_ (.B1(_1625_),
    .Y(_1026_),
    .A1(_1603_),
    .A2(_0261_));
 sg13g2_a21oi_1 _3807_ (.A1(net17),
    .A2(_1026_),
    .Y(_1027_),
    .B1(_1720_));
 sg13g2_nor3_1 _3808_ (.A(net106),
    .B(_0805_),
    .C(_1027_),
    .Y(_1028_));
 sg13g2_nor3_1 _3809_ (.A(_1965_),
    .B(_0382_),
    .C(_0805_),
    .Y(_1029_));
 sg13g2_nor4_1 _3810_ (.A(_0799_),
    .B(_1025_),
    .C(_1028_),
    .D(_1029_),
    .Y(_1030_));
 sg13g2_inv_1 _3811_ (.Y(_1031_),
    .A(_0607_));
 sg13g2_o21ai_1 _3812_ (.B1(_0683_),
    .Y(_1032_),
    .A1(net193),
    .A2(_0705_));
 sg13g2_nand4_1 _3813_ (.B(_0847_),
    .C(_0585_),
    .A(_1031_),
    .Y(_1033_),
    .D(_1032_));
 sg13g2_o21ai_1 _3814_ (.B1(net116),
    .Y(_1035_),
    .A1(_1646_),
    .A2(_1653_));
 sg13g2_a21o_1 _3815_ (.A2(_0084_),
    .A1(_0202_),
    .B1(net15),
    .X(_1036_));
 sg13g2_a21oi_1 _3816_ (.A1(_1035_),
    .A2(_1036_),
    .Y(_1037_),
    .B1(net94));
 sg13g2_a21oi_1 _3817_ (.A1(_0190_),
    .A2(_0090_),
    .Y(_1038_),
    .B1(_1499_));
 sg13g2_o21ai_1 _3818_ (.B1(net73),
    .Y(_1039_),
    .A1(_1772_),
    .A2(_0693_));
 sg13g2_a21oi_1 _3819_ (.A1(_1807_),
    .A2(_1039_),
    .Y(_1040_),
    .B1(net114));
 sg13g2_o21ai_1 _3820_ (.B1(_1040_),
    .Y(_1041_),
    .A1(net11),
    .A2(_1038_));
 sg13g2_nor4_1 _3821_ (.A(net101),
    .B(_1025_),
    .C(_1037_),
    .D(_1041_),
    .Y(_1042_));
 sg13g2_or4_1 _3822_ (.A(_1024_),
    .B(_1030_),
    .C(_1033_),
    .D(_1042_),
    .X(_1043_));
 sg13g2_or4_1 _3823_ (.A(_0883_),
    .B(_0944_),
    .C(_0994_),
    .D(_1043_),
    .X(_1044_));
 sg13g2_a221oi_1 _3824_ (.B2(_0759_),
    .C1(_1044_),
    .B1(_0510_),
    .A1(_1841_),
    .Y(_1046_),
    .A2(_0200_));
 sg13g2_buf_1 _3825_ (.A(_1046_),
    .X(_1047_));
 sg13g2_buf_1 _3826_ (.A(net2),
    .X(_1048_));
 sg13g2_xnor2_1 _3827_ (.Y(_1049_),
    .A(net102),
    .B(_0185_));
 sg13g2_nand2_1 _3828_ (.Y(_1050_),
    .A(\palette_inst.rrggbb[0] ),
    .B(net200));
 sg13g2_o21ai_1 _3829_ (.B1(_1050_),
    .Y(_1051_),
    .A1(net200),
    .A2(_1049_));
 sg13g2_and2_1 _3830_ (.A(_1047_),
    .B(_1051_),
    .X(_0015_));
 sg13g2_nand2_1 _3831_ (.Y(_1052_),
    .A(net160),
    .B(_1584_));
 sg13g2_xnor2_1 _3832_ (.Y(_1053_),
    .A(_1404_),
    .B(_1052_));
 sg13g2_xnor2_1 _3833_ (.Y(_1054_),
    .A(_1574_),
    .B(net77));
 sg13g2_nor2_1 _3834_ (.A(_0185_),
    .B(_1054_),
    .Y(_1056_));
 sg13g2_xor2_1 _3835_ (.B(_1056_),
    .A(_1053_),
    .X(_1057_));
 sg13g2_nand2_1 _3836_ (.Y(_1058_),
    .A(net200),
    .B(\palette_inst.rrggbb[1] ));
 sg13g2_o21ai_1 _3837_ (.B1(_1058_),
    .Y(_1059_),
    .A1(net200),
    .A2(_1057_));
 sg13g2_and2_1 _3838_ (.A(_1047_),
    .B(_1059_),
    .X(_0016_));
 sg13g2_o21ai_1 _3839_ (.B1(_1053_),
    .Y(_1060_),
    .A1(net130),
    .A2(_0185_));
 sg13g2_nand2_1 _3840_ (.Y(_1061_),
    .A(_1574_),
    .B(_1060_));
 sg13g2_nor2_1 _3841_ (.A(net126),
    .B(_0185_),
    .Y(_1062_));
 sg13g2_or2_1 _3842_ (.X(_1063_),
    .B(_1053_),
    .A(_1062_));
 sg13g2_buf_1 _3843_ (.A(_1063_),
    .X(_1064_));
 sg13g2_nand2_1 _3844_ (.Y(_1066_),
    .A(_1061_),
    .B(_1064_));
 sg13g2_nand2_1 _3845_ (.Y(_1067_),
    .A(_1187_),
    .B(_1052_));
 sg13g2_o21ai_1 _3846_ (.B1(_1067_),
    .Y(_1068_),
    .A1(net154),
    .A2(_1052_));
 sg13g2_nand2_1 _3847_ (.Y(_1069_),
    .A(_1430_),
    .B(_1434_));
 sg13g2_xnor2_1 _3848_ (.Y(_1070_),
    .A(_0771_),
    .B(_1069_));
 sg13g2_xnor2_1 _3849_ (.Y(_1071_),
    .A(net132),
    .B(_1070_));
 sg13g2_xor2_1 _3850_ (.B(_1071_),
    .A(_1068_),
    .X(_1072_));
 sg13g2_xnor2_1 _3851_ (.Y(_1073_),
    .A(_1066_),
    .B(_1072_));
 sg13g2_nand2_1 _3852_ (.Y(_1074_),
    .A(net200),
    .B(\palette_inst.rrggbb[2] ));
 sg13g2_o21ai_1 _3853_ (.B1(_1074_),
    .Y(_1075_),
    .A1(net200),
    .A2(_1073_));
 sg13g2_and2_1 _3854_ (.A(_1047_),
    .B(_1075_),
    .X(_0017_));
 sg13g2_nand3_1 _3855_ (.B(_1064_),
    .C(_1068_),
    .A(_1061_),
    .Y(_1077_));
 sg13g2_a21oi_1 _3856_ (.A1(_1061_),
    .A2(_1064_),
    .Y(_1078_),
    .B1(_1068_));
 sg13g2_a21o_1 _3857_ (.A2(_1077_),
    .A1(_1071_),
    .B1(_1078_),
    .X(_1079_));
 sg13g2_xnor2_1 _3858_ (.Y(_1080_),
    .A(net181),
    .B(_1489_));
 sg13g2_nor2_1 _3859_ (.A(net132),
    .B(_1070_),
    .Y(_1081_));
 sg13g2_a21oi_1 _3860_ (.A1(_1238_),
    .A2(_1070_),
    .Y(_1082_),
    .B1(_1081_));
 sg13g2_xnor2_1 _3861_ (.Y(_1083_),
    .A(_1080_),
    .B(_1082_));
 sg13g2_xnor2_1 _3862_ (.Y(_1084_),
    .A(net70),
    .B(_1083_));
 sg13g2_xnor2_1 _3863_ (.Y(_1085_),
    .A(_1079_),
    .B(_1084_));
 sg13g2_nand2_1 _3864_ (.Y(_1087_),
    .A(net200),
    .B(\palette_inst.rrggbb[3] ));
 sg13g2_o21ai_1 _3865_ (.B1(_1087_),
    .Y(_1088_),
    .A1(_1048_),
    .A2(_1085_));
 sg13g2_and2_1 _3866_ (.A(_1047_),
    .B(_1088_),
    .X(_0018_));
 sg13g2_nand2b_1 _3867_ (.Y(_1089_),
    .B(net200),
    .A_N(\palette_inst.rrggbb[4] ));
 sg13g2_nor2_1 _3868_ (.A(_1079_),
    .B(_1082_),
    .Y(_1090_));
 sg13g2_nand3_1 _3869_ (.B(net91),
    .C(_1090_),
    .A(net25),
    .Y(_1091_));
 sg13g2_or4_1 _3870_ (.A(net177),
    .B(net25),
    .C(net91),
    .D(_1090_),
    .X(_1092_));
 sg13g2_and2_1 _3871_ (.A(net177),
    .B(net25),
    .X(_1093_));
 sg13g2_and2_1 _3872_ (.A(net177),
    .B(net91),
    .X(_1094_));
 sg13g2_o21ai_1 _3873_ (.B1(_1090_),
    .Y(_1095_),
    .A1(_1093_),
    .A2(_1094_));
 sg13g2_nand3_1 _3874_ (.B(_1092_),
    .C(_1095_),
    .A(_1091_),
    .Y(_1097_));
 sg13g2_and2_1 _3875_ (.A(_1079_),
    .B(_1082_),
    .X(_1098_));
 sg13g2_nand3_1 _3876_ (.B(net70),
    .C(_1098_),
    .A(net14),
    .Y(_1099_));
 sg13g2_nand3b_1 _3877_ (.B(_1093_),
    .C(net91),
    .Y(_1100_),
    .A_N(_1098_));
 sg13g2_nor2_1 _3878_ (.A(_1243_),
    .B(net25),
    .Y(_1101_));
 sg13g2_nor2_1 _3879_ (.A(_1243_),
    .B(net91),
    .Y(_1102_));
 sg13g2_o21ai_1 _3880_ (.B1(_1098_),
    .Y(_1103_),
    .A1(_1101_),
    .A2(_1102_));
 sg13g2_nand3_1 _3881_ (.B(_1100_),
    .C(_1103_),
    .A(_1099_),
    .Y(_1104_));
 sg13g2_xnor2_1 _3882_ (.Y(_1105_),
    .A(_0793_),
    .B(_0918_));
 sg13g2_xnor2_1 _3883_ (.Y(_1106_),
    .A(net69),
    .B(_1105_));
 sg13g2_or4_1 _3884_ (.A(net2),
    .B(_1097_),
    .C(_1104_),
    .D(_1106_),
    .X(_1108_));
 sg13g2_nor2b_1 _3885_ (.A(net2),
    .B_N(_1106_),
    .Y(_1109_));
 sg13g2_o21ai_1 _3886_ (.B1(_1109_),
    .Y(_1110_),
    .A1(_1097_),
    .A2(_1104_));
 sg13g2_and4_1 _3887_ (.A(_1047_),
    .B(_1089_),
    .C(_1108_),
    .D(_1110_),
    .X(_0019_));
 sg13g2_nand2b_1 _3888_ (.Y(_1111_),
    .B(_1048_),
    .A_N(\palette_inst.rrggbb[5] ));
 sg13g2_and2_1 _3889_ (.A(_1047_),
    .B(_1111_),
    .X(_0020_));
 sg13g2_inv_1 _3890_ (.Y(_1112_),
    .A(_1278_));
 sg13g2_nand2_1 _3891_ (.Y(_1113_),
    .A(_0013_),
    .B(_1112_));
 sg13g2_nand2_1 _3892_ (.Y(_1114_),
    .A(\color_index[0] ),
    .B(_1278_));
 sg13g2_a21oi_1 _3893_ (.A1(_1113_),
    .A2(_1114_),
    .Y(_0021_),
    .B1(net184));
 sg13g2_nand2_1 _3894_ (.Y(_1116_),
    .A(\color_index[0] ),
    .B(_1112_));
 sg13g2_xnor2_1 _3895_ (.Y(_1117_),
    .A(\color_index[1] ),
    .B(_1116_));
 sg13g2_and2_1 _3896_ (.A(_1298_),
    .B(_1117_),
    .X(_0022_));
 sg13g2_nand2_1 _3897_ (.Y(_1118_),
    .A(\color_index[2] ),
    .B(_1278_));
 sg13g2_xor2_1 _3898_ (.B(_1279_),
    .A(_0007_),
    .X(_1119_));
 sg13g2_nand2_1 _3899_ (.Y(_1120_),
    .A(_1112_),
    .B(_1119_));
 sg13g2_a21oi_1 _3900_ (.A1(_1118_),
    .A2(_1120_),
    .Y(_0023_),
    .B1(net184));
 sg13g2_buf_1 _3901_ (.A(_1276_),
    .X(_1121_));
 sg13g2_buf_1 _3902_ (.A(_1170_),
    .X(_1122_));
 sg13g2_a21oi_1 _3903_ (.A1(net147),
    .A2(_1255_),
    .Y(_1123_),
    .B1(_1122_));
 sg13g2_buf_1 _3904_ (.A(_1276_),
    .X(_1125_));
 sg13g2_inv_2 _3905_ (.Y(_1126_),
    .A(net146));
 sg13g2_nor4_1 _3906_ (.A(_0006_),
    .B(_1126_),
    .C(_1235_),
    .D(_1248_),
    .Y(_1127_));
 sg13g2_o21ai_1 _3907_ (.B1(net191),
    .Y(_0024_),
    .A1(_1123_),
    .A2(_1127_));
 sg13g2_nor3_1 _3908_ (.A(_0009_),
    .B(_1126_),
    .C(_1096_),
    .Y(_1128_));
 sg13g2_buf_1 _3909_ (.A(_0869_),
    .X(_1129_));
 sg13g2_a21oi_1 _3910_ (.A1(net147),
    .A2(_1141_),
    .Y(_1130_),
    .B1(net172));
 sg13g2_nor3_1 _3911_ (.A(net184),
    .B(_1128_),
    .C(_1130_),
    .Y(_0025_));
 sg13g2_nand2_1 _3912_ (.Y(_1131_),
    .A(_0011_),
    .B(net147));
 sg13g2_nand2_1 _3913_ (.Y(_1132_),
    .A(net186),
    .B(_1126_));
 sg13g2_a21oi_1 _3914_ (.A1(_1131_),
    .A2(_1132_),
    .Y(_0026_),
    .B1(net184));
 sg13g2_xor2_1 _3915_ (.B(net173),
    .A(_0011_),
    .X(_1134_));
 sg13g2_nand2_1 _3916_ (.Y(_1135_),
    .A(net146),
    .B(_1134_));
 sg13g2_xor2_1 _3917_ (.B(_1135_),
    .A(net187),
    .X(_1136_));
 sg13g2_nor2_1 _3918_ (.A(net174),
    .B(_1136_),
    .Y(_0027_));
 sg13g2_nor3_1 _3919_ (.A(net187),
    .B(net186),
    .C(net173),
    .Y(_1137_));
 sg13g2_a21oi_1 _3920_ (.A1(net173),
    .A2(_1233_),
    .Y(_1138_),
    .B1(_1137_));
 sg13g2_nand2b_1 _3921_ (.Y(_1139_),
    .B(net146),
    .A_N(_1138_));
 sg13g2_xnor2_1 _3922_ (.Y(_1140_),
    .A(_1574_),
    .B(_1139_));
 sg13g2_nor2_1 _3923_ (.A(net174),
    .B(_1140_),
    .Y(_0028_));
 sg13g2_inv_1 _3924_ (.Y(_1142_),
    .A(net173));
 sg13g2_nor2_1 _3925_ (.A(_1206_),
    .B(net186),
    .Y(_1143_));
 sg13g2_o21ai_1 _3926_ (.B1(_1574_),
    .Y(_1144_),
    .A1(net173),
    .A2(_1143_));
 sg13g2_o21ai_1 _3927_ (.B1(_1144_),
    .Y(_1145_),
    .A1(_1142_),
    .A2(_1233_));
 sg13g2_xnor2_1 _3928_ (.Y(_1146_),
    .A(_1142_),
    .B(_1145_));
 sg13g2_nand2_1 _3929_ (.Y(_1147_),
    .A(net147),
    .B(_1146_));
 sg13g2_xnor2_1 _3930_ (.Y(_1148_),
    .A(_1250_),
    .B(_1147_));
 sg13g2_nand2_1 _3931_ (.Y(_0029_),
    .A(net191),
    .B(_1148_));
 sg13g2_buf_1 _3932_ (.A(net184),
    .X(_1149_));
 sg13g2_nor2_1 _3933_ (.A(net179),
    .B(_1197_),
    .Y(_1150_));
 sg13g2_nand2_1 _3934_ (.Y(_1152_),
    .A(_1150_),
    .B(_1137_));
 sg13g2_o21ai_1 _3935_ (.B1(_1152_),
    .Y(_1153_),
    .A1(_1142_),
    .A2(_1235_));
 sg13g2_nand2_1 _3936_ (.Y(_1154_),
    .A(net147),
    .B(_1153_));
 sg13g2_xnor2_1 _3937_ (.Y(_1155_),
    .A(_1239_),
    .B(_1154_));
 sg13g2_nor2_1 _3938_ (.A(net171),
    .B(_1155_),
    .Y(_0030_));
 sg13g2_a21oi_1 _3939_ (.A1(_1150_),
    .A2(_1143_),
    .Y(_1156_),
    .B1(net173));
 sg13g2_a21oi_1 _3940_ (.A1(net173),
    .A2(_1235_),
    .Y(_1157_),
    .B1(_1239_));
 sg13g2_nor2_1 _3941_ (.A(_1156_),
    .B(_1157_),
    .Y(_1158_));
 sg13g2_nor2_1 _3942_ (.A(_1142_),
    .B(_1158_),
    .Y(_1159_));
 sg13g2_nor2_1 _3943_ (.A(net178),
    .B(_1152_),
    .Y(_1160_));
 sg13g2_o21ai_1 _3944_ (.B1(net146),
    .Y(_1162_),
    .A1(_1159_),
    .A2(_1160_));
 sg13g2_xor2_1 _3945_ (.B(_1162_),
    .A(net177),
    .X(_1163_));
 sg13g2_nor2_1 _3946_ (.A(net171),
    .B(_1163_),
    .Y(_0031_));
 sg13g2_nor3_1 _3947_ (.A(net177),
    .B(net178),
    .C(_1152_),
    .Y(_1164_));
 sg13g2_a21oi_1 _3948_ (.A1(net177),
    .A2(_1159_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_nor2_1 _3949_ (.A(_1126_),
    .B(_1165_),
    .Y(_1166_));
 sg13g2_xnor2_1 _3950_ (.Y(_1167_),
    .A(_1241_),
    .B(_1166_));
 sg13g2_nand2_1 _3951_ (.Y(_0032_),
    .A(net191),
    .B(_1167_));
 sg13g2_nor2b_1 _3952_ (.A(_1252_),
    .B_N(_1145_),
    .Y(_1168_));
 sg13g2_nand4_1 _3953_ (.B(net177),
    .C(net178),
    .A(_1241_),
    .Y(_1169_),
    .D(_1122_));
 sg13g2_nor3_1 _3954_ (.A(_1250_),
    .B(_1145_),
    .C(_1169_),
    .Y(_1171_));
 sg13g2_o21ai_1 _3955_ (.B1(net146),
    .Y(_1172_),
    .A1(_1168_),
    .A2(_1171_));
 sg13g2_xnor2_1 _3956_ (.Y(_1173_),
    .A(_0927_),
    .B(_1172_));
 sg13g2_nand2_1 _3957_ (.Y(_0033_),
    .A(net191),
    .B(_1173_));
 sg13g2_mux2_1 _3958_ (.A0(_1168_),
    .A1(_1171_),
    .S(_1245_),
    .X(_1174_));
 sg13g2_nand2_1 _3959_ (.Y(_1175_),
    .A(net146),
    .B(_1174_));
 sg13g2_xor2_1 _3960_ (.B(_1175_),
    .A(_1244_),
    .X(_1176_));
 sg13g2_nor2_1 _3961_ (.A(net171),
    .B(_1176_),
    .Y(_0034_));
 sg13g2_nand3_1 _3962_ (.B(_1247_),
    .C(_1157_),
    .A(net173),
    .Y(_1177_));
 sg13g2_nand3_1 _3963_ (.B(_1253_),
    .C(_1158_),
    .A(_1251_),
    .Y(_1178_));
 sg13g2_a21oi_1 _3964_ (.A1(_1177_),
    .A2(_1178_),
    .Y(_1180_),
    .B1(_1126_));
 sg13g2_xnor2_1 _3965_ (.Y(_1181_),
    .A(_1236_),
    .B(_1180_));
 sg13g2_nor2_1 _3966_ (.A(net171),
    .B(_1181_),
    .Y(_0035_));
 sg13g2_nand2_1 _3967_ (.Y(_1182_),
    .A(_0913_),
    .B(net147));
 sg13g2_nand2_1 _3968_ (.Y(_1183_),
    .A(net188),
    .B(_1126_));
 sg13g2_a21oi_1 _3969_ (.A1(_1182_),
    .A2(_1183_),
    .Y(_0036_),
    .B1(net184));
 sg13g2_xor2_1 _3970_ (.B(net172),
    .A(_0913_),
    .X(_1184_));
 sg13g2_nand2_1 _3971_ (.Y(_1185_),
    .A(_1121_),
    .B(_1184_));
 sg13g2_xnor2_1 _3972_ (.Y(_1186_),
    .A(_1393_),
    .B(_1185_));
 sg13g2_nor2_1 _3973_ (.A(net171),
    .B(_1186_),
    .Y(_0037_));
 sg13g2_nand3_1 _3974_ (.B(_1065_),
    .C(net172),
    .A(net189),
    .Y(_1188_));
 sg13g2_nand2b_1 _3975_ (.Y(_1189_),
    .B(_1677_),
    .A_N(net172));
 sg13g2_a21oi_1 _3976_ (.A1(_1188_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_1126_));
 sg13g2_xnor2_1 _3977_ (.Y(_1191_),
    .A(_1045_),
    .B(_1190_));
 sg13g2_nor2_1 _3978_ (.A(net171),
    .B(_1191_),
    .Y(_0038_));
 sg13g2_o21ai_1 _3979_ (.B1(_0869_),
    .Y(_1192_),
    .A1(_1393_),
    .A2(_1107_));
 sg13g2_nor2_1 _3980_ (.A(_0869_),
    .B(_1677_),
    .Y(_1193_));
 sg13g2_a21oi_1 _3981_ (.A1(_1045_),
    .A2(_1192_),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_xor2_1 _3982_ (.B(_1194_),
    .A(net172),
    .X(_1195_));
 sg13g2_a21oi_1 _3983_ (.A1(net147),
    .A2(_1195_),
    .Y(_1196_),
    .B1(net190));
 sg13g2_and3_1 _3984_ (.X(_1198_),
    .A(net190),
    .B(net147),
    .C(_1195_));
 sg13g2_o21ai_1 _3985_ (.B1(net191),
    .Y(_0039_),
    .A1(_1196_),
    .A2(_1198_));
 sg13g2_nor2_1 _3986_ (.A(net188),
    .B(_1129_),
    .Y(_1199_));
 sg13g2_a22oi_1 _3987_ (.Y(_1200_),
    .B1(_1133_),
    .B2(_1199_),
    .A2(_1086_),
    .A1(_1129_));
 sg13g2_nor2_1 _3988_ (.A(_1126_),
    .B(_1200_),
    .Y(_1201_));
 sg13g2_xnor2_1 _3989_ (.Y(_1202_),
    .A(_1001_),
    .B(_1201_));
 sg13g2_nor2_1 _3990_ (.A(net171),
    .B(_1202_),
    .Y(_0040_));
 sg13g2_a21oi_1 _3991_ (.A1(_1107_),
    .A2(_1133_),
    .Y(_1203_),
    .B1(_0869_));
 sg13g2_a21oi_1 _3992_ (.A1(_0869_),
    .A2(_1076_),
    .Y(_1204_),
    .B1(_1012_));
 sg13g2_nor2_2 _3993_ (.A(_1203_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_xor2_1 _3994_ (.B(_1205_),
    .A(net172),
    .X(_1207_));
 sg13g2_nand2_1 _3995_ (.Y(_1208_),
    .A(net146),
    .B(_1207_));
 sg13g2_xor2_1 _3996_ (.B(_1208_),
    .A(net180),
    .X(_1209_));
 sg13g2_nor2_1 _3997_ (.A(net171),
    .B(_1209_),
    .Y(_0041_));
 sg13g2_and2_1 _3998_ (.A(net180),
    .B(_0869_),
    .X(_1210_));
 sg13g2_nor2_1 _3999_ (.A(net180),
    .B(net172),
    .Y(_1211_));
 sg13g2_mux2_1 _4000_ (.A0(_1210_),
    .A1(_1211_),
    .S(_1205_),
    .X(_1212_));
 sg13g2_nand2_1 _4001_ (.Y(_1213_),
    .A(net146),
    .B(_1212_));
 sg13g2_xor2_1 _4002_ (.B(_1213_),
    .A(_0880_),
    .X(_1214_));
 sg13g2_nand2_1 _4003_ (.Y(_0042_),
    .A(net191),
    .B(_1214_));
 sg13g2_nand2_1 _4004_ (.Y(_1216_),
    .A(_0880_),
    .B(_1210_));
 sg13g2_nand2_1 _4005_ (.Y(_1217_),
    .A(_1001_),
    .B(net190));
 sg13g2_nor3_1 _4006_ (.A(_1194_),
    .B(_1216_),
    .C(_1217_),
    .Y(_1218_));
 sg13g2_nor2_1 _4007_ (.A(net190),
    .B(net172),
    .Y(_1219_));
 sg13g2_and3_1 _4008_ (.X(_1220_),
    .A(_1124_),
    .B(_1194_),
    .C(_1219_));
 sg13g2_o21ai_1 _4009_ (.B1(_1125_),
    .Y(_1221_),
    .A1(_1218_),
    .A2(_1220_));
 sg13g2_xnor2_1 _4010_ (.Y(_1222_),
    .A(_0888_),
    .B(_1221_));
 sg13g2_nand2_1 _4011_ (.Y(_0043_),
    .A(net191),
    .B(_1222_));
 sg13g2_mux2_1 _4012_ (.A0(_1218_),
    .A1(_1220_),
    .S(_0888_),
    .X(_1223_));
 sg13g2_nand2_1 _4013_ (.Y(_1224_),
    .A(_1121_),
    .B(_1223_));
 sg13g2_xnor2_1 _4014_ (.Y(_1226_),
    .A(_0979_),
    .B(_1224_));
 sg13g2_nor2_1 _4015_ (.A(_1149_),
    .B(_1226_),
    .Y(_0044_));
 sg13g2_nor3_1 _4016_ (.A(_0979_),
    .B(_0888_),
    .C(_1216_),
    .Y(_1227_));
 sg13g2_nor3_1 _4017_ (.A(_0968_),
    .B(_0990_),
    .C(_0880_),
    .Y(_1228_));
 sg13g2_and2_1 _4018_ (.A(_1211_),
    .B(_1228_),
    .X(_1229_));
 sg13g2_mux2_1 _4019_ (.A0(_1227_),
    .A1(_1229_),
    .S(_1205_),
    .X(_1230_));
 sg13g2_nand2_1 _4020_ (.Y(_1231_),
    .A(_1125_),
    .B(_1230_));
 sg13g2_xor2_1 _4021_ (.B(_1231_),
    .A(_0957_),
    .X(_1232_));
 sg13g2_nor2_1 _4022_ (.A(_1149_),
    .B(_1232_),
    .Y(_0045_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \B[0]$_SDFF_PN0__217  (.L_HI(net217));
 sg13g2_buf_1 _4025_ (.A(net201),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4026_ (.A(net202),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4027_ (.A(net203),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4028_ (.A(net204),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4029_ (.A(net205),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4030_ (.A(net206),
    .X(uio_oe[5]));
 sg13g2_buf_1 _4031_ (.A(net207),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4032_ (.A(net208),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4033_ (.A(net209),
    .X(uio_out[0]));
 sg13g2_buf_1 _4034_ (.A(net210),
    .X(uio_out[1]));
 sg13g2_buf_1 _4035_ (.A(net211),
    .X(uio_out[2]));
 sg13g2_buf_1 _4036_ (.A(net212),
    .X(uio_out[3]));
 sg13g2_buf_1 _4037_ (.A(net213),
    .X(uio_out[4]));
 sg13g2_buf_1 _4038_ (.A(net214),
    .X(uio_out[5]));
 sg13g2_buf_1 _4039_ (.A(net215),
    .X(uio_out[6]));
 sg13g2_buf_1 _4040_ (.A(net216),
    .X(uio_out[7]));
 sg13g2_buf_1 _4041_ (.A(\vga_sync_gen.vsync ),
    .X(net6));
 sg13g2_buf_1 _4042_ (.A(hsync),
    .X(net10));
 sg13g2_dfrbp_1 \color_index[0]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net223),
    .D(_0021_),
    .Q_N(_0013_),
    .Q(\color_index[0] ));
 sg13g2_dfrbp_1 \color_index[1]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net224),
    .D(_0022_),
    .Q_N(_0008_),
    .Q(\color_index[1] ));
 sg13g2_dfrbp_1 \color_index[2]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net225),
    .D(_0023_),
    .Q_N(_0007_),
    .Q(\color_index[2] ));
 sg13g2_dfrbp_1 \dir_x$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net226),
    .D(_0024_),
    .Q_N(_0006_),
    .Q(dir_x));
 sg13g2_dfrbp_1 \dir_y$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net227),
    .D(_0025_),
    .Q_N(_0009_),
    .Q(dir_y));
 sg13g2_dfrbp_1 \logo_left[0]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net228),
    .D(_0026_),
    .Q_N(_0011_),
    .Q(\logo_left[0] ));
 sg13g2_dfrbp_1 \logo_left[1]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net229),
    .D(_0027_),
    .Q_N(_2032_),
    .Q(\logo_left[1] ));
 sg13g2_dfrbp_1 \logo_left[2]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net230),
    .D(_0028_),
    .Q_N(_2031_),
    .Q(\logo_left[2] ));
 sg13g2_dfrbp_1 \logo_left[3]$_SDFFE_PN1P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net231),
    .D(_0029_),
    .Q_N(_2030_),
    .Q(\logo_left[3] ));
 sg13g2_dfrbp_1 \logo_left[4]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net232),
    .D(_0030_),
    .Q_N(_2029_),
    .Q(\logo_left[4] ));
 sg13g2_dfrbp_1 \logo_left[5]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net233),
    .D(_0031_),
    .Q_N(_2028_),
    .Q(\logo_left[5] ));
 sg13g2_dfrbp_1 \logo_left[6]$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net234),
    .D(_0032_),
    .Q_N(_2027_),
    .Q(\logo_left[6] ));
 sg13g2_dfrbp_1 \logo_left[7]$_SDFFE_PN1P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net235),
    .D(_0033_),
    .Q_N(_2026_),
    .Q(\logo_left[7] ));
 sg13g2_dfrbp_1 \logo_left[8]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net236),
    .D(_0034_),
    .Q_N(_2025_),
    .Q(\logo_left[8] ));
 sg13g2_dfrbp_1 \logo_left[9]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net237),
    .D(_0035_),
    .Q_N(_2024_),
    .Q(\logo_left[9] ));
 sg13g2_dfrbp_1 \logo_top[0]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net238),
    .D(_0036_),
    .Q_N(_0012_),
    .Q(\logo_top[0] ));
 sg13g2_dfrbp_1 \logo_top[1]$_SDFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net239),
    .D(_0037_),
    .Q_N(_2023_),
    .Q(\logo_top[1] ));
 sg13g2_dfrbp_1 \logo_top[2]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net240),
    .D(_0038_),
    .Q_N(_2022_),
    .Q(\logo_top[2] ));
 sg13g2_dfrbp_1 \logo_top[3]$_SDFFE_PN1P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net241),
    .D(_0039_),
    .Q_N(_2021_),
    .Q(\logo_top[3] ));
 sg13g2_dfrbp_1 \logo_top[4]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net242),
    .D(_0040_),
    .Q_N(_2020_),
    .Q(\logo_top[4] ));
 sg13g2_dfrbp_1 \logo_top[5]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net243),
    .D(_0041_),
    .Q_N(_2019_),
    .Q(\logo_top[5] ));
 sg13g2_dfrbp_1 \logo_top[6]$_SDFFE_PN1P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net244),
    .D(_0042_),
    .Q_N(_2018_),
    .Q(\logo_top[6] ));
 sg13g2_dfrbp_1 \logo_top[7]$_SDFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net245),
    .D(_0043_),
    .Q_N(_2017_),
    .Q(\logo_top[7] ));
 sg13g2_dfrbp_1 \logo_top[8]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net246),
    .D(_0044_),
    .Q_N(_2016_),
    .Q(\logo_top[8] ));
 sg13g2_dfrbp_1 \logo_top[9]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net247),
    .D(_0045_),
    .Q_N(_2039_),
    .Q(\logo_top[9] ));
 sg13g2_dfrbp_1 \pallete_color[0]$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net248),
    .D(_0000_),
    .Q_N(_2040_),
    .Q(\palette_inst.rrggbb[0] ));
 sg13g2_dfrbp_1 \pallete_color[1]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net249),
    .D(_0001_),
    .Q_N(_2041_),
    .Q(\palette_inst.rrggbb[1] ));
 sg13g2_dfrbp_1 \pallete_color[2]$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net250),
    .D(_0002_),
    .Q_N(_2042_),
    .Q(\palette_inst.rrggbb[2] ));
 sg13g2_dfrbp_1 \pallete_color[3]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net251),
    .D(_0003_),
    .Q_N(_2015_),
    .Q(\palette_inst.rrggbb[3] ));
 sg13g2_dfrbp_1 \pallete_color[4]$_SDFF_PP1_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net252),
    .D(_0046_),
    .Q_N(_2014_),
    .Q(\palette_inst.rrggbb[4] ));
 sg13g2_dfrbp_1 \pallete_color[5]$_SDFF_PP1_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net253),
    .D(_0047_),
    .Q_N(_2013_),
    .Q(\palette_inst.rrggbb[5] ));
 sg13g2_dfrbp_1 \prev_y[0]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net254),
    .D(_0048_),
    .Q_N(_2012_),
    .Q(\prev_y[0] ));
 sg13g2_dfrbp_1 \prev_y[1]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net255),
    .D(_0049_),
    .Q_N(_2011_),
    .Q(\prev_y[1] ));
 sg13g2_dfrbp_1 \prev_y[2]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net256),
    .D(_0050_),
    .Q_N(_2010_),
    .Q(\prev_y[2] ));
 sg13g2_dfrbp_1 \prev_y[3]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net257),
    .D(_0051_),
    .Q_N(_2009_),
    .Q(\prev_y[3] ));
 sg13g2_dfrbp_1 \prev_y[4]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net258),
    .D(_0052_),
    .Q_N(_2008_),
    .Q(\prev_y[4] ));
 sg13g2_dfrbp_1 \prev_y[5]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net259),
    .D(_0053_),
    .Q_N(_2007_),
    .Q(\prev_y[5] ));
 sg13g2_dfrbp_1 \prev_y[6]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net260),
    .D(_0054_),
    .Q_N(_2006_),
    .Q(\prev_y[6] ));
 sg13g2_dfrbp_1 \prev_y[7]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net261),
    .D(_0055_),
    .Q_N(_2005_),
    .Q(\prev_y[7] ));
 sg13g2_dfrbp_1 \prev_y[8]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net262),
    .D(_0056_),
    .Q_N(_2004_),
    .Q(\prev_y[8] ));
 sg13g2_dfrbp_1 \prev_y[9]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net263),
    .D(_0057_),
    .Q_N(_2003_),
    .Q(\prev_y[9] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net264),
    .D(_0058_),
    .Q_N(_0014_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net265),
    .D(_0059_),
    .Q_N(_2002_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net266),
    .D(_0060_),
    .Q_N(_2001_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net267),
    .D(_0061_),
    .Q_N(_2000_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net268),
    .D(_0062_),
    .Q_N(_1999_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net269),
    .D(_0063_),
    .Q_N(_1998_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net270),
    .D(_0064_),
    .Q_N(_1997_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net271),
    .D(_0065_),
    .Q_N(_1996_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net272),
    .D(_0066_),
    .Q_N(_1995_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net273),
    .D(_0067_),
    .Q_N(_2043_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 \vga_sync_gen.hsync$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net274),
    .D(_0004_),
    .Q_N(_1994_),
    .Q(hsync));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net275),
    .D(_0068_),
    .Q_N(_0010_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net276),
    .D(_0069_),
    .Q_N(_1993_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net277),
    .D(_0070_),
    .Q_N(_1992_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net278),
    .D(_0071_),
    .Q_N(_1991_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net279),
    .D(_0072_),
    .Q_N(_1990_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net280),
    .D(_0073_),
    .Q_N(_1989_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net281),
    .D(_0074_),
    .Q_N(_1988_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net282),
    .D(_0075_),
    .Q_N(_1987_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net283),
    .D(_0076_),
    .Q_N(_1986_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net284),
    .D(_0077_),
    .Q_N(_2044_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 \vga_sync_gen.vsync$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net285),
    .D(_0005_),
    .Q_N(_1985_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout11 (.A(_1818_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_1780_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_1720_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_1718_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1562_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0219_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_1981_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_1968_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_1927_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1910_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1864_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1817_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1813_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1807_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1798_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1774_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1717_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1701_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1670_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1615_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1594_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1561_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1525_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1517_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1508_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1484_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0325_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0149_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0099_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1926_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1906_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1900_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1869_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1801_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1791_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1779_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1775_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1766_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1764_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1716_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1709_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1690_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1669_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1614_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1583_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1582_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1560_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1507_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1493_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1483_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0207_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0122_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1975_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1833_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1778_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1772_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1765_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1763_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1759_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1748_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1725_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1712_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1706_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1703_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1671_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1644_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1630_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1623_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1611_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1604_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1600_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1520_),
    .X(net82));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_1509_));
 sg13g2_buf_2 fanout84 (.A(_1492_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1482_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0392_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0189_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0162_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0111_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1965_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1945_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1924_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1916_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1914_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1875_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1860_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1846_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1805_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1789_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1771_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1747_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1730_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1702_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1661_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1656_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1640_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1629_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1609_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1603_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1599_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1592_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_1543_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_1519_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_1392_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0249_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0090_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1978_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1944_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1917_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_1882_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_1872_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1856_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_1770_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_1696_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_1668_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_1660_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1652_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1639_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1619_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1602_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1532_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1391_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_1318_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_1947_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1893_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1859_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1823_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1795_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_1788_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_1769_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_1638_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_1608_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_1579_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_1557_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1540_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_1125_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_1121_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_1887_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_1768_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_1727_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_1700_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_1634_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_1621_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_1554_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_1511_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_1707_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_1691_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_1659_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_1606_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_1430_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_1421_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_1626_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_1605_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_1477_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_1458_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_1420_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_1407_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0094_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_1761_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_1423_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_1149_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_1129_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_1122_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_1292_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_1267_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_1264_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_1243_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_1238_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_1187_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_0902_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_0760_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_0541_),
    .X(net182));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_1298_));
 sg13g2_buf_2 fanout184 (.A(_1291_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_1242_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_1215_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_1206_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_1065_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_1055_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_1034_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_0858_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_0771_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_0694_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_0640_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_0629_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_0596_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_0574_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_0563_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_0552_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_1048_),
    .X(net200));
 sg13g2_tielo _4025__201 (.L_LO(net201));
 sg13g2_tielo _4026__202 (.L_LO(net202));
 sg13g2_tielo _4027__203 (.L_LO(net203));
 sg13g2_tielo _4028__204 (.L_LO(net204));
 sg13g2_tielo _4029__205 (.L_LO(net205));
 sg13g2_tielo _4030__206 (.L_LO(net206));
 sg13g2_tielo _4031__207 (.L_LO(net207));
 sg13g2_tielo _4032__208 (.L_LO(net208));
 sg13g2_tielo _4033__209 (.L_LO(net209));
 sg13g2_tielo _4034__210 (.L_LO(net210));
 sg13g2_tielo _4035__211 (.L_LO(net211));
 sg13g2_tielo _4036__212 (.L_LO(net212));
 sg13g2_tielo _4037__213 (.L_LO(net213));
 sg13g2_tielo _4038__214 (.L_LO(net214));
 sg13g2_tielo _4039__215 (.L_LO(net215));
 sg13g2_tielo _4040__216 (.L_LO(net216));
 sg13g2_tiehi \B[1]$_SDFF_PN0__218  (.L_HI(net218));
 sg13g2_tiehi \G[0]$_SDFF_PN0__219  (.L_HI(net219));
 sg13g2_tiehi \G[1]$_SDFF_PN0__220  (.L_HI(net220));
 sg13g2_tiehi \R[0]$_SDFF_PN0__221  (.L_HI(net221));
 sg13g2_tiehi \R[1]$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \color_index[0]$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \color_index[1]$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \color_index[2]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \dir_x$_SDFFE_PN1P__226  (.L_HI(net226));
 sg13g2_tiehi \dir_y$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \logo_left[0]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \logo_left[1]$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \logo_left[2]$_SDFFE_PN0P__230  (.L_HI(net230));
 sg13g2_tiehi \logo_left[3]$_SDFFE_PN1P__231  (.L_HI(net231));
 sg13g2_tiehi \logo_left[4]$_SDFFE_PN0P__232  (.L_HI(net232));
 sg13g2_tiehi \logo_left[5]$_SDFFE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \logo_left[6]$_SDFFE_PN1P__234  (.L_HI(net234));
 sg13g2_tiehi \logo_left[7]$_SDFFE_PN1P__235  (.L_HI(net235));
 sg13g2_tiehi \logo_left[8]$_SDFFE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \logo_left[9]$_SDFFE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \logo_top[0]$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \logo_top[1]$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \logo_top[2]$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \logo_top[3]$_SDFFE_PN1P__241  (.L_HI(net241));
 sg13g2_tiehi \logo_top[4]$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \logo_top[5]$_SDFFE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \logo_top[6]$_SDFFE_PN1P__244  (.L_HI(net244));
 sg13g2_tiehi \logo_top[7]$_SDFFE_PN1P__245  (.L_HI(net245));
 sg13g2_tiehi \logo_top[8]$_SDFFE_PN0P__246  (.L_HI(net246));
 sg13g2_tiehi \logo_top[9]$_SDFFE_PN0P__247  (.L_HI(net247));
 sg13g2_tiehi \pallete_color[0]$_DFF_P__248  (.L_HI(net248));
 sg13g2_tiehi \pallete_color[1]$_DFF_P__249  (.L_HI(net249));
 sg13g2_tiehi \pallete_color[2]$_DFF_P__250  (.L_HI(net250));
 sg13g2_tiehi \pallete_color[3]$_DFF_P__251  (.L_HI(net251));
 sg13g2_tiehi \pallete_color[4]$_SDFF_PP1__252  (.L_HI(net252));
 sg13g2_tiehi \pallete_color[5]$_SDFF_PP1__253  (.L_HI(net253));
 sg13g2_tiehi \prev_y[0]$_DFFE_PP__254  (.L_HI(net254));
 sg13g2_tiehi \prev_y[1]$_DFFE_PP__255  (.L_HI(net255));
 sg13g2_tiehi \prev_y[2]$_DFFE_PP__256  (.L_HI(net256));
 sg13g2_tiehi \prev_y[3]$_DFFE_PP__257  (.L_HI(net257));
 sg13g2_tiehi \prev_y[4]$_DFFE_PP__258  (.L_HI(net258));
 sg13g2_tiehi \prev_y[5]$_DFFE_PP__259  (.L_HI(net259));
 sg13g2_tiehi \prev_y[6]$_DFFE_PP__260  (.L_HI(net260));
 sg13g2_tiehi \prev_y[7]$_DFFE_PP__261  (.L_HI(net261));
 sg13g2_tiehi \prev_y[8]$_DFFE_PP__262  (.L_HI(net262));
 sg13g2_tiehi \prev_y[9]$_DFFE_PP__263  (.L_HI(net263));
 sg13g2_tiehi \vga_sync_gen.hpos[0]$_SDFF_PP0__264  (.L_HI(net264));
 sg13g2_tiehi \vga_sync_gen.hpos[1]$_SDFF_PP0__265  (.L_HI(net265));
 sg13g2_tiehi \vga_sync_gen.hpos[2]$_SDFF_PP0__266  (.L_HI(net266));
 sg13g2_tiehi \vga_sync_gen.hpos[3]$_SDFF_PP0__267  (.L_HI(net267));
 sg13g2_tiehi \vga_sync_gen.hpos[4]$_SDFF_PP0__268  (.L_HI(net268));
 sg13g2_tiehi \vga_sync_gen.hpos[5]$_SDFF_PP0__269  (.L_HI(net269));
 sg13g2_tiehi \vga_sync_gen.hpos[6]$_SDFF_PP0__270  (.L_HI(net270));
 sg13g2_tiehi \vga_sync_gen.hpos[7]$_SDFF_PP0__271  (.L_HI(net271));
 sg13g2_tiehi \vga_sync_gen.hpos[8]$_SDFF_PP0__272  (.L_HI(net272));
 sg13g2_tiehi \vga_sync_gen.hpos[9]$_SDFF_PP0__273  (.L_HI(net273));
 sg13g2_tiehi \vga_sync_gen.hsync$_DFF_P__274  (.L_HI(net274));
 sg13g2_tiehi \vga_sync_gen.vpos[0]$_SDFFCE_PP0P__275  (.L_HI(net275));
 sg13g2_tiehi \vga_sync_gen.vpos[1]$_SDFFCE_PP0P__276  (.L_HI(net276));
 sg13g2_tiehi \vga_sync_gen.vpos[2]$_SDFFCE_PP0P__277  (.L_HI(net277));
 sg13g2_tiehi \vga_sync_gen.vpos[3]$_SDFFCE_PP0P__278  (.L_HI(net278));
 sg13g2_tiehi \vga_sync_gen.vpos[4]$_SDFFCE_PP0P__279  (.L_HI(net279));
 sg13g2_tiehi \vga_sync_gen.vpos[5]$_SDFFCE_PP0P__280  (.L_HI(net280));
 sg13g2_tiehi \vga_sync_gen.vpos[6]$_SDFFCE_PP0P__281  (.L_HI(net281));
 sg13g2_tiehi \vga_sync_gen.vpos[7]$_SDFFCE_PP0P__282  (.L_HI(net282));
 sg13g2_tiehi \vga_sync_gen.vpos[8]$_SDFFCE_PP0P__283  (.L_HI(net283));
 sg13g2_tiehi \vga_sync_gen.vpos[9]$_SDFFCE_PP0P__284  (.L_HI(net284));
 sg13g2_tiehi \vga_sync_gen.vsync$_DFF_P__285  (.L_HI(net285));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0004_));
 sg13g2_antennanp ANTENNA_2 (.A(_1015_));
 sg13g2_antennanp ANTENNA_3 (.A(_1015_));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(_0004_));
 sg13g2_antennanp ANTENNA_7 (.A(clk));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(_0004_));
 sg13g2_antennanp ANTENNA_10 (.A(clk));
 sg13g2_antennanp ANTENNA_11 (.A(clk));
 sg13g2_antennanp ANTENNA_12 (.A(_0004_));
 sg13g2_antennanp ANTENNA_13 (.A(clk));
 sg13g2_antennanp ANTENNA_14 (.A(clk));
 sg13g2_antennanp ANTENNA_15 (.A(_0004_));
 sg13g2_antennanp ANTENNA_16 (.A(clk));
 sg13g2_antennanp ANTENNA_17 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_fill_1 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_96 ();
 sg13g2_decap_8 FILLER_1_103 ();
 sg13g2_decap_8 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_fill_2 FILLER_1_124 ();
 sg13g2_fill_1 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_131 ();
 sg13g2_decap_8 FILLER_1_138 ();
 sg13g2_fill_2 FILLER_1_154 ();
 sg13g2_fill_1 FILLER_1_156 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_4 FILLER_2_77 ();
 sg13g2_decap_4 FILLER_2_111 ();
 sg13g2_fill_1 FILLER_2_115 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_fill_2 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_222 ();
 sg13g2_decap_8 FILLER_2_229 ();
 sg13g2_decap_8 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_243 ();
 sg13g2_decap_8 FILLER_2_250 ();
 sg13g2_decap_8 FILLER_2_257 ();
 sg13g2_decap_8 FILLER_2_264 ();
 sg13g2_decap_8 FILLER_2_271 ();
 sg13g2_decap_8 FILLER_2_278 ();
 sg13g2_decap_8 FILLER_2_285 ();
 sg13g2_decap_8 FILLER_2_292 ();
 sg13g2_decap_8 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_306 ();
 sg13g2_decap_8 FILLER_2_313 ();
 sg13g2_decap_8 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_4 FILLER_3_77 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_86 ();
 sg13g2_decap_8 FILLER_3_93 ();
 sg13g2_decap_8 FILLER_3_100 ();
 sg13g2_decap_8 FILLER_3_111 ();
 sg13g2_decap_8 FILLER_3_118 ();
 sg13g2_decap_8 FILLER_3_125 ();
 sg13g2_decap_8 FILLER_3_132 ();
 sg13g2_decap_8 FILLER_3_139 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_4 FILLER_3_161 ();
 sg13g2_fill_1 FILLER_3_165 ();
 sg13g2_decap_4 FILLER_3_170 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_fill_2 FILLER_3_191 ();
 sg13g2_fill_1 FILLER_3_193 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_decap_8 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_253 ();
 sg13g2_decap_8 FILLER_3_260 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_decap_8 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_85 ();
 sg13g2_decap_8 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_99 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_137 ();
 sg13g2_decap_4 FILLER_4_151 ();
 sg13g2_fill_1 FILLER_4_155 ();
 sg13g2_decap_4 FILLER_4_160 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_fill_1 FILLER_4_204 ();
 sg13g2_fill_2 FILLER_4_222 ();
 sg13g2_fill_1 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_234 ();
 sg13g2_decap_8 FILLER_4_241 ();
 sg13g2_decap_8 FILLER_4_248 ();
 sg13g2_decap_8 FILLER_4_255 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_4 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_fill_1 FILLER_5_114 ();
 sg13g2_fill_2 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_176 ();
 sg13g2_fill_1 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_fill_2 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_4 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_311 ();
 sg13g2_fill_2 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_decap_8 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_5_414 ();
 sg13g2_decap_8 FILLER_5_421 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_111 ();
 sg13g2_decap_8 FILLER_6_120 ();
 sg13g2_decap_8 FILLER_6_127 ();
 sg13g2_decap_4 FILLER_6_134 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_decap_4 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_157 ();
 sg13g2_decap_8 FILLER_6_164 ();
 sg13g2_decap_4 FILLER_6_171 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_fill_1 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_decap_8 FILLER_6_212 ();
 sg13g2_decap_8 FILLER_6_219 ();
 sg13g2_decap_8 FILLER_6_226 ();
 sg13g2_decap_8 FILLER_6_233 ();
 sg13g2_decap_4 FILLER_6_240 ();
 sg13g2_fill_2 FILLER_6_253 ();
 sg13g2_fill_1 FILLER_6_255 ();
 sg13g2_decap_4 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_fill_1 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_88 ();
 sg13g2_decap_4 FILLER_7_95 ();
 sg13g2_fill_1 FILLER_7_99 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_4 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_143 ();
 sg13g2_decap_8 FILLER_7_150 ();
 sg13g2_decap_8 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_164 ();
 sg13g2_fill_2 FILLER_7_171 ();
 sg13g2_fill_1 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_7_190 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_223 ();
 sg13g2_decap_4 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_decap_4 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_254 ();
 sg13g2_decap_8 FILLER_7_261 ();
 sg13g2_decap_8 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_282 ();
 sg13g2_decap_4 FILLER_7_289 ();
 sg13g2_fill_1 FILLER_7_293 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_4 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_decap_4 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_4 FILLER_8_95 ();
 sg13g2_decap_4 FILLER_8_142 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_fill_1 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_fill_2 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_4 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_fill_2 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_fill_1 FILLER_8_291 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_4 FILLER_8_374 ();
 sg13g2_fill_1 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_415 ();
 sg13g2_decap_8 FILLER_8_422 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_89 ();
 sg13g2_decap_8 FILLER_9_96 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_fill_1 FILLER_9_110 ();
 sg13g2_decap_8 FILLER_9_115 ();
 sg13g2_decap_4 FILLER_9_134 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_171 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_decap_4 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_4 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_264 ();
 sg13g2_fill_2 FILLER_9_293 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_1 FILLER_9_351 ();
 sg13g2_fill_1 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_fill_1 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_4 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_8 FILLER_10_92 ();
 sg13g2_decap_4 FILLER_10_99 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_4 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_decap_4 FILLER_10_150 ();
 sg13g2_fill_1 FILLER_10_166 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_fill_2 FILLER_10_266 ();
 sg13g2_decap_4 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_358 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_4 FILLER_11_63 ();
 sg13g2_fill_1 FILLER_11_67 ();
 sg13g2_decap_4 FILLER_11_86 ();
 sg13g2_decap_8 FILLER_11_99 ();
 sg13g2_decap_8 FILLER_11_106 ();
 sg13g2_decap_8 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_120 ();
 sg13g2_decap_8 FILLER_11_127 ();
 sg13g2_fill_1 FILLER_11_138 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_decap_8 FILLER_11_152 ();
 sg13g2_fill_2 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_4 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_195 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_211 ();
 sg13g2_decap_8 FILLER_11_223 ();
 sg13g2_decap_4 FILLER_11_230 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_340 ();
 sg13g2_decap_4 FILLER_11_351 ();
 sg13g2_decap_4 FILLER_11_359 ();
 sg13g2_fill_1 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_decap_4 FILLER_12_87 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_decap_4 FILLER_12_96 ();
 sg13g2_decap_8 FILLER_12_108 ();
 sg13g2_decap_8 FILLER_12_115 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_135 ();
 sg13g2_decap_4 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_150 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_171 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_decap_8 FILLER_12_185 ();
 sg13g2_decap_8 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_decap_4 FILLER_12_252 ();
 sg13g2_fill_2 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_4 FILLER_12_326 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_4 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_351 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_fill_2 FILLER_12_372 ();
 sg13g2_fill_1 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_decap_8 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_414 ();
 sg13g2_decap_8 FILLER_12_421 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_4 FILLER_13_102 ();
 sg13g2_fill_2 FILLER_13_106 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_decap_4 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_159 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_4 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_fill_1 FILLER_13_310 ();
 sg13g2_decap_4 FILLER_13_316 ();
 sg13g2_decap_4 FILLER_13_330 ();
 sg13g2_decap_4 FILLER_13_339 ();
 sg13g2_fill_1 FILLER_13_343 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_351 ();
 sg13g2_fill_2 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_4 FILLER_13_375 ();
 sg13g2_fill_1 FILLER_13_379 ();
 sg13g2_fill_2 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_4 FILLER_14_67 ();
 sg13g2_fill_2 FILLER_14_71 ();
 sg13g2_decap_8 FILLER_14_118 ();
 sg13g2_decap_8 FILLER_14_125 ();
 sg13g2_decap_8 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_decap_4 FILLER_14_146 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_decap_4 FILLER_14_161 ();
 sg13g2_fill_2 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_4 FILLER_14_182 ();
 sg13g2_fill_1 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_204 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_fill_2 FILLER_14_217 ();
 sg13g2_decap_4 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_fill_1 FILLER_14_294 ();
 sg13g2_decap_4 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_317 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_fill_2 FILLER_14_344 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_4 FILLER_14_424 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_48 ();
 sg13g2_decap_4 FILLER_15_55 ();
 sg13g2_decap_4 FILLER_15_67 ();
 sg13g2_fill_1 FILLER_15_71 ();
 sg13g2_fill_2 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_216 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_4 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_269 ();
 sg13g2_decap_4 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_decap_4 FILLER_15_309 ();
 sg13g2_decap_4 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_330 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_93 ();
 sg13g2_fill_2 FILLER_16_101 ();
 sg13g2_fill_1 FILLER_16_141 ();
 sg13g2_decap_4 FILLER_16_146 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_decap_4 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_decap_4 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_246 ();
 sg13g2_decap_4 FILLER_16_259 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_4 FILLER_16_317 ();
 sg13g2_fill_1 FILLER_16_321 ();
 sg13g2_decap_4 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_decap_4 FILLER_16_346 ();
 sg13g2_decap_4 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_50 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_fill_1 FILLER_17_89 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_decap_8 FILLER_17_125 ();
 sg13g2_decap_8 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_139 ();
 sg13g2_decap_8 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_decap_8 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_decap_4 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_decap_4 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_decap_4 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_decap_4 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_4 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_decap_4 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_8 FILLER_17_404 ();
 sg13g2_decap_8 FILLER_17_411 ();
 sg13g2_decap_8 FILLER_17_418 ();
 sg13g2_decap_4 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_55 ();
 sg13g2_decap_8 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_fill_2 FILLER_18_80 ();
 sg13g2_fill_2 FILLER_18_87 ();
 sg13g2_fill_2 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_decap_8 FILLER_18_104 ();
 sg13g2_decap_8 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_decap_8 FILLER_18_132 ();
 sg13g2_decap_8 FILLER_18_139 ();
 sg13g2_decap_8 FILLER_18_146 ();
 sg13g2_decap_8 FILLER_18_153 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_decap_4 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_229 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_decap_4 FILLER_18_280 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_384 ();
 sg13g2_fill_1 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_159 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_decap_4 FILLER_19_281 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_290 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_decap_8 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_38 ();
 sg13g2_decap_8 FILLER_20_45 ();
 sg13g2_decap_8 FILLER_20_52 ();
 sg13g2_decap_4 FILLER_20_59 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_4 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_decap_4 FILLER_20_143 ();
 sg13g2_fill_2 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_170 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_288 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_4 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_decap_4 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_54 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_69 ();
 sg13g2_decap_8 FILLER_21_87 ();
 sg13g2_decap_4 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_106 ();
 sg13g2_decap_8 FILLER_21_113 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_decap_4 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_decap_4 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_4 FILLER_21_298 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_4 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_decap_4 FILLER_21_370 ();
 sg13g2_decap_4 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_78 ();
 sg13g2_decap_8 FILLER_22_85 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_decap_8 FILLER_22_183 ();
 sg13g2_decap_8 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_197 ();
 sg13g2_decap_4 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_208 ();
 sg13g2_decap_4 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_decap_4 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_242 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_359 ();
 sg13g2_decap_4 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_58 ();
 sg13g2_decap_8 FILLER_23_65 ();
 sg13g2_decap_8 FILLER_23_72 ();
 sg13g2_decap_8 FILLER_23_79 ();
 sg13g2_decap_4 FILLER_23_86 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_152 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_8 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_223 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_decap_4 FILLER_23_330 ();
 sg13g2_fill_2 FILLER_23_342 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_decap_4 FILLER_23_350 ();
 sg13g2_decap_4 FILLER_23_358 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_416 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_decap_8 FILLER_24_55 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_decap_4 FILLER_24_94 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_decap_8 FILLER_24_111 ();
 sg13g2_decap_8 FILLER_24_139 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_decap_8 FILLER_24_180 ();
 sg13g2_decap_8 FILLER_24_187 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_323 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_374 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_4 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_decap_4 FILLER_25_85 ();
 sg13g2_decap_8 FILLER_25_93 ();
 sg13g2_decap_4 FILLER_25_100 ();
 sg13g2_decap_8 FILLER_25_108 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_decap_8 FILLER_25_176 ();
 sg13g2_decap_4 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_decap_4 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_decap_4 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_8 FILLER_25_404 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_50 ();
 sg13g2_decap_8 FILLER_26_57 ();
 sg13g2_decap_8 FILLER_26_64 ();
 sg13g2_fill_2 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_decap_8 FILLER_26_115 ();
 sg13g2_decap_8 FILLER_26_122 ();
 sg13g2_decap_8 FILLER_26_129 ();
 sg13g2_decap_8 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_150 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_4 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_decap_4 FILLER_26_346 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_fill_1 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_26_409 ();
 sg13g2_decap_8 FILLER_26_416 ();
 sg13g2_decap_8 FILLER_26_423 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_177 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_decap_4 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_decap_4 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_decap_4 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_27_412 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_decap_8 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_171 ();
 sg13g2_decap_4 FILLER_28_178 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_decap_4 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_4 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_205 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_4 FILLER_29_349 ();
 sg13g2_decap_4 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_4 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_4 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_decap_8 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_136 ();
 sg13g2_decap_4 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_204 ();
 sg13g2_decap_4 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_decap_4 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_decap_4 FILLER_30_354 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_4 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_8 FILLER_30_404 ();
 sg13g2_decap_8 FILLER_30_411 ();
 sg13g2_decap_8 FILLER_30_418 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_fill_2 FILLER_31_68 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_83 ();
 sg13g2_fill_2 FILLER_31_97 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_135 ();
 sg13g2_decap_4 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_153 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_decap_8 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_312 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_128 ();
 sg13g2_decap_4 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_176 ();
 sg13g2_decap_8 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_decap_4 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_255 ();
 sg13g2_decap_4 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_decap_4 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_decap_4 FILLER_32_366 ();
 sg13g2_decap_4 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_decap_4 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_57 ();
 sg13g2_decap_8 FILLER_33_64 ();
 sg13g2_decap_8 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_85 ();
 sg13g2_decap_4 FILLER_33_118 ();
 sg13g2_decap_4 FILLER_33_153 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_decap_4 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_decap_4 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_286 ();
 sg13g2_decap_8 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_314 ();
 sg13g2_decap_8 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_333 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_decap_4 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_decap_4 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_108 ();
 sg13g2_decap_8 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_decap_8 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_169 ();
 sg13g2_decap_4 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_259 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_decap_4 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_2 FILLER_34_319 ();
 sg13g2_decap_4 FILLER_34_327 ();
 sg13g2_fill_2 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_fill_2 FILLER_34_374 ();
 sg13g2_decap_4 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_decap_4 FILLER_34_426 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_fill_2 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_2 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_80 ();
 sg13g2_decap_4 FILLER_35_85 ();
 sg13g2_fill_1 FILLER_35_89 ();
 sg13g2_fill_1 FILLER_35_94 ();
 sg13g2_decap_8 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_106 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_decap_4 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_261 ();
 sg13g2_decap_4 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_decap_4 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_decap_8 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_37 ();
 sg13g2_fill_1 FILLER_36_68 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_181 ();
 sg13g2_decap_8 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_257 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_decap_4 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_36_412 ();
 sg13g2_decap_8 FILLER_36_419 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_25 ();
 sg13g2_decap_8 FILLER_37_52 ();
 sg13g2_decap_4 FILLER_37_59 ();
 sg13g2_fill_2 FILLER_37_83 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_fill_1 FILLER_37_111 ();
 sg13g2_decap_8 FILLER_37_120 ();
 sg13g2_decap_4 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_285 ();
 sg13g2_decap_4 FILLER_37_292 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_4 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_2 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_362 ();
 sg13g2_decap_4 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_8 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_decap_8 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_40 ();
 sg13g2_decap_8 FILLER_38_47 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_decap_4 FILLER_38_73 ();
 sg13g2_fill_1 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_decap_4 FILLER_38_109 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_decap_4 FILLER_38_118 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_decap_4 FILLER_38_128 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_decap_8 FILLER_38_150 ();
 sg13g2_decap_8 FILLER_38_157 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_4 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_decap_4 FILLER_38_260 ();
 sg13g2_decap_4 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_decap_4 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_decap_4 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_53 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_decap_4 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_71 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_fill_2 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_94 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_decap_8 FILLER_39_143 ();
 sg13g2_decap_8 FILLER_39_150 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_fill_2 FILLER_39_166 ();
 sg13g2_fill_1 FILLER_39_176 ();
 sg13g2_fill_1 FILLER_39_181 ();
 sg13g2_decap_8 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_193 ();
 sg13g2_decap_4 FILLER_39_200 ();
 sg13g2_decap_8 FILLER_39_208 ();
 sg13g2_decap_4 FILLER_39_215 ();
 sg13g2_fill_2 FILLER_39_219 ();
 sg13g2_decap_4 FILLER_39_225 ();
 sg13g2_fill_1 FILLER_39_229 ();
 sg13g2_decap_8 FILLER_39_239 ();
 sg13g2_fill_2 FILLER_39_246 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_fill_2 FILLER_39_259 ();
 sg13g2_decap_4 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_278 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_fill_2 FILLER_39_314 ();
 sg13g2_decap_4 FILLER_39_329 ();
 sg13g2_fill_2 FILLER_39_338 ();
 sg13g2_decap_4 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_353 ();
 sg13g2_fill_2 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_380 ();
 sg13g2_fill_2 FILLER_39_398 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_fill_2 FILLER_39_427 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_79 ();
 sg13g2_decap_4 FILLER_40_86 ();
 sg13g2_decap_8 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_4 FILLER_40_109 ();
 sg13g2_fill_2 FILLER_40_113 ();
 sg13g2_fill_2 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_4 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_226 ();
 sg13g2_decap_4 FILLER_40_235 ();
 sg13g2_decap_8 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_261 ();
 sg13g2_decap_8 FILLER_40_268 ();
 sg13g2_decap_4 FILLER_40_275 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_decap_8 FILLER_40_288 ();
 sg13g2_decap_4 FILLER_40_295 ();
 sg13g2_fill_2 FILLER_40_299 ();
 sg13g2_decap_4 FILLER_40_307 ();
 sg13g2_fill_1 FILLER_40_311 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_fill_2 FILLER_40_331 ();
 sg13g2_decap_8 FILLER_40_338 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_387 ();
 sg13g2_decap_4 FILLER_40_400 ();
 sg13g2_decap_8 FILLER_40_409 ();
 sg13g2_decap_8 FILLER_40_416 ();
 sg13g2_decap_8 FILLER_40_423 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_4 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_51 ();
 sg13g2_decap_8 FILLER_41_62 ();
 sg13g2_decap_4 FILLER_41_69 ();
 sg13g2_decap_4 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_102 ();
 sg13g2_decap_8 FILLER_41_128 ();
 sg13g2_decap_4 FILLER_41_135 ();
 sg13g2_fill_2 FILLER_41_139 ();
 sg13g2_decap_8 FILLER_41_146 ();
 sg13g2_decap_8 FILLER_41_153 ();
 sg13g2_decap_8 FILLER_41_160 ();
 sg13g2_decap_4 FILLER_41_167 ();
 sg13g2_fill_2 FILLER_41_171 ();
 sg13g2_decap_8 FILLER_41_177 ();
 sg13g2_decap_8 FILLER_41_184 ();
 sg13g2_decap_8 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_decap_8 FILLER_41_204 ();
 sg13g2_decap_4 FILLER_41_211 ();
 sg13g2_fill_1 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_234 ();
 sg13g2_fill_2 FILLER_41_241 ();
 sg13g2_fill_2 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_decap_8 FILLER_41_263 ();
 sg13g2_decap_4 FILLER_41_270 ();
 sg13g2_fill_1 FILLER_41_279 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_decap_4 FILLER_41_291 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_302 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_328 ();
 sg13g2_decap_4 FILLER_41_335 ();
 sg13g2_fill_2 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_fill_2 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_363 ();
 sg13g2_fill_1 FILLER_41_370 ();
 sg13g2_decap_8 FILLER_41_375 ();
 sg13g2_fill_1 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_decap_8 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_41_415 ();
 sg13g2_decap_8 FILLER_41_422 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_fill_1 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_48 ();
 sg13g2_fill_1 FILLER_42_50 ();
 sg13g2_decap_8 FILLER_42_59 ();
 sg13g2_decap_8 FILLER_42_66 ();
 sg13g2_fill_2 FILLER_42_73 ();
 sg13g2_decap_8 FILLER_42_79 ();
 sg13g2_fill_1 FILLER_42_91 ();
 sg13g2_fill_1 FILLER_42_102 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_decap_4 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_decap_8 FILLER_42_128 ();
 sg13g2_decap_4 FILLER_42_135 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_165 ();
 sg13g2_decap_8 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_179 ();
 sg13g2_decap_8 FILLER_42_186 ();
 sg13g2_decap_8 FILLER_42_193 ();
 sg13g2_decap_8 FILLER_42_200 ();
 sg13g2_decap_8 FILLER_42_207 ();
 sg13g2_decap_8 FILLER_42_214 ();
 sg13g2_decap_8 FILLER_42_221 ();
 sg13g2_decap_4 FILLER_42_228 ();
 sg13g2_fill_1 FILLER_42_232 ();
 sg13g2_decap_4 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_250 ();
 sg13g2_fill_1 FILLER_42_257 ();
 sg13g2_fill_1 FILLER_42_265 ();
 sg13g2_fill_1 FILLER_42_307 ();
 sg13g2_decap_8 FILLER_42_319 ();
 sg13g2_decap_8 FILLER_42_326 ();
 sg13g2_decap_4 FILLER_42_333 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_342 ();
 sg13g2_decap_8 FILLER_42_353 ();
 sg13g2_fill_1 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_386 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_419 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_37 ();
 sg13g2_decap_4 FILLER_43_44 ();
 sg13g2_decap_8 FILLER_43_52 ();
 sg13g2_decap_8 FILLER_43_59 ();
 sg13g2_decap_8 FILLER_43_66 ();
 sg13g2_decap_8 FILLER_43_73 ();
 sg13g2_decap_8 FILLER_43_80 ();
 sg13g2_fill_2 FILLER_43_87 ();
 sg13g2_fill_1 FILLER_43_89 ();
 sg13g2_fill_2 FILLER_43_102 ();
 sg13g2_fill_2 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_130 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_decap_8 FILLER_43_170 ();
 sg13g2_decap_8 FILLER_43_177 ();
 sg13g2_decap_8 FILLER_43_184 ();
 sg13g2_decap_8 FILLER_43_191 ();
 sg13g2_decap_8 FILLER_43_198 ();
 sg13g2_decap_8 FILLER_43_209 ();
 sg13g2_decap_8 FILLER_43_216 ();
 sg13g2_decap_4 FILLER_43_223 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_decap_8 FILLER_43_233 ();
 sg13g2_decap_8 FILLER_43_240 ();
 sg13g2_fill_1 FILLER_43_247 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_4 FILLER_43_268 ();
 sg13g2_fill_1 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_279 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_300 ();
 sg13g2_decap_8 FILLER_43_309 ();
 sg13g2_decap_8 FILLER_43_316 ();
 sg13g2_decap_8 FILLER_43_323 ();
 sg13g2_decap_8 FILLER_43_330 ();
 sg13g2_fill_2 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_339 ();
 sg13g2_decap_4 FILLER_43_345 ();
 sg13g2_fill_2 FILLER_43_349 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_4 FILLER_43_378 ();
 sg13g2_fill_2 FILLER_43_386 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_fill_2 FILLER_43_427 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_78 ();
 sg13g2_fill_1 FILLER_44_80 ();
 sg13g2_fill_2 FILLER_44_86 ();
 sg13g2_fill_1 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_106 ();
 sg13g2_decap_8 FILLER_44_113 ();
 sg13g2_decap_8 FILLER_44_120 ();
 sg13g2_decap_8 FILLER_44_127 ();
 sg13g2_decap_8 FILLER_44_134 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_159 ();
 sg13g2_decap_8 FILLER_44_170 ();
 sg13g2_decap_8 FILLER_44_177 ();
 sg13g2_decap_8 FILLER_44_184 ();
 sg13g2_decap_8 FILLER_44_191 ();
 sg13g2_decap_4 FILLER_44_198 ();
 sg13g2_decap_4 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_231 ();
 sg13g2_decap_4 FILLER_44_245 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_257 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_fill_2 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_fill_1 FILLER_44_290 ();
 sg13g2_fill_2 FILLER_44_295 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_321 ();
 sg13g2_fill_2 FILLER_44_328 ();
 sg13g2_decap_8 FILLER_44_335 ();
 sg13g2_decap_4 FILLER_44_342 ();
 sg13g2_fill_1 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_356 ();
 sg13g2_decap_4 FILLER_44_362 ();
 sg13g2_fill_1 FILLER_44_380 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_4 FILLER_44_424 ();
 sg13g2_fill_2 FILLER_44_428 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_64 ();
 sg13g2_fill_1 FILLER_45_66 ();
 sg13g2_decap_4 FILLER_45_85 ();
 sg13g2_fill_1 FILLER_45_89 ();
 sg13g2_fill_2 FILLER_45_99 ();
 sg13g2_decap_8 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_113 ();
 sg13g2_decap_8 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_decap_8 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_164 ();
 sg13g2_decap_8 FILLER_45_171 ();
 sg13g2_decap_8 FILLER_45_178 ();
 sg13g2_decap_8 FILLER_45_195 ();
 sg13g2_decap_8 FILLER_45_202 ();
 sg13g2_decap_8 FILLER_45_209 ();
 sg13g2_decap_4 FILLER_45_216 ();
 sg13g2_fill_1 FILLER_45_220 ();
 sg13g2_decap_4 FILLER_45_253 ();
 sg13g2_fill_1 FILLER_45_262 ();
 sg13g2_decap_8 FILLER_45_267 ();
 sg13g2_fill_1 FILLER_45_274 ();
 sg13g2_decap_8 FILLER_45_286 ();
 sg13g2_fill_1 FILLER_45_293 ();
 sg13g2_decap_4 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_4 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_353 ();
 sg13g2_fill_2 FILLER_45_359 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_fill_2 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_375 ();
 sg13g2_fill_2 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_45_393 ();
 sg13g2_decap_8 FILLER_45_400 ();
 sg13g2_decap_8 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_45_414 ();
 sg13g2_decap_8 FILLER_45_421 ();
 sg13g2_fill_2 FILLER_45_428 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_4 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_25 ();
 sg13g2_decap_8 FILLER_46_30 ();
 sg13g2_decap_8 FILLER_46_37 ();
 sg13g2_decap_8 FILLER_46_44 ();
 sg13g2_decap_8 FILLER_46_51 ();
 sg13g2_decap_8 FILLER_46_58 ();
 sg13g2_decap_4 FILLER_46_65 ();
 sg13g2_decap_4 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_decap_8 FILLER_46_99 ();
 sg13g2_decap_8 FILLER_46_106 ();
 sg13g2_decap_8 FILLER_46_113 ();
 sg13g2_decap_8 FILLER_46_120 ();
 sg13g2_decap_8 FILLER_46_127 ();
 sg13g2_decap_8 FILLER_46_134 ();
 sg13g2_decap_8 FILLER_46_141 ();
 sg13g2_decap_8 FILLER_46_148 ();
 sg13g2_decap_4 FILLER_46_155 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_decap_8 FILLER_46_166 ();
 sg13g2_decap_8 FILLER_46_173 ();
 sg13g2_decap_8 FILLER_46_180 ();
 sg13g2_decap_8 FILLER_46_187 ();
 sg13g2_decap_8 FILLER_46_194 ();
 sg13g2_decap_8 FILLER_46_201 ();
 sg13g2_decap_8 FILLER_46_208 ();
 sg13g2_decap_8 FILLER_46_215 ();
 sg13g2_decap_4 FILLER_46_222 ();
 sg13g2_fill_2 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_246 ();
 sg13g2_fill_2 FILLER_46_255 ();
 sg13g2_fill_1 FILLER_46_257 ();
 sg13g2_fill_2 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_300 ();
 sg13g2_fill_2 FILLER_46_307 ();
 sg13g2_fill_2 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_321 ();
 sg13g2_fill_2 FILLER_46_327 ();
 sg13g2_fill_1 FILLER_46_329 ();
 sg13g2_fill_2 FILLER_46_336 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_344 ();
 sg13g2_fill_1 FILLER_46_357 ();
 sg13g2_fill_2 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_decap_8 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_46_415 ();
 sg13g2_decap_8 FILLER_46_422 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_58 ();
 sg13g2_decap_8 FILLER_47_65 ();
 sg13g2_decap_8 FILLER_47_72 ();
 sg13g2_decap_4 FILLER_47_79 ();
 sg13g2_fill_1 FILLER_47_97 ();
 sg13g2_decap_8 FILLER_47_106 ();
 sg13g2_decap_8 FILLER_47_113 ();
 sg13g2_decap_8 FILLER_47_120 ();
 sg13g2_fill_1 FILLER_47_127 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_135 ();
 sg13g2_decap_4 FILLER_47_141 ();
 sg13g2_fill_1 FILLER_47_145 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_4 FILLER_47_175 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_decap_8 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_195 ();
 sg13g2_decap_4 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_206 ();
 sg13g2_decap_8 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_219 ();
 sg13g2_fill_1 FILLER_47_226 ();
 sg13g2_decap_8 FILLER_47_239 ();
 sg13g2_decap_4 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_250 ();
 sg13g2_fill_2 FILLER_47_264 ();
 sg13g2_decap_8 FILLER_47_276 ();
 sg13g2_decap_4 FILLER_47_283 ();
 sg13g2_decap_8 FILLER_47_305 ();
 sg13g2_decap_8 FILLER_47_312 ();
 sg13g2_decap_8 FILLER_47_319 ();
 sg13g2_decap_8 FILLER_47_326 ();
 sg13g2_fill_2 FILLER_47_333 ();
 sg13g2_fill_1 FILLER_47_335 ();
 sg13g2_decap_4 FILLER_47_353 ();
 sg13g2_fill_1 FILLER_47_357 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_decap_4 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_fill_1 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_403 ();
 sg13g2_decap_8 FILLER_47_410 ();
 sg13g2_decap_8 FILLER_47_417 ();
 sg13g2_decap_4 FILLER_47_424 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_decap_8 FILLER_48_12 ();
 sg13g2_fill_1 FILLER_48_19 ();
 sg13g2_decap_4 FILLER_48_26 ();
 sg13g2_fill_1 FILLER_48_30 ();
 sg13g2_decap_4 FILLER_48_37 ();
 sg13g2_decap_8 FILLER_48_71 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_decap_8 FILLER_48_99 ();
 sg13g2_decap_4 FILLER_48_106 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_fill_2 FILLER_48_137 ();
 sg13g2_decap_4 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_184 ();
 sg13g2_decap_8 FILLER_48_191 ();
 sg13g2_decap_8 FILLER_48_198 ();
 sg13g2_decap_8 FILLER_48_205 ();
 sg13g2_decap_8 FILLER_48_212 ();
 sg13g2_decap_8 FILLER_48_219 ();
 sg13g2_decap_4 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_234 ();
 sg13g2_fill_2 FILLER_48_242 ();
 sg13g2_fill_1 FILLER_48_244 ();
 sg13g2_decap_8 FILLER_48_254 ();
 sg13g2_decap_8 FILLER_48_261 ();
 sg13g2_decap_8 FILLER_48_268 ();
 sg13g2_decap_8 FILLER_48_275 ();
 sg13g2_decap_8 FILLER_48_282 ();
 sg13g2_decap_4 FILLER_48_289 ();
 sg13g2_fill_2 FILLER_48_293 ();
 sg13g2_decap_8 FILLER_48_300 ();
 sg13g2_fill_2 FILLER_48_307 ();
 sg13g2_decap_8 FILLER_48_314 ();
 sg13g2_decap_4 FILLER_48_321 ();
 sg13g2_fill_2 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_decap_4 FILLER_48_350 ();
 sg13g2_fill_1 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_360 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_8 FILLER_48_404 ();
 sg13g2_decap_8 FILLER_48_411 ();
 sg13g2_decap_8 FILLER_48_418 ();
 sg13g2_decap_4 FILLER_48_425 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_14 ();
 sg13g2_decap_4 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_37 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_52 ();
 sg13g2_decap_8 FILLER_49_57 ();
 sg13g2_decap_8 FILLER_49_64 ();
 sg13g2_decap_4 FILLER_49_71 ();
 sg13g2_fill_1 FILLER_49_75 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_4 FILLER_49_168 ();
 sg13g2_fill_2 FILLER_49_172 ();
 sg13g2_decap_4 FILLER_49_183 ();
 sg13g2_fill_2 FILLER_49_187 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_1 FILLER_49_230 ();
 sg13g2_fill_2 FILLER_49_235 ();
 sg13g2_fill_1 FILLER_49_237 ();
 sg13g2_fill_2 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_262 ();
 sg13g2_decap_4 FILLER_49_269 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_290 ();
 sg13g2_decap_8 FILLER_49_297 ();
 sg13g2_decap_4 FILLER_49_304 ();
 sg13g2_fill_1 FILLER_49_308 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_2 FILLER_49_339 ();
 sg13g2_fill_2 FILLER_49_350 ();
 sg13g2_fill_1 FILLER_49_352 ();
 sg13g2_decap_4 FILLER_49_367 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_decap_4 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_4 FILLER_49_424 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_4 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_69 ();
 sg13g2_decap_8 FILLER_50_76 ();
 sg13g2_fill_2 FILLER_50_83 ();
 sg13g2_decap_4 FILLER_50_102 ();
 sg13g2_fill_1 FILLER_50_106 ();
 sg13g2_fill_2 FILLER_50_111 ();
 sg13g2_decap_8 FILLER_50_118 ();
 sg13g2_decap_8 FILLER_50_125 ();
 sg13g2_decap_8 FILLER_50_132 ();
 sg13g2_decap_8 FILLER_50_139 ();
 sg13g2_decap_8 FILLER_50_146 ();
 sg13g2_decap_8 FILLER_50_153 ();
 sg13g2_decap_8 FILLER_50_160 ();
 sg13g2_decap_4 FILLER_50_167 ();
 sg13g2_fill_2 FILLER_50_171 ();
 sg13g2_decap_8 FILLER_50_186 ();
 sg13g2_decap_8 FILLER_50_193 ();
 sg13g2_decap_8 FILLER_50_200 ();
 sg13g2_decap_8 FILLER_50_207 ();
 sg13g2_decap_8 FILLER_50_214 ();
 sg13g2_decap_4 FILLER_50_221 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_fill_2 FILLER_50_240 ();
 sg13g2_fill_1 FILLER_50_242 ();
 sg13g2_fill_1 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_284 ();
 sg13g2_decap_4 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_decap_8 FILLER_50_316 ();
 sg13g2_fill_2 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_325 ();
 sg13g2_decap_8 FILLER_50_335 ();
 sg13g2_fill_2 FILLER_50_342 ();
 sg13g2_fill_1 FILLER_50_344 ();
 sg13g2_fill_2 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_367 ();
 sg13g2_fill_1 FILLER_50_374 ();
 sg13g2_fill_2 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_8 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_50_412 ();
 sg13g2_decap_8 FILLER_50_419 ();
 sg13g2_decap_4 FILLER_50_426 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_fill_1 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_68 ();
 sg13g2_decap_8 FILLER_51_75 ();
 sg13g2_decap_8 FILLER_51_82 ();
 sg13g2_decap_4 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_fill_2 FILLER_51_136 ();
 sg13g2_decap_8 FILLER_51_145 ();
 sg13g2_decap_8 FILLER_51_152 ();
 sg13g2_decap_8 FILLER_51_163 ();
 sg13g2_decap_8 FILLER_51_170 ();
 sg13g2_fill_2 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_179 ();
 sg13g2_fill_2 FILLER_51_184 ();
 sg13g2_decap_8 FILLER_51_191 ();
 sg13g2_decap_8 FILLER_51_198 ();
 sg13g2_decap_8 FILLER_51_205 ();
 sg13g2_decap_8 FILLER_51_212 ();
 sg13g2_fill_1 FILLER_51_228 ();
 sg13g2_fill_1 FILLER_51_234 ();
 sg13g2_decap_8 FILLER_51_244 ();
 sg13g2_fill_2 FILLER_51_275 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_decap_8 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_298 ();
 sg13g2_fill_1 FILLER_51_311 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_decap_8 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_331 ();
 sg13g2_fill_2 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_345 ();
 sg13g2_fill_1 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_51_353 ();
 sg13g2_fill_2 FILLER_51_360 ();
 sg13g2_fill_1 FILLER_51_362 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_384 ();
 sg13g2_decap_8 FILLER_51_395 ();
 sg13g2_decap_8 FILLER_51_402 ();
 sg13g2_decap_8 FILLER_51_409 ();
 sg13g2_decap_8 FILLER_51_416 ();
 sg13g2_decap_8 FILLER_51_423 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_50 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_83 ();
 sg13g2_decap_8 FILLER_52_90 ();
 sg13g2_decap_8 FILLER_52_97 ();
 sg13g2_decap_8 FILLER_52_108 ();
 sg13g2_decap_8 FILLER_52_115 ();
 sg13g2_decap_8 FILLER_52_122 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_decap_8 FILLER_52_160 ();
 sg13g2_fill_2 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_169 ();
 sg13g2_decap_8 FILLER_52_180 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_decap_8 FILLER_52_192 ();
 sg13g2_decap_8 FILLER_52_199 ();
 sg13g2_decap_8 FILLER_52_206 ();
 sg13g2_fill_2 FILLER_52_213 ();
 sg13g2_fill_1 FILLER_52_215 ();
 sg13g2_decap_4 FILLER_52_221 ();
 sg13g2_fill_2 FILLER_52_225 ();
 sg13g2_fill_1 FILLER_52_232 ();
 sg13g2_fill_1 FILLER_52_239 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_decap_8 FILLER_52_271 ();
 sg13g2_decap_4 FILLER_52_278 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_4 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_298 ();
 sg13g2_decap_4 FILLER_52_321 ();
 sg13g2_decap_4 FILLER_52_330 ();
 sg13g2_decap_4 FILLER_52_339 ();
 sg13g2_fill_2 FILLER_52_343 ();
 sg13g2_fill_1 FILLER_52_361 ();
 sg13g2_decap_4 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_fill_2 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_380 ();
 sg13g2_decap_8 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_52_415 ();
 sg13g2_decap_8 FILLER_52_422 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_40 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_4 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_81 ();
 sg13g2_fill_2 FILLER_53_86 ();
 sg13g2_decap_8 FILLER_53_92 ();
 sg13g2_decap_8 FILLER_53_99 ();
 sg13g2_decap_4 FILLER_53_106 ();
 sg13g2_fill_2 FILLER_53_110 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_145 ();
 sg13g2_decap_8 FILLER_53_152 ();
 sg13g2_decap_4 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_163 ();
 sg13g2_decap_8 FILLER_53_184 ();
 sg13g2_decap_8 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_198 ();
 sg13g2_decap_8 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_212 ();
 sg13g2_decap_8 FILLER_53_219 ();
 sg13g2_decap_4 FILLER_53_226 ();
 sg13g2_fill_1 FILLER_53_230 ();
 sg13g2_decap_4 FILLER_53_246 ();
 sg13g2_fill_2 FILLER_53_254 ();
 sg13g2_decap_8 FILLER_53_260 ();
 sg13g2_decap_8 FILLER_53_267 ();
 sg13g2_decap_4 FILLER_53_274 ();
 sg13g2_fill_1 FILLER_53_278 ();
 sg13g2_decap_8 FILLER_53_283 ();
 sg13g2_decap_8 FILLER_53_296 ();
 sg13g2_decap_8 FILLER_53_303 ();
 sg13g2_decap_8 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_317 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_decap_8 FILLER_53_330 ();
 sg13g2_decap_8 FILLER_53_337 ();
 sg13g2_decap_4 FILLER_53_344 ();
 sg13g2_fill_1 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_365 ();
 sg13g2_fill_2 FILLER_53_372 ();
 sg13g2_fill_1 FILLER_53_374 ();
 sg13g2_fill_1 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_decap_8 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_53_415 ();
 sg13g2_decap_8 FILLER_53_422 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_40 ();
 sg13g2_decap_8 FILLER_54_47 ();
 sg13g2_decap_8 FILLER_54_54 ();
 sg13g2_fill_1 FILLER_54_61 ();
 sg13g2_decap_8 FILLER_54_66 ();
 sg13g2_decap_8 FILLER_54_73 ();
 sg13g2_decap_4 FILLER_54_80 ();
 sg13g2_fill_1 FILLER_54_84 ();
 sg13g2_fill_1 FILLER_54_97 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_4 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_180 ();
 sg13g2_decap_8 FILLER_54_187 ();
 sg13g2_decap_8 FILLER_54_194 ();
 sg13g2_decap_8 FILLER_54_201 ();
 sg13g2_decap_8 FILLER_54_208 ();
 sg13g2_decap_4 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_219 ();
 sg13g2_fill_1 FILLER_54_229 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_246 ();
 sg13g2_fill_1 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_267 ();
 sg13g2_decap_4 FILLER_54_272 ();
 sg13g2_fill_1 FILLER_54_276 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_fill_2 FILLER_54_304 ();
 sg13g2_fill_1 FILLER_54_306 ();
 sg13g2_decap_4 FILLER_54_317 ();
 sg13g2_fill_1 FILLER_54_321 ();
 sg13g2_decap_8 FILLER_54_326 ();
 sg13g2_fill_2 FILLER_54_333 ();
 sg13g2_decap_8 FILLER_54_339 ();
 sg13g2_fill_2 FILLER_54_346 ();
 sg13g2_fill_1 FILLER_54_348 ();
 sg13g2_decap_4 FILLER_54_354 ();
 sg13g2_fill_1 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_363 ();
 sg13g2_decap_8 FILLER_54_370 ();
 sg13g2_fill_2 FILLER_54_382 ();
 sg13g2_decap_8 FILLER_54_388 ();
 sg13g2_decap_8 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_decap_8 FILLER_54_409 ();
 sg13g2_decap_8 FILLER_54_416 ();
 sg13g2_decap_8 FILLER_54_423 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_20 ();
 sg13g2_decap_4 FILLER_55_27 ();
 sg13g2_fill_1 FILLER_55_39 ();
 sg13g2_fill_2 FILLER_55_45 ();
 sg13g2_fill_2 FILLER_55_51 ();
 sg13g2_fill_1 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_92 ();
 sg13g2_decap_4 FILLER_55_113 ();
 sg13g2_decap_8 FILLER_55_125 ();
 sg13g2_fill_2 FILLER_55_132 ();
 sg13g2_decap_8 FILLER_55_159 ();
 sg13g2_decap_4 FILLER_55_166 ();
 sg13g2_decap_8 FILLER_55_178 ();
 sg13g2_decap_8 FILLER_55_195 ();
 sg13g2_decap_8 FILLER_55_202 ();
 sg13g2_decap_8 FILLER_55_209 ();
 sg13g2_decap_8 FILLER_55_216 ();
 sg13g2_decap_4 FILLER_55_223 ();
 sg13g2_decap_4 FILLER_55_238 ();
 sg13g2_fill_2 FILLER_55_242 ();
 sg13g2_decap_4 FILLER_55_262 ();
 sg13g2_fill_1 FILLER_55_266 ();
 sg13g2_fill_2 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_fill_2 FILLER_55_337 ();
 sg13g2_decap_4 FILLER_55_348 ();
 sg13g2_decap_4 FILLER_55_367 ();
 sg13g2_fill_2 FILLER_55_385 ();
 sg13g2_fill_1 FILLER_55_387 ();
 sg13g2_fill_2 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_398 ();
 sg13g2_decap_8 FILLER_55_405 ();
 sg13g2_decap_8 FILLER_55_412 ();
 sg13g2_decap_8 FILLER_55_419 ();
 sg13g2_decap_4 FILLER_55_426 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_4 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_32 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_decap_8 FILLER_56_54 ();
 sg13g2_decap_8 FILLER_56_61 ();
 sg13g2_decap_8 FILLER_56_68 ();
 sg13g2_decap_8 FILLER_56_75 ();
 sg13g2_decap_8 FILLER_56_82 ();
 sg13g2_decap_8 FILLER_56_89 ();
 sg13g2_decap_8 FILLER_56_96 ();
 sg13g2_fill_2 FILLER_56_103 ();
 sg13g2_fill_1 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_110 ();
 sg13g2_decap_8 FILLER_56_117 ();
 sg13g2_fill_2 FILLER_56_124 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_142 ();
 sg13g2_decap_8 FILLER_56_149 ();
 sg13g2_decap_8 FILLER_56_156 ();
 sg13g2_decap_8 FILLER_56_163 ();
 sg13g2_decap_8 FILLER_56_170 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_decap_8 FILLER_56_184 ();
 sg13g2_decap_8 FILLER_56_191 ();
 sg13g2_decap_8 FILLER_56_198 ();
 sg13g2_decap_8 FILLER_56_205 ();
 sg13g2_decap_4 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_216 ();
 sg13g2_decap_8 FILLER_56_221 ();
 sg13g2_fill_1 FILLER_56_233 ();
 sg13g2_decap_8 FILLER_56_241 ();
 sg13g2_fill_2 FILLER_56_248 ();
 sg13g2_fill_1 FILLER_56_260 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_decap_8 FILLER_56_298 ();
 sg13g2_decap_8 FILLER_56_305 ();
 sg13g2_fill_2 FILLER_56_312 ();
 sg13g2_decap_8 FILLER_56_324 ();
 sg13g2_fill_1 FILLER_56_331 ();
 sg13g2_fill_1 FILLER_56_336 ();
 sg13g2_fill_2 FILLER_56_342 ();
 sg13g2_fill_1 FILLER_56_363 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_56_412 ();
 sg13g2_decap_8 FILLER_56_419 ();
 sg13g2_decap_4 FILLER_56_426 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_decap_8 FILLER_57_55 ();
 sg13g2_decap_8 FILLER_57_62 ();
 sg13g2_decap_8 FILLER_57_69 ();
 sg13g2_decap_8 FILLER_57_76 ();
 sg13g2_decap_8 FILLER_57_83 ();
 sg13g2_decap_8 FILLER_57_90 ();
 sg13g2_decap_8 FILLER_57_97 ();
 sg13g2_decap_8 FILLER_57_104 ();
 sg13g2_decap_8 FILLER_57_111 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_4 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_180 ();
 sg13g2_decap_8 FILLER_57_187 ();
 sg13g2_decap_8 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_201 ();
 sg13g2_decap_8 FILLER_57_208 ();
 sg13g2_decap_4 FILLER_57_215 ();
 sg13g2_fill_2 FILLER_57_219 ();
 sg13g2_fill_1 FILLER_57_226 ();
 sg13g2_decap_4 FILLER_57_239 ();
 sg13g2_decap_4 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_258 ();
 sg13g2_decap_8 FILLER_57_265 ();
 sg13g2_decap_8 FILLER_57_272 ();
 sg13g2_decap_8 FILLER_57_279 ();
 sg13g2_decap_4 FILLER_57_286 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_decap_8 FILLER_57_296 ();
 sg13g2_decap_8 FILLER_57_303 ();
 sg13g2_decap_4 FILLER_57_310 ();
 sg13g2_decap_4 FILLER_57_320 ();
 sg13g2_fill_2 FILLER_57_324 ();
 sg13g2_decap_8 FILLER_57_330 ();
 sg13g2_decap_8 FILLER_57_337 ();
 sg13g2_decap_8 FILLER_57_344 ();
 sg13g2_fill_2 FILLER_57_351 ();
 sg13g2_decap_8 FILLER_57_358 ();
 sg13g2_fill_1 FILLER_57_365 ();
 sg13g2_decap_4 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_fill_2 FILLER_57_386 ();
 sg13g2_fill_1 FILLER_57_396 ();
 sg13g2_decap_8 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_57_412 ();
 sg13g2_decap_8 FILLER_57_419 ();
 sg13g2_decap_4 FILLER_57_426 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_11 ();
 sg13g2_decap_8 FILLER_58_18 ();
 sg13g2_decap_4 FILLER_58_25 ();
 sg13g2_fill_1 FILLER_58_29 ();
 sg13g2_decap_8 FILLER_58_39 ();
 sg13g2_fill_2 FILLER_58_46 ();
 sg13g2_fill_2 FILLER_58_53 ();
 sg13g2_fill_1 FILLER_58_55 ();
 sg13g2_decap_8 FILLER_58_87 ();
 sg13g2_decap_8 FILLER_58_94 ();
 sg13g2_decap_8 FILLER_58_101 ();
 sg13g2_decap_8 FILLER_58_108 ();
 sg13g2_fill_1 FILLER_58_115 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_122 ();
 sg13g2_fill_2 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_145 ();
 sg13g2_decap_8 FILLER_58_152 ();
 sg13g2_decap_8 FILLER_58_159 ();
 sg13g2_decap_8 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_58_173 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_fill_1 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_198 ();
 sg13g2_decap_8 FILLER_58_205 ();
 sg13g2_fill_2 FILLER_58_212 ();
 sg13g2_decap_4 FILLER_58_219 ();
 sg13g2_decap_4 FILLER_58_237 ();
 sg13g2_decap_4 FILLER_58_258 ();
 sg13g2_decap_8 FILLER_58_276 ();
 sg13g2_decap_4 FILLER_58_283 ();
 sg13g2_fill_1 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_305 ();
 sg13g2_fill_2 FILLER_58_311 ();
 sg13g2_decap_8 FILLER_58_317 ();
 sg13g2_decap_8 FILLER_58_324 ();
 sg13g2_decap_4 FILLER_58_331 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_decap_4 FILLER_58_341 ();
 sg13g2_fill_2 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_359 ();
 sg13g2_fill_1 FILLER_58_361 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_decap_4 FILLER_58_376 ();
 sg13g2_decap_8 FILLER_58_390 ();
 sg13g2_decap_8 FILLER_58_397 ();
 sg13g2_decap_8 FILLER_58_404 ();
 sg13g2_decap_8 FILLER_58_411 ();
 sg13g2_decap_8 FILLER_58_418 ();
 sg13g2_decap_4 FILLER_58_425 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_1 FILLER_59_31 ();
 sg13g2_decap_8 FILLER_59_41 ();
 sg13g2_fill_1 FILLER_59_48 ();
 sg13g2_decap_4 FILLER_59_59 ();
 sg13g2_decap_8 FILLER_59_67 ();
 sg13g2_decap_4 FILLER_59_74 ();
 sg13g2_fill_1 FILLER_59_78 ();
 sg13g2_fill_1 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_115 ();
 sg13g2_fill_1 FILLER_59_120 ();
 sg13g2_fill_2 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_fill_2 FILLER_59_137 ();
 sg13g2_decap_8 FILLER_59_155 ();
 sg13g2_decap_8 FILLER_59_162 ();
 sg13g2_fill_2 FILLER_59_169 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_fill_1 FILLER_59_176 ();
 sg13g2_fill_2 FILLER_59_186 ();
 sg13g2_fill_1 FILLER_59_188 ();
 sg13g2_decap_8 FILLER_59_197 ();
 sg13g2_decap_8 FILLER_59_204 ();
 sg13g2_fill_1 FILLER_59_211 ();
 sg13g2_decap_4 FILLER_59_217 ();
 sg13g2_fill_2 FILLER_59_221 ();
 sg13g2_fill_1 FILLER_59_238 ();
 sg13g2_decap_4 FILLER_59_244 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_fill_1 FILLER_59_266 ();
 sg13g2_fill_1 FILLER_59_273 ();
 sg13g2_fill_2 FILLER_59_279 ();
 sg13g2_decap_8 FILLER_59_291 ();
 sg13g2_decap_4 FILLER_59_298 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_324 ();
 sg13g2_decap_8 FILLER_59_330 ();
 sg13g2_decap_4 FILLER_59_337 ();
 sg13g2_fill_2 FILLER_59_341 ();
 sg13g2_fill_2 FILLER_59_370 ();
 sg13g2_decap_8 FILLER_59_376 ();
 sg13g2_decap_8 FILLER_59_383 ();
 sg13g2_fill_2 FILLER_59_390 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_fill_2 FILLER_59_427 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_18 ();
 sg13g2_fill_1 FILLER_60_29 ();
 sg13g2_decap_8 FILLER_60_34 ();
 sg13g2_decap_4 FILLER_60_41 ();
 sg13g2_fill_2 FILLER_60_45 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_fill_2 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_79 ();
 sg13g2_fill_1 FILLER_60_116 ();
 sg13g2_decap_8 FILLER_60_121 ();
 sg13g2_decap_8 FILLER_60_128 ();
 sg13g2_fill_2 FILLER_60_135 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_decap_8 FILLER_60_157 ();
 sg13g2_decap_8 FILLER_60_169 ();
 sg13g2_decap_4 FILLER_60_176 ();
 sg13g2_decap_8 FILLER_60_188 ();
 sg13g2_decap_8 FILLER_60_195 ();
 sg13g2_decap_8 FILLER_60_202 ();
 sg13g2_decap_8 FILLER_60_209 ();
 sg13g2_decap_8 FILLER_60_216 ();
 sg13g2_decap_4 FILLER_60_223 ();
 sg13g2_fill_2 FILLER_60_227 ();
 sg13g2_decap_8 FILLER_60_237 ();
 sg13g2_decap_8 FILLER_60_244 ();
 sg13g2_decap_4 FILLER_60_267 ();
 sg13g2_fill_2 FILLER_60_271 ();
 sg13g2_decap_8 FILLER_60_288 ();
 sg13g2_decap_8 FILLER_60_295 ();
 sg13g2_decap_8 FILLER_60_302 ();
 sg13g2_fill_1 FILLER_60_309 ();
 sg13g2_decap_4 FILLER_60_315 ();
 sg13g2_fill_1 FILLER_60_319 ();
 sg13g2_fill_1 FILLER_60_334 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_2 FILLER_60_348 ();
 sg13g2_decap_4 FILLER_60_382 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_decap_8 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_60_414 ();
 sg13g2_decap_8 FILLER_60_421 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_fill_1 FILLER_61_21 ();
 sg13g2_decap_4 FILLER_61_27 ();
 sg13g2_decap_8 FILLER_61_45 ();
 sg13g2_fill_2 FILLER_61_52 ();
 sg13g2_decap_4 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_69 ();
 sg13g2_decap_8 FILLER_61_76 ();
 sg13g2_fill_2 FILLER_61_83 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_101 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_decap_4 FILLER_61_127 ();
 sg13g2_fill_2 FILLER_61_131 ();
 sg13g2_decap_4 FILLER_61_142 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_decap_8 FILLER_61_153 ();
 sg13g2_decap_8 FILLER_61_160 ();
 sg13g2_decap_8 FILLER_61_167 ();
 sg13g2_decap_8 FILLER_61_174 ();
 sg13g2_decap_8 FILLER_61_181 ();
 sg13g2_decap_8 FILLER_61_188 ();
 sg13g2_decap_8 FILLER_61_195 ();
 sg13g2_decap_8 FILLER_61_202 ();
 sg13g2_decap_8 FILLER_61_209 ();
 sg13g2_decap_8 FILLER_61_216 ();
 sg13g2_decap_8 FILLER_61_223 ();
 sg13g2_decap_8 FILLER_61_230 ();
 sg13g2_decap_8 FILLER_61_237 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_259 ();
 sg13g2_decap_4 FILLER_61_264 ();
 sg13g2_fill_1 FILLER_61_268 ();
 sg13g2_decap_8 FILLER_61_284 ();
 sg13g2_decap_8 FILLER_61_291 ();
 sg13g2_decap_8 FILLER_61_298 ();
 sg13g2_decap_4 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_decap_8 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_decap_8 FILLER_61_355 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_fill_2 FILLER_61_383 ();
 sg13g2_decap_4 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_61_403 ();
 sg13g2_decap_8 FILLER_61_410 ();
 sg13g2_decap_8 FILLER_61_417 ();
 sg13g2_decap_4 FILLER_61_424 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_25 ();
 sg13g2_decap_4 FILLER_62_43 ();
 sg13g2_fill_2 FILLER_62_47 ();
 sg13g2_decap_4 FILLER_62_62 ();
 sg13g2_fill_1 FILLER_62_66 ();
 sg13g2_decap_8 FILLER_62_82 ();
 sg13g2_decap_8 FILLER_62_89 ();
 sg13g2_decap_8 FILLER_62_96 ();
 sg13g2_fill_2 FILLER_62_103 ();
 sg13g2_fill_1 FILLER_62_105 ();
 sg13g2_decap_4 FILLER_62_111 ();
 sg13g2_decap_8 FILLER_62_118 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_decap_8 FILLER_62_136 ();
 sg13g2_decap_8 FILLER_62_143 ();
 sg13g2_decap_8 FILLER_62_150 ();
 sg13g2_decap_8 FILLER_62_157 ();
 sg13g2_decap_8 FILLER_62_164 ();
 sg13g2_decap_8 FILLER_62_171 ();
 sg13g2_decap_8 FILLER_62_178 ();
 sg13g2_decap_8 FILLER_62_185 ();
 sg13g2_decap_4 FILLER_62_192 ();
 sg13g2_fill_2 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_fill_1 FILLER_62_209 ();
 sg13g2_decap_8 FILLER_62_216 ();
 sg13g2_fill_1 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_230 ();
 sg13g2_decap_8 FILLER_62_237 ();
 sg13g2_fill_1 FILLER_62_249 ();
 sg13g2_decap_4 FILLER_62_255 ();
 sg13g2_decap_8 FILLER_62_264 ();
 sg13g2_decap_8 FILLER_62_271 ();
 sg13g2_decap_8 FILLER_62_278 ();
 sg13g2_decap_4 FILLER_62_285 ();
 sg13g2_decap_8 FILLER_62_299 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_decap_4 FILLER_62_313 ();
 sg13g2_fill_2 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_fill_2 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_decap_8 FILLER_62_347 ();
 sg13g2_decap_4 FILLER_62_354 ();
 sg13g2_decap_8 FILLER_62_362 ();
 sg13g2_decap_8 FILLER_62_369 ();
 sg13g2_decap_4 FILLER_62_376 ();
 sg13g2_fill_2 FILLER_62_380 ();
 sg13g2_fill_2 FILLER_62_386 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_401 ();
 sg13g2_decap_8 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_62_415 ();
 sg13g2_decap_8 FILLER_62_422 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_37 ();
 sg13g2_decap_8 FILLER_63_44 ();
 sg13g2_decap_8 FILLER_63_51 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_72 ();
 sg13g2_decap_8 FILLER_63_90 ();
 sg13g2_decap_8 FILLER_63_97 ();
 sg13g2_decap_8 FILLER_63_104 ();
 sg13g2_decap_8 FILLER_63_111 ();
 sg13g2_decap_8 FILLER_63_118 ();
 sg13g2_decap_4 FILLER_63_125 ();
 sg13g2_decap_8 FILLER_63_135 ();
 sg13g2_decap_8 FILLER_63_142 ();
 sg13g2_decap_8 FILLER_63_149 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_decap_4 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_165 ();
 sg13g2_fill_2 FILLER_63_182 ();
 sg13g2_fill_1 FILLER_63_184 ();
 sg13g2_decap_8 FILLER_63_190 ();
 sg13g2_decap_8 FILLER_63_197 ();
 sg13g2_decap_8 FILLER_63_204 ();
 sg13g2_decap_8 FILLER_63_211 ();
 sg13g2_decap_4 FILLER_63_218 ();
 sg13g2_decap_4 FILLER_63_226 ();
 sg13g2_fill_1 FILLER_63_230 ();
 sg13g2_decap_4 FILLER_63_237 ();
 sg13g2_decap_4 FILLER_63_256 ();
 sg13g2_decap_8 FILLER_63_264 ();
 sg13g2_decap_4 FILLER_63_271 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_313 ();
 sg13g2_fill_2 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_334 ();
 sg13g2_decap_4 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_345 ();
 sg13g2_decap_8 FILLER_63_351 ();
 sg13g2_fill_2 FILLER_63_358 ();
 sg13g2_decap_4 FILLER_63_377 ();
 sg13g2_fill_2 FILLER_63_385 ();
 sg13g2_fill_1 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_decap_8 FILLER_63_403 ();
 sg13g2_decap_8 FILLER_63_410 ();
 sg13g2_decap_8 FILLER_63_417 ();
 sg13g2_decap_4 FILLER_63_424 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_4 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_39 ();
 sg13g2_decap_8 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_94 ();
 sg13g2_decap_8 FILLER_64_101 ();
 sg13g2_decap_8 FILLER_64_108 ();
 sg13g2_decap_8 FILLER_64_115 ();
 sg13g2_decap_8 FILLER_64_122 ();
 sg13g2_fill_2 FILLER_64_129 ();
 sg13g2_fill_1 FILLER_64_131 ();
 sg13g2_decap_8 FILLER_64_138 ();
 sg13g2_decap_8 FILLER_64_149 ();
 sg13g2_decap_4 FILLER_64_156 ();
 sg13g2_fill_2 FILLER_64_164 ();
 sg13g2_fill_1 FILLER_64_166 ();
 sg13g2_decap_8 FILLER_64_185 ();
 sg13g2_decap_8 FILLER_64_192 ();
 sg13g2_decap_8 FILLER_64_199 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_fill_2 FILLER_64_218 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_decap_4 FILLER_64_263 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_278 ();
 sg13g2_decap_8 FILLER_64_285 ();
 sg13g2_decap_4 FILLER_64_296 ();
 sg13g2_decap_8 FILLER_64_309 ();
 sg13g2_decap_4 FILLER_64_316 ();
 sg13g2_decap_8 FILLER_64_325 ();
 sg13g2_decap_8 FILLER_64_332 ();
 sg13g2_decap_4 FILLER_64_343 ();
 sg13g2_fill_1 FILLER_64_353 ();
 sg13g2_fill_1 FILLER_64_361 ();
 sg13g2_fill_1 FILLER_64_368 ();
 sg13g2_fill_2 FILLER_64_375 ();
 sg13g2_fill_2 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_decap_8 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_64_414 ();
 sg13g2_decap_8 FILLER_64_421 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_81 ();
 sg13g2_decap_8 FILLER_65_88 ();
 sg13g2_decap_8 FILLER_65_95 ();
 sg13g2_decap_8 FILLER_65_102 ();
 sg13g2_decap_8 FILLER_65_109 ();
 sg13g2_decap_8 FILLER_65_116 ();
 sg13g2_fill_2 FILLER_65_123 ();
 sg13g2_decap_4 FILLER_65_133 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_fill_1 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_181 ();
 sg13g2_decap_8 FILLER_65_188 ();
 sg13g2_decap_8 FILLER_65_195 ();
 sg13g2_decap_8 FILLER_65_202 ();
 sg13g2_decap_8 FILLER_65_209 ();
 sg13g2_decap_8 FILLER_65_216 ();
 sg13g2_fill_1 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_decap_4 FILLER_65_237 ();
 sg13g2_fill_2 FILLER_65_241 ();
 sg13g2_decap_8 FILLER_65_248 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_decap_8 FILLER_65_261 ();
 sg13g2_decap_8 FILLER_65_268 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_decap_8 FILLER_65_282 ();
 sg13g2_fill_2 FILLER_65_289 ();
 sg13g2_decap_8 FILLER_65_296 ();
 sg13g2_decap_8 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_326 ();
 sg13g2_decap_4 FILLER_65_335 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_4 FILLER_65_357 ();
 sg13g2_fill_2 FILLER_65_361 ();
 sg13g2_decap_4 FILLER_65_373 ();
 sg13g2_fill_1 FILLER_65_377 ();
 sg13g2_fill_2 FILLER_65_384 ();
 sg13g2_fill_1 FILLER_65_386 ();
 sg13g2_decap_4 FILLER_65_392 ();
 sg13g2_fill_1 FILLER_65_396 ();
 sg13g2_decap_8 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_65_412 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_decap_4 FILLER_65_426 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_4 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_fill_2 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_51 ();
 sg13g2_decap_8 FILLER_66_60 ();
 sg13g2_decap_4 FILLER_66_67 ();
 sg13g2_fill_2 FILLER_66_71 ();
 sg13g2_decap_8 FILLER_66_121 ();
 sg13g2_decap_8 FILLER_66_128 ();
 sg13g2_decap_8 FILLER_66_135 ();
 sg13g2_decap_8 FILLER_66_142 ();
 sg13g2_decap_8 FILLER_66_149 ();
 sg13g2_decap_8 FILLER_66_156 ();
 sg13g2_decap_8 FILLER_66_163 ();
 sg13g2_decap_4 FILLER_66_170 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_decap_8 FILLER_66_180 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_decap_8 FILLER_66_197 ();
 sg13g2_decap_8 FILLER_66_204 ();
 sg13g2_decap_8 FILLER_66_211 ();
 sg13g2_decap_8 FILLER_66_218 ();
 sg13g2_decap_8 FILLER_66_225 ();
 sg13g2_fill_2 FILLER_66_237 ();
 sg13g2_fill_2 FILLER_66_245 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_decap_8 FILLER_66_264 ();
 sg13g2_fill_2 FILLER_66_271 ();
 sg13g2_fill_1 FILLER_66_273 ();
 sg13g2_fill_2 FILLER_66_283 ();
 sg13g2_fill_1 FILLER_66_285 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_fill_1 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_315 ();
 sg13g2_fill_1 FILLER_66_325 ();
 sg13g2_fill_2 FILLER_66_331 ();
 sg13g2_fill_1 FILLER_66_333 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_decap_4 FILLER_66_345 ();
 sg13g2_fill_2 FILLER_66_349 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_decap_4 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_404 ();
 sg13g2_decap_8 FILLER_66_411 ();
 sg13g2_decap_8 FILLER_66_418 ();
 sg13g2_decap_4 FILLER_66_425 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_decap_8 FILLER_67_52 ();
 sg13g2_decap_4 FILLER_67_59 ();
 sg13g2_fill_1 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_69 ();
 sg13g2_decap_8 FILLER_67_76 ();
 sg13g2_decap_8 FILLER_67_83 ();
 sg13g2_decap_8 FILLER_67_90 ();
 sg13g2_decap_4 FILLER_67_97 ();
 sg13g2_fill_1 FILLER_67_101 ();
 sg13g2_decap_8 FILLER_67_106 ();
 sg13g2_decap_8 FILLER_67_113 ();
 sg13g2_fill_2 FILLER_67_120 ();
 sg13g2_fill_1 FILLER_67_122 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_4 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_158 ();
 sg13g2_decap_8 FILLER_67_163 ();
 sg13g2_decap_8 FILLER_67_170 ();
 sg13g2_decap_8 FILLER_67_177 ();
 sg13g2_decap_8 FILLER_67_184 ();
 sg13g2_decap_8 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_198 ();
 sg13g2_decap_4 FILLER_67_205 ();
 sg13g2_fill_1 FILLER_67_209 ();
 sg13g2_decap_8 FILLER_67_214 ();
 sg13g2_fill_2 FILLER_67_221 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_decap_4 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_232 ();
 sg13g2_fill_2 FILLER_67_257 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_265 ();
 sg13g2_fill_2 FILLER_67_271 ();
 sg13g2_fill_1 FILLER_67_284 ();
 sg13g2_decap_8 FILLER_67_290 ();
 sg13g2_fill_1 FILLER_67_297 ();
 sg13g2_decap_4 FILLER_67_313 ();
 sg13g2_fill_2 FILLER_67_317 ();
 sg13g2_decap_4 FILLER_67_324 ();
 sg13g2_fill_1 FILLER_67_338 ();
 sg13g2_decap_8 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_354 ();
 sg13g2_decap_8 FILLER_67_361 ();
 sg13g2_decap_8 FILLER_67_368 ();
 sg13g2_fill_1 FILLER_67_375 ();
 sg13g2_fill_1 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_391 ();
 sg13g2_fill_1 FILLER_67_398 ();
 sg13g2_decap_8 FILLER_67_404 ();
 sg13g2_decap_8 FILLER_67_411 ();
 sg13g2_decap_8 FILLER_67_418 ();
 sg13g2_decap_4 FILLER_67_425 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_decap_8 FILLER_68_44 ();
 sg13g2_decap_4 FILLER_68_51 ();
 sg13g2_decap_8 FILLER_68_83 ();
 sg13g2_decap_8 FILLER_68_90 ();
 sg13g2_decap_8 FILLER_68_97 ();
 sg13g2_decap_8 FILLER_68_104 ();
 sg13g2_decap_8 FILLER_68_111 ();
 sg13g2_decap_8 FILLER_68_118 ();
 sg13g2_decap_8 FILLER_68_125 ();
 sg13g2_fill_1 FILLER_68_132 ();
 sg13g2_decap_8 FILLER_68_136 ();
 sg13g2_decap_8 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_150 ();
 sg13g2_decap_8 FILLER_68_177 ();
 sg13g2_decap_8 FILLER_68_184 ();
 sg13g2_decap_8 FILLER_68_191 ();
 sg13g2_decap_8 FILLER_68_198 ();
 sg13g2_decap_8 FILLER_68_205 ();
 sg13g2_decap_8 FILLER_68_212 ();
 sg13g2_decap_8 FILLER_68_219 ();
 sg13g2_decap_8 FILLER_68_226 ();
 sg13g2_fill_2 FILLER_68_233 ();
 sg13g2_fill_2 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_decap_4 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_264 ();
 sg13g2_fill_2 FILLER_68_269 ();
 sg13g2_decap_8 FILLER_68_276 ();
 sg13g2_decap_4 FILLER_68_283 ();
 sg13g2_fill_2 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_319 ();
 sg13g2_decap_4 FILLER_68_326 ();
 sg13g2_decap_4 FILLER_68_335 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_decap_8 FILLER_68_345 ();
 sg13g2_decap_8 FILLER_68_352 ();
 sg13g2_fill_2 FILLER_68_359 ();
 sg13g2_fill_1 FILLER_68_361 ();
 sg13g2_decap_8 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_386 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_8 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_68_412 ();
 sg13g2_decap_8 FILLER_68_419 ();
 sg13g2_decap_4 FILLER_68_426 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_32 ();
 sg13g2_decap_4 FILLER_69_39 ();
 sg13g2_fill_2 FILLER_69_43 ();
 sg13g2_decap_8 FILLER_69_61 ();
 sg13g2_fill_2 FILLER_69_68 ();
 sg13g2_fill_2 FILLER_69_80 ();
 sg13g2_decap_4 FILLER_69_108 ();
 sg13g2_fill_1 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_fill_2 FILLER_69_168 ();
 sg13g2_fill_1 FILLER_69_178 ();
 sg13g2_decap_8 FILLER_69_187 ();
 sg13g2_decap_8 FILLER_69_194 ();
 sg13g2_decap_8 FILLER_69_201 ();
 sg13g2_decap_8 FILLER_69_208 ();
 sg13g2_decap_4 FILLER_69_215 ();
 sg13g2_decap_4 FILLER_69_224 ();
 sg13g2_fill_2 FILLER_69_228 ();
 sg13g2_decap_4 FILLER_69_239 ();
 sg13g2_fill_1 FILLER_69_243 ();
 sg13g2_decap_8 FILLER_69_248 ();
 sg13g2_decap_8 FILLER_69_255 ();
 sg13g2_decap_8 FILLER_69_262 ();
 sg13g2_decap_8 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_276 ();
 sg13g2_decap_8 FILLER_69_282 ();
 sg13g2_fill_2 FILLER_69_289 ();
 sg13g2_decap_8 FILLER_69_300 ();
 sg13g2_decap_4 FILLER_69_318 ();
 sg13g2_fill_2 FILLER_69_322 ();
 sg13g2_fill_1 FILLER_69_338 ();
 sg13g2_fill_2 FILLER_69_344 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_2 FILLER_69_360 ();
 sg13g2_fill_1 FILLER_69_362 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_fill_2 FILLER_69_388 ();
 sg13g2_fill_2 FILLER_69_400 ();
 sg13g2_decap_8 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_69_414 ();
 sg13g2_decap_8 FILLER_69_421 ();
 sg13g2_fill_2 FILLER_69_428 ();
 sg13g2_decap_8 FILLER_70_26 ();
 sg13g2_decap_4 FILLER_70_45 ();
 sg13g2_fill_1 FILLER_70_49 ();
 sg13g2_fill_2 FILLER_70_70 ();
 sg13g2_fill_1 FILLER_70_72 ();
 sg13g2_fill_1 FILLER_70_77 ();
 sg13g2_decap_4 FILLER_70_86 ();
 sg13g2_decap_8 FILLER_70_94 ();
 sg13g2_decap_8 FILLER_70_101 ();
 sg13g2_decap_8 FILLER_70_108 ();
 sg13g2_fill_2 FILLER_70_115 ();
 sg13g2_fill_1 FILLER_70_117 ();
 sg13g2_fill_2 FILLER_70_129 ();
 sg13g2_fill_2 FILLER_70_141 ();
 sg13g2_fill_2 FILLER_70_177 ();
 sg13g2_decap_8 FILLER_70_192 ();
 sg13g2_decap_8 FILLER_70_199 ();
 sg13g2_decap_8 FILLER_70_206 ();
 sg13g2_decap_8 FILLER_70_213 ();
 sg13g2_decap_8 FILLER_70_220 ();
 sg13g2_decap_8 FILLER_70_227 ();
 sg13g2_fill_2 FILLER_70_234 ();
 sg13g2_fill_1 FILLER_70_236 ();
 sg13g2_decap_4 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_249 ();
 sg13g2_decap_8 FILLER_70_261 ();
 sg13g2_decap_4 FILLER_70_268 ();
 sg13g2_decap_4 FILLER_70_282 ();
 sg13g2_decap_4 FILLER_70_304 ();
 sg13g2_fill_2 FILLER_70_308 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_fill_1 FILLER_70_347 ();
 sg13g2_fill_1 FILLER_70_353 ();
 sg13g2_decap_4 FILLER_70_367 ();
 sg13g2_fill_2 FILLER_70_371 ();
 sg13g2_fill_1 FILLER_70_411 ();
 sg13g2_fill_2 FILLER_70_417 ();
 sg13g2_decap_8 FILLER_70_423 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_13 ();
 sg13g2_decap_8 FILLER_71_20 ();
 sg13g2_decap_8 FILLER_71_27 ();
 sg13g2_decap_4 FILLER_71_60 ();
 sg13g2_fill_2 FILLER_71_64 ();
 sg13g2_decap_8 FILLER_71_92 ();
 sg13g2_decap_8 FILLER_71_99 ();
 sg13g2_decap_8 FILLER_71_106 ();
 sg13g2_fill_2 FILLER_71_113 ();
 sg13g2_decap_4 FILLER_71_123 ();
 sg13g2_fill_1 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_138 ();
 sg13g2_decap_8 FILLER_71_143 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_decap_8 FILLER_71_155 ();
 sg13g2_decap_8 FILLER_71_162 ();
 sg13g2_decap_8 FILLER_71_169 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_188 ();
 sg13g2_decap_8 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_202 ();
 sg13g2_decap_8 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_8 FILLER_71_221 ();
 sg13g2_decap_4 FILLER_71_228 ();
 sg13g2_fill_2 FILLER_71_232 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_267 ();
 sg13g2_fill_2 FILLER_71_280 ();
 sg13g2_fill_2 FILLER_71_293 ();
 sg13g2_decap_8 FILLER_71_303 ();
 sg13g2_decap_8 FILLER_71_310 ();
 sg13g2_decap_4 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_321 ();
 sg13g2_fill_2 FILLER_71_332 ();
 sg13g2_decap_4 FILLER_71_345 ();
 sg13g2_fill_2 FILLER_71_349 ();
 sg13g2_decap_8 FILLER_71_356 ();
 sg13g2_fill_2 FILLER_71_363 ();
 sg13g2_fill_1 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_398 ();
 sg13g2_decap_8 FILLER_71_405 ();
 sg13g2_decap_8 FILLER_71_412 ();
 sg13g2_decap_8 FILLER_71_419 ();
 sg13g2_decap_4 FILLER_71_426 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_4 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_45 ();
 sg13g2_decap_8 FILLER_72_60 ();
 sg13g2_decap_8 FILLER_72_67 ();
 sg13g2_decap_8 FILLER_72_74 ();
 sg13g2_decap_4 FILLER_72_81 ();
 sg13g2_fill_1 FILLER_72_85 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_4 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_222 ();
 sg13g2_decap_8 FILLER_72_229 ();
 sg13g2_decap_8 FILLER_72_236 ();
 sg13g2_fill_2 FILLER_72_251 ();
 sg13g2_fill_1 FILLER_72_253 ();
 sg13g2_decap_4 FILLER_72_271 ();
 sg13g2_fill_2 FILLER_72_275 ();
 sg13g2_decap_8 FILLER_72_285 ();
 sg13g2_decap_4 FILLER_72_292 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_4 FILLER_72_315 ();
 sg13g2_fill_2 FILLER_72_319 ();
 sg13g2_decap_8 FILLER_72_334 ();
 sg13g2_decap_8 FILLER_72_341 ();
 sg13g2_fill_1 FILLER_72_348 ();
 sg13g2_decap_8 FILLER_72_355 ();
 sg13g2_fill_2 FILLER_72_362 ();
 sg13g2_fill_1 FILLER_72_364 ();
 sg13g2_fill_2 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_72_388 ();
 sg13g2_decap_8 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_72_409 ();
 sg13g2_decap_8 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_21 ();
 sg13g2_decap_4 FILLER_73_30 ();
 sg13g2_decap_8 FILLER_73_44 ();
 sg13g2_decap_8 FILLER_73_51 ();
 sg13g2_decap_8 FILLER_73_58 ();
 sg13g2_decap_8 FILLER_73_65 ();
 sg13g2_decap_8 FILLER_73_72 ();
 sg13g2_decap_8 FILLER_73_79 ();
 sg13g2_decap_8 FILLER_73_86 ();
 sg13g2_fill_2 FILLER_73_93 ();
 sg13g2_fill_1 FILLER_73_95 ();
 sg13g2_decap_8 FILLER_73_104 ();
 sg13g2_decap_8 FILLER_73_111 ();
 sg13g2_fill_2 FILLER_73_123 ();
 sg13g2_decap_4 FILLER_73_133 ();
 sg13g2_fill_2 FILLER_73_137 ();
 sg13g2_fill_2 FILLER_73_165 ();
 sg13g2_fill_1 FILLER_73_167 ();
 sg13g2_fill_1 FILLER_73_181 ();
 sg13g2_decap_8 FILLER_73_191 ();
 sg13g2_decap_8 FILLER_73_198 ();
 sg13g2_decap_8 FILLER_73_205 ();
 sg13g2_decap_8 FILLER_73_212 ();
 sg13g2_fill_2 FILLER_73_219 ();
 sg13g2_decap_8 FILLER_73_225 ();
 sg13g2_decap_8 FILLER_73_232 ();
 sg13g2_decap_4 FILLER_73_239 ();
 sg13g2_fill_1 FILLER_73_243 ();
 sg13g2_decap_8 FILLER_73_256 ();
 sg13g2_decap_8 FILLER_73_263 ();
 sg13g2_decap_8 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_fill_2 FILLER_73_283 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_decap_8 FILLER_73_293 ();
 sg13g2_decap_8 FILLER_73_300 ();
 sg13g2_decap_8 FILLER_73_307 ();
 sg13g2_decap_8 FILLER_73_314 ();
 sg13g2_decap_8 FILLER_73_321 ();
 sg13g2_decap_8 FILLER_73_328 ();
 sg13g2_decap_8 FILLER_73_335 ();
 sg13g2_fill_2 FILLER_73_342 ();
 sg13g2_decap_8 FILLER_73_354 ();
 sg13g2_decap_8 FILLER_73_361 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_fill_2 FILLER_73_375 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_decap_8 FILLER_73_384 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_8 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_73_412 ();
 sg13g2_decap_8 FILLER_73_419 ();
 sg13g2_decap_4 FILLER_73_426 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_26 ();
 sg13g2_fill_2 FILLER_74_33 ();
 sg13g2_fill_1 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_62 ();
 sg13g2_decap_8 FILLER_74_69 ();
 sg13g2_decap_8 FILLER_74_76 ();
 sg13g2_decap_8 FILLER_74_83 ();
 sg13g2_decap_8 FILLER_74_90 ();
 sg13g2_fill_2 FILLER_74_112 ();
 sg13g2_decap_4 FILLER_74_122 ();
 sg13g2_decap_8 FILLER_74_131 ();
 sg13g2_decap_8 FILLER_74_138 ();
 sg13g2_fill_1 FILLER_74_145 ();
 sg13g2_decap_8 FILLER_74_150 ();
 sg13g2_decap_8 FILLER_74_157 ();
 sg13g2_decap_8 FILLER_74_164 ();
 sg13g2_fill_2 FILLER_74_171 ();
 sg13g2_decap_8 FILLER_74_183 ();
 sg13g2_decap_4 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_199 ();
 sg13g2_decap_8 FILLER_74_205 ();
 sg13g2_decap_8 FILLER_74_212 ();
 sg13g2_decap_8 FILLER_74_219 ();
 sg13g2_decap_8 FILLER_74_226 ();
 sg13g2_decap_8 FILLER_74_233 ();
 sg13g2_decap_8 FILLER_74_240 ();
 sg13g2_decap_8 FILLER_74_247 ();
 sg13g2_decap_4 FILLER_74_270 ();
 sg13g2_decap_4 FILLER_74_282 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_2 FILLER_74_297 ();
 sg13g2_decap_8 FILLER_74_304 ();
 sg13g2_decap_4 FILLER_74_311 ();
 sg13g2_fill_2 FILLER_74_315 ();
 sg13g2_decap_4 FILLER_74_320 ();
 sg13g2_decap_8 FILLER_74_330 ();
 sg13g2_decap_8 FILLER_74_337 ();
 sg13g2_decap_8 FILLER_74_344 ();
 sg13g2_decap_8 FILLER_74_351 ();
 sg13g2_fill_1 FILLER_74_362 ();
 sg13g2_decap_4 FILLER_74_367 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_decap_8 FILLER_74_404 ();
 sg13g2_decap_8 FILLER_74_411 ();
 sg13g2_decap_8 FILLER_74_418 ();
 sg13g2_decap_4 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_30 ();
 sg13g2_decap_4 FILLER_75_37 ();
 sg13g2_fill_1 FILLER_75_41 ();
 sg13g2_fill_1 FILLER_75_54 ();
 sg13g2_fill_2 FILLER_75_108 ();
 sg13g2_decap_8 FILLER_75_118 ();
 sg13g2_decap_8 FILLER_75_125 ();
 sg13g2_fill_1 FILLER_75_132 ();
 sg13g2_decap_8 FILLER_75_159 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_185 ();
 sg13g2_fill_2 FILLER_75_192 ();
 sg13g2_fill_1 FILLER_75_194 ();
 sg13g2_decap_8 FILLER_75_221 ();
 sg13g2_decap_8 FILLER_75_228 ();
 sg13g2_decap_8 FILLER_75_235 ();
 sg13g2_decap_8 FILLER_75_242 ();
 sg13g2_fill_2 FILLER_75_249 ();
 sg13g2_fill_1 FILLER_75_251 ();
 sg13g2_fill_2 FILLER_75_257 ();
 sg13g2_fill_1 FILLER_75_259 ();
 sg13g2_fill_2 FILLER_75_265 ();
 sg13g2_fill_2 FILLER_75_278 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_fill_2 FILLER_75_294 ();
 sg13g2_fill_2 FILLER_75_312 ();
 sg13g2_decap_8 FILLER_75_330 ();
 sg13g2_fill_2 FILLER_75_337 ();
 sg13g2_fill_2 FILLER_75_356 ();
 sg13g2_fill_2 FILLER_75_363 ();
 sg13g2_fill_2 FILLER_75_370 ();
 sg13g2_fill_2 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_384 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_8 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_75_412 ();
 sg13g2_decap_8 FILLER_75_419 ();
 sg13g2_decap_4 FILLER_75_426 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_15 ();
 sg13g2_decap_8 FILLER_76_22 ();
 sg13g2_decap_4 FILLER_76_29 ();
 sg13g2_fill_2 FILLER_76_33 ();
 sg13g2_decap_8 FILLER_76_53 ();
 sg13g2_decap_8 FILLER_76_60 ();
 sg13g2_decap_4 FILLER_76_67 ();
 sg13g2_decap_8 FILLER_76_75 ();
 sg13g2_decap_8 FILLER_76_82 ();
 sg13g2_fill_2 FILLER_76_89 ();
 sg13g2_decap_4 FILLER_76_95 ();
 sg13g2_fill_1 FILLER_76_106 ();
 sg13g2_fill_2 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_118 ();
 sg13g2_decap_8 FILLER_76_125 ();
 sg13g2_decap_4 FILLER_76_132 ();
 sg13g2_fill_1 FILLER_76_136 ();
 sg13g2_decap_8 FILLER_76_141 ();
 sg13g2_decap_8 FILLER_76_148 ();
 sg13g2_decap_8 FILLER_76_155 ();
 sg13g2_decap_8 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_169 ();
 sg13g2_decap_8 FILLER_76_176 ();
 sg13g2_decap_4 FILLER_76_183 ();
 sg13g2_fill_1 FILLER_76_187 ();
 sg13g2_decap_4 FILLER_76_193 ();
 sg13g2_fill_1 FILLER_76_197 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_fill_2 FILLER_76_210 ();
 sg13g2_fill_1 FILLER_76_212 ();
 sg13g2_decap_4 FILLER_76_218 ();
 sg13g2_fill_1 FILLER_76_222 ();
 sg13g2_decap_8 FILLER_76_228 ();
 sg13g2_decap_8 FILLER_76_235 ();
 sg13g2_decap_8 FILLER_76_242 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_76_256 ();
 sg13g2_decap_4 FILLER_76_263 ();
 sg13g2_fill_1 FILLER_76_267 ();
 sg13g2_decap_4 FILLER_76_273 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_fill_1 FILLER_76_302 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_fill_1 FILLER_76_347 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_fill_2 FILLER_76_362 ();
 sg13g2_decap_4 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_decap_8 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_44 ();
 sg13g2_decap_8 FILLER_77_51 ();
 sg13g2_decap_8 FILLER_77_58 ();
 sg13g2_decap_8 FILLER_77_65 ();
 sg13g2_decap_8 FILLER_77_72 ();
 sg13g2_fill_1 FILLER_77_79 ();
 sg13g2_fill_2 FILLER_77_85 ();
 sg13g2_fill_1 FILLER_77_87 ();
 sg13g2_decap_4 FILLER_77_96 ();
 sg13g2_fill_2 FILLER_77_100 ();
 sg13g2_decap_8 FILLER_77_132 ();
 sg13g2_decap_8 FILLER_77_139 ();
 sg13g2_decap_8 FILLER_77_146 ();
 sg13g2_decap_4 FILLER_77_153 ();
 sg13g2_decap_8 FILLER_77_172 ();
 sg13g2_decap_8 FILLER_77_179 ();
 sg13g2_decap_8 FILLER_77_186 ();
 sg13g2_decap_8 FILLER_77_193 ();
 sg13g2_decap_8 FILLER_77_200 ();
 sg13g2_decap_8 FILLER_77_207 ();
 sg13g2_decap_8 FILLER_77_214 ();
 sg13g2_decap_8 FILLER_77_221 ();
 sg13g2_decap_8 FILLER_77_228 ();
 sg13g2_decap_8 FILLER_77_235 ();
 sg13g2_decap_8 FILLER_77_242 ();
 sg13g2_decap_8 FILLER_77_249 ();
 sg13g2_decap_8 FILLER_77_256 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_decap_8 FILLER_77_270 ();
 sg13g2_decap_8 FILLER_77_277 ();
 sg13g2_decap_8 FILLER_77_284 ();
 sg13g2_decap_4 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_295 ();
 sg13g2_fill_2 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_318 ();
 sg13g2_decap_4 FILLER_77_324 ();
 sg13g2_fill_1 FILLER_77_328 ();
 sg13g2_fill_2 FILLER_77_351 ();
 sg13g2_fill_2 FILLER_77_367 ();
 sg13g2_decap_8 FILLER_77_373 ();
 sg13g2_decap_8 FILLER_77_380 ();
 sg13g2_decap_8 FILLER_77_387 ();
 sg13g2_decap_8 FILLER_77_394 ();
 sg13g2_decap_8 FILLER_77_401 ();
 sg13g2_decap_8 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_77_415 ();
 sg13g2_decap_8 FILLER_77_422 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_25 ();
 sg13g2_decap_8 FILLER_78_32 ();
 sg13g2_decap_8 FILLER_78_39 ();
 sg13g2_decap_8 FILLER_78_46 ();
 sg13g2_decap_8 FILLER_78_53 ();
 sg13g2_decap_8 FILLER_78_60 ();
 sg13g2_decap_4 FILLER_78_67 ();
 sg13g2_fill_1 FILLER_78_71 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_fill_2 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_118 ();
 sg13g2_decap_8 FILLER_78_125 ();
 sg13g2_fill_2 FILLER_78_132 ();
 sg13g2_fill_2 FILLER_78_216 ();
 sg13g2_decap_4 FILLER_78_222 ();
 sg13g2_fill_1 FILLER_78_226 ();
 sg13g2_decap_8 FILLER_78_253 ();
 sg13g2_decap_8 FILLER_78_260 ();
 sg13g2_decap_8 FILLER_78_267 ();
 sg13g2_decap_8 FILLER_78_274 ();
 sg13g2_decap_8 FILLER_78_281 ();
 sg13g2_decap_8 FILLER_78_288 ();
 sg13g2_decap_8 FILLER_78_295 ();
 sg13g2_decap_4 FILLER_78_302 ();
 sg13g2_decap_8 FILLER_78_310 ();
 sg13g2_decap_8 FILLER_78_317 ();
 sg13g2_fill_2 FILLER_78_324 ();
 sg13g2_decap_8 FILLER_78_330 ();
 sg13g2_decap_8 FILLER_78_337 ();
 sg13g2_decap_8 FILLER_78_344 ();
 sg13g2_decap_8 FILLER_78_351 ();
 sg13g2_decap_8 FILLER_78_358 ();
 sg13g2_decap_8 FILLER_78_365 ();
 sg13g2_decap_8 FILLER_78_372 ();
 sg13g2_decap_8 FILLER_78_379 ();
 sg13g2_decap_8 FILLER_78_386 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_decap_8 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_78_414 ();
 sg13g2_decap_8 FILLER_78_421 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_fill_2 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_83 ();
 sg13g2_fill_1 FILLER_79_87 ();
 sg13g2_decap_8 FILLER_79_92 ();
 sg13g2_decap_8 FILLER_79_99 ();
 sg13g2_decap_8 FILLER_79_106 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_fill_1 FILLER_79_120 ();
 sg13g2_decap_8 FILLER_79_125 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_4 FILLER_79_139 ();
 sg13g2_fill_2 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_184 ();
 sg13g2_decap_8 FILLER_79_195 ();
 sg13g2_decap_4 FILLER_79_202 ();
 sg13g2_fill_1 FILLER_79_206 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_fill_2 FILLER_79_427 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_74 ();
 sg13g2_fill_2 FILLER_80_80 ();
 sg13g2_fill_1 FILLER_80_90 ();
 sg13g2_fill_2 FILLER_80_119 ();
 sg13g2_fill_2 FILLER_80_125 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_fill_2 FILLER_80_144 ();
 sg13g2_fill_2 FILLER_80_170 ();
 sg13g2_fill_1 FILLER_80_172 ();
 sg13g2_fill_1 FILLER_80_177 ();
 sg13g2_decap_4 FILLER_80_182 ();
 sg13g2_fill_2 FILLER_80_198 ();
 sg13g2_fill_1 FILLER_80_200 ();
 sg13g2_fill_2 FILLER_80_209 ();
 sg13g2_fill_1 FILLER_80_211 ();
 sg13g2_fill_1 FILLER_80_220 ();
 sg13g2_fill_2 FILLER_80_225 ();
 sg13g2_fill_1 FILLER_80_227 ();
 sg13g2_fill_2 FILLER_80_240 ();
 sg13g2_decap_4 FILLER_80_246 ();
 sg13g2_decap_4 FILLER_80_254 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_355 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_decap_4 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_decap_8 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_8 FILLER_80_404 ();
 sg13g2_decap_8 FILLER_80_411 ();
 sg13g2_decap_8 FILLER_80_418 ();
 sg13g2_decap_4 FILLER_80_425 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
