module tt_um_stochastic_addmultiply_CL123abc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire SN_Bit_1;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire clknet_leaf_0_clk;
 wire net95;
 wire \add_avg[0] ;
 wire \add_avg[1] ;
 wire \add_avg[2] ;
 wire \add_avg[3] ;
 wire \add_avg[4] ;
 wire \add_avg[5] ;
 wire \add_avg[6] ;
 wire \add_avg[7] ;
 wire \add_avg[8] ;
 wire add_bit_out;
 wire \add_output.bitseq[0] ;
 wire \add_output.bitseq[1] ;
 wire \add_output.bitseq[2] ;
 wire \add_output.bitseq[3] ;
 wire \add_output.bitseq[4] ;
 wire \add_output.bitseq[5] ;
 wire \add_output.bitseq[6] ;
 wire \add_output.bitseq[7] ;
 wire \add_output.bitseq[8] ;
 wire \add_output.counter[0] ;
 wire \add_output.counter[1] ;
 wire \add_output.counter[2] ;
 wire \add_output.counter[3] ;
 wire \add_up_counter.clk_counter[0] ;
 wire \add_up_counter.clk_counter[10] ;
 wire \add_up_counter.clk_counter[11] ;
 wire \add_up_counter.clk_counter[12] ;
 wire \add_up_counter.clk_counter[13] ;
 wire \add_up_counter.clk_counter[14] ;
 wire \add_up_counter.clk_counter[15] ;
 wire \add_up_counter.clk_counter[16] ;
 wire \add_up_counter.clk_counter[17] ;
 wire \add_up_counter.clk_counter[1] ;
 wire \add_up_counter.clk_counter[2] ;
 wire \add_up_counter.clk_counter[3] ;
 wire \add_up_counter.clk_counter[4] ;
 wire \add_up_counter.clk_counter[5] ;
 wire \add_up_counter.clk_counter[6] ;
 wire \add_up_counter.clk_counter[7] ;
 wire \add_up_counter.clk_counter[8] ;
 wire \add_up_counter.clk_counter[9] ;
 wire \add_up_counter.prob_counter[0] ;
 wire \add_up_counter.prob_counter[10] ;
 wire \add_up_counter.prob_counter[11] ;
 wire \add_up_counter.prob_counter[12] ;
 wire \add_up_counter.prob_counter[13] ;
 wire \add_up_counter.prob_counter[14] ;
 wire \add_up_counter.prob_counter[15] ;
 wire \add_up_counter.prob_counter[16] ;
 wire \add_up_counter.prob_counter[1] ;
 wire \add_up_counter.prob_counter[2] ;
 wire \add_up_counter.prob_counter[3] ;
 wire \add_up_counter.prob_counter[4] ;
 wire \add_up_counter.prob_counter[5] ;
 wire \add_up_counter.prob_counter[6] ;
 wire \add_up_counter.prob_counter[7] ;
 wire \add_up_counter.prob_counter[8] ;
 wire \add_up_counter.prob_counter[9] ;
 wire \global_SN_gen.Input_1[0] ;
 wire \global_SN_gen.Input_1[1] ;
 wire \global_SN_gen.Input_1[2] ;
 wire \global_SN_gen.Input_1[3] ;
 wire \global_SN_gen.Input_1[4] ;
 wire \global_SN_gen.Input_1[5] ;
 wire \global_SN_gen.Input_1[6] ;
 wire \global_SN_gen.Input_1[7] ;
 wire \global_SN_gen.Input_1[8] ;
 wire \global_SN_gen.Input_2[0] ;
 wire \global_SN_gen.Input_2[1] ;
 wire \global_SN_gen.Input_2[2] ;
 wire \global_SN_gen.Input_2[3] ;
 wire \global_SN_gen.Input_2[4] ;
 wire \global_SN_gen.Input_2[5] ;
 wire \global_SN_gen.Input_2[6] ;
 wire \global_SN_gen.Input_2[7] ;
 wire \global_SN_gen.Input_2[8] ;
 wire \global_SN_gen.lfsr[0] ;
 wire \global_SN_gen.lfsr[10] ;
 wire \global_SN_gen.lfsr[11] ;
 wire \global_SN_gen.lfsr[12] ;
 wire \global_SN_gen.lfsr[13] ;
 wire \global_SN_gen.lfsr[14] ;
 wire \global_SN_gen.lfsr[15] ;
 wire \global_SN_gen.lfsr[16] ;
 wire \global_SN_gen.lfsr[17] ;
 wire \global_SN_gen.lfsr[18] ;
 wire \global_SN_gen.lfsr[19] ;
 wire \global_SN_gen.lfsr[1] ;
 wire \global_SN_gen.lfsr[20] ;
 wire \global_SN_gen.lfsr[21] ;
 wire \global_SN_gen.lfsr[22] ;
 wire \global_SN_gen.lfsr[23] ;
 wire \global_SN_gen.lfsr[24] ;
 wire \global_SN_gen.lfsr[25] ;
 wire \global_SN_gen.lfsr[26] ;
 wire \global_SN_gen.lfsr[27] ;
 wire \global_SN_gen.lfsr[28] ;
 wire \global_SN_gen.lfsr[29] ;
 wire \global_SN_gen.lfsr[2] ;
 wire \global_SN_gen.lfsr[30] ;
 wire \global_SN_gen.lfsr[3] ;
 wire \global_SN_gen.lfsr[4] ;
 wire \global_SN_gen.lfsr[5] ;
 wire \global_SN_gen.lfsr[6] ;
 wire \global_SN_gen.lfsr[7] ;
 wire \global_SN_gen.lfsr[8] ;
 wire \global_SN_gen.lfsr[9] ;
 wire \global_input.adjustment[0] ;
 wire \global_input.adjustment[1] ;
 wire \global_input.adjustment[2] ;
 wire \global_input.adjustment[3] ;
 wire \global_input.adjustment[4] ;
 wire \global_input.loop ;
 wire \global_input.output_bitcounter_1[0] ;
 wire \global_input.output_bitcounter_1[1] ;
 wire \global_input.output_bitcounter_1[2] ;
 wire \global_input.output_bitcounter_1[3] ;
 wire \global_input.output_bitcounter_1[4] ;
 wire \global_input.output_bitcounter_1[5] ;
 wire \global_input.output_bitcounter_1[6] ;
 wire \global_input.output_bitcounter_1[7] ;
 wire \global_input.output_bitcounter_1[8] ;
 wire \global_input.output_bitcounter_2[0] ;
 wire \global_input.output_bitcounter_2[1] ;
 wire \global_input.output_bitcounter_2[2] ;
 wire \global_input.output_bitcounter_2[3] ;
 wire \global_input.output_bitcounter_2[4] ;
 wire \global_input.output_bitcounter_2[5] ;
 wire \global_input.output_bitcounter_2[6] ;
 wire \global_input.output_bitcounter_2[7] ;
 wire \global_input.output_bitcounter_2[8] ;
 wire \global_input.output_case[0] ;
 wire \global_input.output_case[1] ;
 wire \global_input.output_case[2] ;
 wire \global_input.output_case[3] ;
 wire \mul_avg[0] ;
 wire \mul_avg[1] ;
 wire \mul_avg[2] ;
 wire \mul_avg[3] ;
 wire \mul_avg[4] ;
 wire \mul_avg[5] ;
 wire \mul_avg[6] ;
 wire \mul_avg[7] ;
 wire \mul_avg[8] ;
 wire mul_bit_out;
 wire \mul_output.bitseq[0] ;
 wire \mul_output.bitseq[1] ;
 wire \mul_output.bitseq[2] ;
 wire \mul_output.bitseq[3] ;
 wire \mul_output.bitseq[4] ;
 wire \mul_output.bitseq[5] ;
 wire \mul_output.bitseq[6] ;
 wire \mul_output.bitseq[7] ;
 wire \mul_output.bitseq[8] ;
 wire \mul_output.counter[0] ;
 wire \mul_output.counter[1] ;
 wire \mul_output.counter[2] ;
 wire \mul_output.counter[3] ;
 wire \mul_up_counter.prob_counter[0] ;
 wire \mul_up_counter.prob_counter[10] ;
 wire \mul_up_counter.prob_counter[11] ;
 wire \mul_up_counter.prob_counter[12] ;
 wire \mul_up_counter.prob_counter[13] ;
 wire \mul_up_counter.prob_counter[14] ;
 wire \mul_up_counter.prob_counter[15] ;
 wire \mul_up_counter.prob_counter[16] ;
 wire \mul_up_counter.prob_counter[1] ;
 wire \mul_up_counter.prob_counter[2] ;
 wire \mul_up_counter.prob_counter[3] ;
 wire \mul_up_counter.prob_counter[4] ;
 wire \mul_up_counter.prob_counter[5] ;
 wire \mul_up_counter.prob_counter[6] ;
 wire \mul_up_counter.prob_counter[7] ;
 wire \mul_up_counter.prob_counter[8] ;
 wire \mul_up_counter.prob_counter[9] ;
 wire \smul.SN_Bit_Q ;
 wire \smul_avg[0] ;
 wire \smul_avg[1] ;
 wire \smul_avg[2] ;
 wire \smul_avg[3] ;
 wire \smul_avg[4] ;
 wire \smul_avg[5] ;
 wire \smul_avg[6] ;
 wire \smul_avg[7] ;
 wire \smul_avg[8] ;
 wire smul_bit_out;
 wire \smul_output.bitseq[0] ;
 wire \smul_output.bitseq[1] ;
 wire \smul_output.bitseq[2] ;
 wire \smul_output.bitseq[3] ;
 wire \smul_output.bitseq[4] ;
 wire \smul_output.bitseq[5] ;
 wire \smul_output.bitseq[6] ;
 wire \smul_output.bitseq[7] ;
 wire \smul_output.bitseq[8] ;
 wire \smul_output.counter[0] ;
 wire \smul_output.counter[1] ;
 wire \smul_output.counter[2] ;
 wire \smul_output.counter[3] ;
 wire \smul_up_counter.prob_counter[0] ;
 wire \smul_up_counter.prob_counter[10] ;
 wire \smul_up_counter.prob_counter[11] ;
 wire \smul_up_counter.prob_counter[12] ;
 wire \smul_up_counter.prob_counter[13] ;
 wire \smul_up_counter.prob_counter[14] ;
 wire \smul_up_counter.prob_counter[15] ;
 wire \smul_up_counter.prob_counter[16] ;
 wire \smul_up_counter.prob_counter[1] ;
 wire \smul_up_counter.prob_counter[2] ;
 wire \smul_up_counter.prob_counter[3] ;
 wire \smul_up_counter.prob_counter[4] ;
 wire \smul_up_counter.prob_counter[5] ;
 wire \smul_up_counter.prob_counter[6] ;
 wire \smul_up_counter.prob_counter[7] ;
 wire \smul_up_counter.prob_counter[8] ;
 wire \smul_up_counter.prob_counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _0910_ (.Y(_0232_),
    .A(\global_SN_gen.Input_1[8] ));
 sg13g2_inv_1 _0911_ (.Y(_0233_),
    .A(\global_SN_gen.Input_1[1] ));
 sg13g2_nand2b_1 _0912_ (.Y(_0234_),
    .B(\global_SN_gen.Input_1[0] ),
    .A_N(\global_SN_gen.lfsr[0] ));
 sg13g2_a21oi_1 _0913_ (.A1(_0233_),
    .A2(\global_SN_gen.lfsr[1] ),
    .Y(_0235_),
    .B1(_0234_));
 sg13g2_nand2b_1 _0914_ (.Y(_0236_),
    .B(\global_SN_gen.Input_1[2] ),
    .A_N(\global_SN_gen.lfsr[2] ));
 sg13g2_o21ai_1 _0915_ (.B1(_0236_),
    .Y(_0237_),
    .A1(_0233_),
    .A2(\global_SN_gen.lfsr[1] ));
 sg13g2_buf_2 _0916_ (.A(\global_SN_gen.Input_1[3] ),
    .X(_0238_));
 sg13g2_xor2_1 _0917_ (.B(\global_SN_gen.lfsr[3] ),
    .A(_0238_),
    .X(_0239_));
 sg13g2_nor2b_1 _0918_ (.A(\global_SN_gen.Input_1[2] ),
    .B_N(\global_SN_gen.lfsr[2] ),
    .Y(_0240_));
 sg13g2_xor2_1 _0919_ (.B(\global_SN_gen.lfsr[4] ),
    .A(\global_SN_gen.Input_1[4] ),
    .X(_0241_));
 sg13g2_nor3_1 _0920_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_o21ai_1 _0921_ (.B1(_0242_),
    .Y(_0243_),
    .A1(_0235_),
    .A2(_0237_));
 sg13g2_nand2b_1 _0922_ (.Y(_0244_),
    .B(_0238_),
    .A_N(\global_SN_gen.lfsr[3] ));
 sg13g2_inv_1 _0923_ (.Y(_0245_),
    .A(\global_SN_gen.Input_1[4] ));
 sg13g2_a21oi_1 _0924_ (.A1(\global_SN_gen.lfsr[4] ),
    .A2(_0244_),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_nand2b_1 _0925_ (.Y(_0247_),
    .B(\global_SN_gen.Input_1[6] ),
    .A_N(\global_SN_gen.lfsr[6] ));
 sg13g2_nand2b_1 _0926_ (.Y(_0248_),
    .B(\global_SN_gen.Input_1[7] ),
    .A_N(\global_SN_gen.lfsr[7] ));
 sg13g2_nand2b_1 _0927_ (.Y(_0249_),
    .B(\global_SN_gen.Input_1[5] ),
    .A_N(\global_SN_gen.lfsr[5] ));
 sg13g2_nand3_1 _0928_ (.B(_0248_),
    .C(_0249_),
    .A(_0247_),
    .Y(_0250_));
 sg13g2_nor2_1 _0929_ (.A(\global_SN_gen.lfsr[4] ),
    .B(_0244_),
    .Y(_0251_));
 sg13g2_nor3_1 _0930_ (.A(_0246_),
    .B(_0250_),
    .C(_0251_),
    .Y(_0252_));
 sg13g2_nor2b_1 _0931_ (.A(\global_SN_gen.Input_1[7] ),
    .B_N(\global_SN_gen.lfsr[7] ),
    .Y(_0253_));
 sg13g2_nor2b_1 _0932_ (.A(\global_SN_gen.Input_1[6] ),
    .B_N(\global_SN_gen.lfsr[6] ),
    .Y(_0254_));
 sg13g2_o21ai_1 _0933_ (.B1(_0248_),
    .Y(_0255_),
    .A1(_0253_),
    .A2(_0254_));
 sg13g2_inv_1 _0934_ (.Y(_0256_),
    .A(\global_SN_gen.Input_1[5] ));
 sg13g2_nand4_1 _0935_ (.B(\global_SN_gen.lfsr[5] ),
    .C(_0247_),
    .A(_0256_),
    .Y(_0257_),
    .D(_0248_));
 sg13g2_nand2_1 _0936_ (.Y(_0258_),
    .A(_0255_),
    .B(_0257_));
 sg13g2_a221oi_1 _0937_ (.B2(_0252_),
    .C1(_0258_),
    .B1(_0243_),
    .A1(_0232_),
    .Y(_0259_),
    .A2(\global_SN_gen.lfsr[8] ));
 sg13g2_nor2_1 _0938_ (.A(_0232_),
    .B(\global_SN_gen.lfsr[8] ),
    .Y(_0260_));
 sg13g2_nor2_1 _0939_ (.A(_0259_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_inv_1 _0940_ (.Y(SN_Bit_1),
    .A(_0261_));
 sg13g2_buf_2 _0941_ (.A(\mul_output.counter[1] ),
    .X(_0262_));
 sg13g2_buf_1 _0942_ (.A(\mul_output.counter[0] ),
    .X(_0263_));
 sg13g2_nor4_2 _0943_ (.A(_0262_),
    .B(_0263_),
    .C(\mul_output.counter[2] ),
    .Y(_0264_),
    .D(\mul_output.counter[3] ));
 sg13g2_buf_1 _0944_ (.A(_0264_),
    .X(_0265_));
 sg13g2_inv_1 _0945_ (.Y(_0131_),
    .A(_0263_));
 sg13g2_inv_1 _0946_ (.Y(_0266_),
    .A(\mul_output.counter[2] ));
 sg13g2_nand2_1 _0947_ (.Y(_0267_),
    .A(_0266_),
    .B(\mul_output.counter[3] ));
 sg13g2_nor3_2 _0948_ (.A(_0262_),
    .B(_0131_),
    .C(_0267_),
    .Y(_0268_));
 sg13g2_buf_1 _0949_ (.A(_0268_),
    .X(_0269_));
 sg13g2_a22oi_1 _0950_ (.Y(_0270_),
    .B1(net30),
    .B2(\mul_output.bitseq[0] ),
    .A2(net33),
    .A1(\mul_avg[1] ));
 sg13g2_nor2_2 _0951_ (.A(_0264_),
    .B(_0268_),
    .Y(_0271_));
 sg13g2_nand2_1 _0952_ (.Y(_0272_),
    .A(\mul_output.bitseq[1] ),
    .B(_0271_));
 sg13g2_nand2_1 _0953_ (.Y(_0028_),
    .A(_0270_),
    .B(_0272_));
 sg13g2_a22oi_1 _0954_ (.Y(_0273_),
    .B1(net30),
    .B2(\mul_output.bitseq[1] ),
    .A2(net33),
    .A1(\mul_avg[2] ));
 sg13g2_nand2_1 _0955_ (.Y(_0274_),
    .A(\mul_output.bitseq[2] ),
    .B(_0271_));
 sg13g2_nand2_1 _0956_ (.Y(_0029_),
    .A(_0273_),
    .B(_0274_));
 sg13g2_a22oi_1 _0957_ (.Y(_0275_),
    .B1(_0269_),
    .B2(\mul_output.bitseq[2] ),
    .A2(net33),
    .A1(\mul_avg[3] ));
 sg13g2_nand2_1 _0958_ (.Y(_0276_),
    .A(\mul_output.bitseq[3] ),
    .B(_0271_));
 sg13g2_nand2_1 _0959_ (.Y(_0030_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_nor2b_1 _0960_ (.A(_0268_),
    .B_N(\mul_output.bitseq[4] ),
    .Y(_0277_));
 sg13g2_a21oi_1 _0961_ (.A1(\mul_output.bitseq[3] ),
    .A2(net30),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_nand2_1 _0962_ (.Y(_0279_),
    .A(\mul_avg[4] ),
    .B(_0265_));
 sg13g2_o21ai_1 _0963_ (.B1(_0279_),
    .Y(_0031_),
    .A1(_0265_),
    .A2(_0278_));
 sg13g2_nor2b_1 _0964_ (.A(_0268_),
    .B_N(\mul_output.bitseq[5] ),
    .Y(_0280_));
 sg13g2_a21oi_1 _0965_ (.A1(\mul_output.bitseq[4] ),
    .A2(_0269_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nand2_1 _0966_ (.Y(_0282_),
    .A(\mul_avg[5] ),
    .B(net33));
 sg13g2_o21ai_1 _0967_ (.B1(_0282_),
    .Y(_0032_),
    .A1(net33),
    .A2(_0281_));
 sg13g2_a22oi_1 _0968_ (.Y(_0283_),
    .B1(net30),
    .B2(\mul_output.bitseq[5] ),
    .A2(_0264_),
    .A1(\mul_avg[6] ));
 sg13g2_nand2_1 _0969_ (.Y(_0284_),
    .A(\mul_output.bitseq[6] ),
    .B(_0271_));
 sg13g2_nand2_1 _0970_ (.Y(_0033_),
    .A(_0283_),
    .B(_0284_));
 sg13g2_a22oi_1 _0971_ (.Y(_0285_),
    .B1(net30),
    .B2(\mul_output.bitseq[6] ),
    .A2(_0264_),
    .A1(\mul_avg[7] ));
 sg13g2_nand2_1 _0972_ (.Y(_0286_),
    .A(\mul_output.bitseq[7] ),
    .B(_0271_));
 sg13g2_nand2_1 _0973_ (.Y(_0034_),
    .A(_0285_),
    .B(_0286_));
 sg13g2_nor2b_1 _0974_ (.A(_0268_),
    .B_N(\mul_output.bitseq[8] ),
    .Y(_0287_));
 sg13g2_a21oi_1 _0975_ (.A1(\mul_output.bitseq[7] ),
    .A2(net30),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_nand2_1 _0976_ (.Y(_0289_),
    .A(\mul_avg[8] ),
    .B(net33));
 sg13g2_o21ai_1 _0977_ (.B1(_0289_),
    .Y(_0035_),
    .A1(net33),
    .A2(_0288_));
 sg13g2_and2_1 _0978_ (.A(\mul_output.bitseq[8] ),
    .B(net30),
    .X(_0036_));
 sg13g2_buf_1 _0979_ (.A(\smul_output.counter[0] ),
    .X(_0290_));
 sg13g2_buf_2 _0980_ (.A(\smul_output.counter[1] ),
    .X(_0291_));
 sg13g2_nor4_2 _0981_ (.A(_0290_),
    .B(_0291_),
    .C(\smul_output.counter[2] ),
    .Y(_0292_),
    .D(\smul_output.counter[3] ));
 sg13g2_buf_1 _0982_ (.A(_0292_),
    .X(_0293_));
 sg13g2_inv_1 _0983_ (.Y(_0294_),
    .A(\smul_output.counter[2] ));
 sg13g2_nand2_1 _0984_ (.Y(_0295_),
    .A(_0294_),
    .B(\smul_output.counter[3] ));
 sg13g2_nand2b_1 _0985_ (.Y(_0296_),
    .B(_0290_),
    .A_N(_0291_));
 sg13g2_nor2_2 _0986_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_buf_1 _0987_ (.A(_0297_),
    .X(_0298_));
 sg13g2_a22oi_1 _0988_ (.Y(_0299_),
    .B1(net29),
    .B2(\smul_output.bitseq[0] ),
    .A2(net32),
    .A1(\smul_avg[1] ));
 sg13g2_nor2_2 _0989_ (.A(_0292_),
    .B(_0297_),
    .Y(_0300_));
 sg13g2_nand2_1 _0990_ (.Y(_0301_),
    .A(\smul_output.bitseq[1] ),
    .B(_0300_));
 sg13g2_nand2_1 _0991_ (.Y(_0037_),
    .A(_0299_),
    .B(_0301_));
 sg13g2_a22oi_1 _0992_ (.Y(_0302_),
    .B1(net29),
    .B2(\smul_output.bitseq[1] ),
    .A2(net32),
    .A1(\smul_avg[2] ));
 sg13g2_nand2_1 _0993_ (.Y(_0303_),
    .A(\smul_output.bitseq[2] ),
    .B(_0300_));
 sg13g2_nand2_1 _0994_ (.Y(_0038_),
    .A(_0302_),
    .B(_0303_));
 sg13g2_a22oi_1 _0995_ (.Y(_0304_),
    .B1(net29),
    .B2(\smul_output.bitseq[2] ),
    .A2(net32),
    .A1(\smul_avg[3] ));
 sg13g2_nand2_1 _0996_ (.Y(_0305_),
    .A(\smul_output.bitseq[3] ),
    .B(_0300_));
 sg13g2_nand2_1 _0997_ (.Y(_0039_),
    .A(_0304_),
    .B(_0305_));
 sg13g2_nor2b_1 _0998_ (.A(_0297_),
    .B_N(\smul_output.bitseq[4] ),
    .Y(_0306_));
 sg13g2_a21oi_1 _0999_ (.A1(\smul_output.bitseq[3] ),
    .A2(net29),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_nand2_1 _1000_ (.Y(_0308_),
    .A(\smul_avg[4] ),
    .B(net32));
 sg13g2_o21ai_1 _1001_ (.B1(_0308_),
    .Y(_0040_),
    .A1(net32),
    .A2(_0307_));
 sg13g2_nor2b_1 _1002_ (.A(_0297_),
    .B_N(\smul_output.bitseq[5] ),
    .Y(_0309_));
 sg13g2_a21oi_1 _1003_ (.A1(\smul_output.bitseq[4] ),
    .A2(net29),
    .Y(_0310_),
    .B1(_0309_));
 sg13g2_nand2_1 _1004_ (.Y(_0311_),
    .A(\smul_avg[5] ),
    .B(net32));
 sg13g2_o21ai_1 _1005_ (.B1(_0311_),
    .Y(_0041_),
    .A1(_0293_),
    .A2(_0310_));
 sg13g2_a22oi_1 _1006_ (.Y(_0312_),
    .B1(net29),
    .B2(\smul_output.bitseq[5] ),
    .A2(_0292_),
    .A1(\smul_avg[6] ));
 sg13g2_nand2_1 _1007_ (.Y(_0313_),
    .A(\smul_output.bitseq[6] ),
    .B(_0300_));
 sg13g2_nand2_1 _1008_ (.Y(_0042_),
    .A(_0312_),
    .B(_0313_));
 sg13g2_a22oi_1 _1009_ (.Y(_0314_),
    .B1(net29),
    .B2(\smul_output.bitseq[6] ),
    .A2(_0292_),
    .A1(\smul_avg[7] ));
 sg13g2_nand2_1 _1010_ (.Y(_0315_),
    .A(\smul_output.bitseq[7] ),
    .B(_0300_));
 sg13g2_nand2_1 _1011_ (.Y(_0043_),
    .A(_0314_),
    .B(_0315_));
 sg13g2_nor2b_1 _1012_ (.A(_0297_),
    .B_N(\smul_output.bitseq[8] ),
    .Y(_0316_));
 sg13g2_a21oi_1 _1013_ (.A1(\smul_output.bitseq[7] ),
    .A2(_0298_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_nand2_1 _1014_ (.Y(_0318_),
    .A(\smul_avg[8] ),
    .B(net32));
 sg13g2_o21ai_1 _1015_ (.B1(_0318_),
    .Y(_0044_),
    .A1(net32),
    .A2(_0317_));
 sg13g2_and2_1 _1016_ (.A(\smul_output.bitseq[8] ),
    .B(net29),
    .X(_0045_));
 sg13g2_buf_2 _1017_ (.A(\add_up_counter.clk_counter[0] ),
    .X(_0319_));
 sg13g2_nor2_1 _1018_ (.A(\add_up_counter.clk_counter[4] ),
    .B(\add_up_counter.clk_counter[6] ),
    .Y(_0320_));
 sg13g2_nor4_1 _1019_ (.A(_0319_),
    .B(\add_up_counter.clk_counter[1] ),
    .C(\add_up_counter.clk_counter[2] ),
    .D(\add_up_counter.clk_counter[3] ),
    .Y(_0321_));
 sg13g2_buf_1 _1020_ (.A(\add_up_counter.clk_counter[9] ),
    .X(_0322_));
 sg13g2_nor4_1 _1021_ (.A(\add_up_counter.clk_counter[5] ),
    .B(\add_up_counter.clk_counter[7] ),
    .C(_0322_),
    .D(\add_up_counter.clk_counter[16] ),
    .Y(_0323_));
 sg13g2_nor4_1 _1022_ (.A(\add_up_counter.clk_counter[8] ),
    .B(\add_up_counter.clk_counter[11] ),
    .C(\add_up_counter.clk_counter[10] ),
    .D(\add_up_counter.clk_counter[13] ),
    .Y(_0324_));
 sg13g2_nand4_1 _1023_ (.B(_0321_),
    .C(_0323_),
    .A(_0320_),
    .Y(_0325_),
    .D(_0324_));
 sg13g2_nor4_2 _1024_ (.A(\add_up_counter.clk_counter[12] ),
    .B(\add_up_counter.clk_counter[15] ),
    .C(\add_up_counter.clk_counter[14] ),
    .Y(_0326_),
    .D(_0325_));
 sg13g2_and2_1 _1025_ (.A(\add_up_counter.clk_counter[17] ),
    .B(_0326_),
    .X(_0327_));
 sg13g2_buf_1 _1026_ (.A(_0327_),
    .X(_0328_));
 sg13g2_buf_1 _1027_ (.A(_0328_),
    .X(_0329_));
 sg13g2_buf_1 _1028_ (.A(net23),
    .X(_0330_));
 sg13g2_nor2_1 _1029_ (.A(_0319_),
    .B(net18),
    .Y(_0000_));
 sg13g2_xor2_1 _1030_ (.B(\add_up_counter.clk_counter[1] ),
    .A(_0319_),
    .X(_0009_));
 sg13g2_nand2_1 _1031_ (.Y(_0331_),
    .A(_0319_),
    .B(\add_up_counter.clk_counter[1] ));
 sg13g2_xnor2_1 _1032_ (.Y(_0010_),
    .A(\add_up_counter.clk_counter[2] ),
    .B(_0331_));
 sg13g2_nand3_1 _1033_ (.B(\add_up_counter.clk_counter[1] ),
    .C(\add_up_counter.clk_counter[2] ),
    .A(_0319_),
    .Y(_0332_));
 sg13g2_xnor2_1 _1034_ (.Y(_0011_),
    .A(\add_up_counter.clk_counter[3] ),
    .B(_0332_));
 sg13g2_inv_1 _1035_ (.Y(_0333_),
    .A(\add_up_counter.clk_counter[3] ));
 sg13g2_nor2_1 _1036_ (.A(_0333_),
    .B(_0332_),
    .Y(_0334_));
 sg13g2_xor2_1 _1037_ (.B(_0334_),
    .A(\add_up_counter.clk_counter[4] ),
    .X(_0012_));
 sg13g2_nand2_1 _1038_ (.Y(_0335_),
    .A(\add_up_counter.clk_counter[4] ),
    .B(_0334_));
 sg13g2_xnor2_1 _1039_ (.Y(_0013_),
    .A(\add_up_counter.clk_counter[5] ),
    .B(_0335_));
 sg13g2_and3_1 _1040_ (.X(_0336_),
    .A(\add_up_counter.clk_counter[4] ),
    .B(\add_up_counter.clk_counter[5] ),
    .C(_0334_));
 sg13g2_xor2_1 _1041_ (.B(_0336_),
    .A(\add_up_counter.clk_counter[6] ),
    .X(_0014_));
 sg13g2_nand2_1 _1042_ (.Y(_0337_),
    .A(\add_up_counter.clk_counter[6] ),
    .B(_0336_));
 sg13g2_xnor2_1 _1043_ (.Y(_0015_),
    .A(\add_up_counter.clk_counter[7] ),
    .B(_0337_));
 sg13g2_nand3_1 _1044_ (.B(\add_up_counter.clk_counter[6] ),
    .C(_0336_),
    .A(\add_up_counter.clk_counter[7] ),
    .Y(_0338_));
 sg13g2_xnor2_1 _1045_ (.Y(_0016_),
    .A(\add_up_counter.clk_counter[8] ),
    .B(_0338_));
 sg13g2_inv_1 _1046_ (.Y(_0339_),
    .A(\add_up_counter.clk_counter[8] ));
 sg13g2_nor2_2 _1047_ (.A(_0339_),
    .B(_0338_),
    .Y(_0340_));
 sg13g2_xor2_1 _1048_ (.B(_0340_),
    .A(_0322_),
    .X(_0017_));
 sg13g2_nand2_1 _1049_ (.Y(_0341_),
    .A(_0322_),
    .B(_0340_));
 sg13g2_xnor2_1 _1050_ (.Y(_0001_),
    .A(\add_up_counter.clk_counter[10] ),
    .B(_0341_));
 sg13g2_nand3_1 _1051_ (.B(\add_up_counter.clk_counter[10] ),
    .C(_0340_),
    .A(_0322_),
    .Y(_0342_));
 sg13g2_xnor2_1 _1052_ (.Y(_0002_),
    .A(\add_up_counter.clk_counter[11] ),
    .B(_0342_));
 sg13g2_nand4_1 _1053_ (.B(\add_up_counter.clk_counter[11] ),
    .C(\add_up_counter.clk_counter[10] ),
    .A(_0322_),
    .Y(_0343_),
    .D(_0340_));
 sg13g2_xnor2_1 _1054_ (.Y(_0003_),
    .A(\add_up_counter.clk_counter[12] ),
    .B(_0343_));
 sg13g2_nand4_1 _1055_ (.B(\add_up_counter.clk_counter[11] ),
    .C(\add_up_counter.clk_counter[10] ),
    .A(_0322_),
    .Y(_0344_),
    .D(\add_up_counter.clk_counter[12] ));
 sg13g2_nor3_2 _1056_ (.A(_0339_),
    .B(_0338_),
    .C(_0344_),
    .Y(_0345_));
 sg13g2_xor2_1 _1057_ (.B(_0345_),
    .A(\add_up_counter.clk_counter[13] ),
    .X(_0004_));
 sg13g2_nand2_1 _1058_ (.Y(_0346_),
    .A(\add_up_counter.clk_counter[13] ),
    .B(_0345_));
 sg13g2_xnor2_1 _1059_ (.Y(_0005_),
    .A(\add_up_counter.clk_counter[14] ),
    .B(_0346_));
 sg13g2_nand3_1 _1060_ (.B(\add_up_counter.clk_counter[14] ),
    .C(_0345_),
    .A(\add_up_counter.clk_counter[13] ),
    .Y(_0347_));
 sg13g2_xnor2_1 _1061_ (.Y(_0006_),
    .A(\add_up_counter.clk_counter[15] ),
    .B(_0347_));
 sg13g2_nand4_1 _1062_ (.B(\add_up_counter.clk_counter[15] ),
    .C(\add_up_counter.clk_counter[14] ),
    .A(\add_up_counter.clk_counter[13] ),
    .Y(_0348_),
    .D(_0345_));
 sg13g2_xnor2_1 _1063_ (.Y(_0007_),
    .A(\add_up_counter.clk_counter[16] ),
    .B(_0348_));
 sg13g2_inv_1 _1064_ (.Y(_0349_),
    .A(\add_up_counter.clk_counter[17] ));
 sg13g2_nor2_1 _1065_ (.A(_0349_),
    .B(_0326_),
    .Y(_0350_));
 sg13g2_inv_1 _1066_ (.Y(_0351_),
    .A(\add_up_counter.clk_counter[16] ));
 sg13g2_nor2_1 _1067_ (.A(_0351_),
    .B(_0348_),
    .Y(_0352_));
 sg13g2_mux2_1 _1068_ (.A0(_0350_),
    .A1(_0349_),
    .S(_0352_),
    .X(_0008_));
 sg13g2_buf_2 _1069_ (.A(\add_output.counter[1] ),
    .X(_0353_));
 sg13g2_buf_1 _1070_ (.A(\add_output.counter[0] ),
    .X(_0354_));
 sg13g2_nor4_2 _1071_ (.A(_0353_),
    .B(_0354_),
    .C(\add_output.counter[2] ),
    .Y(_0355_),
    .D(\add_output.counter[3] ));
 sg13g2_buf_1 _1072_ (.A(_0355_),
    .X(_0356_));
 sg13g2_inv_1 _1073_ (.Y(_0055_),
    .A(_0354_));
 sg13g2_inv_1 _1074_ (.Y(_0357_),
    .A(\add_output.counter[2] ));
 sg13g2_nand2_1 _1075_ (.Y(_0358_),
    .A(_0357_),
    .B(\add_output.counter[3] ));
 sg13g2_nor3_2 _1076_ (.A(_0353_),
    .B(_0055_),
    .C(_0358_),
    .Y(_0359_));
 sg13g2_buf_1 _1077_ (.A(_0359_),
    .X(_0360_));
 sg13g2_a22oi_1 _1078_ (.Y(_0361_),
    .B1(net28),
    .B2(\add_output.bitseq[0] ),
    .A2(net31),
    .A1(\add_avg[1] ));
 sg13g2_nor2_2 _1079_ (.A(_0355_),
    .B(_0359_),
    .Y(_0362_));
 sg13g2_nand2_1 _1080_ (.Y(_0363_),
    .A(\add_output.bitseq[1] ),
    .B(_0362_));
 sg13g2_nand2_1 _1081_ (.Y(_0018_),
    .A(_0361_),
    .B(_0363_));
 sg13g2_a22oi_1 _1082_ (.Y(_0364_),
    .B1(net28),
    .B2(\add_output.bitseq[1] ),
    .A2(net31),
    .A1(\add_avg[2] ));
 sg13g2_nand2_1 _1083_ (.Y(_0365_),
    .A(\add_output.bitseq[2] ),
    .B(_0362_));
 sg13g2_nand2_1 _1084_ (.Y(_0019_),
    .A(_0364_),
    .B(_0365_));
 sg13g2_a22oi_1 _1085_ (.Y(_0366_),
    .B1(net28),
    .B2(\add_output.bitseq[2] ),
    .A2(net31),
    .A1(\add_avg[3] ));
 sg13g2_nand2_1 _1086_ (.Y(_0367_),
    .A(\add_output.bitseq[3] ),
    .B(_0362_));
 sg13g2_nand2_1 _1087_ (.Y(_0020_),
    .A(_0366_),
    .B(_0367_));
 sg13g2_nor2b_1 _1088_ (.A(_0359_),
    .B_N(\add_output.bitseq[4] ),
    .Y(_0368_));
 sg13g2_a21oi_1 _1089_ (.A1(\add_output.bitseq[3] ),
    .A2(_0360_),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_nand2_1 _1090_ (.Y(_0370_),
    .A(\add_avg[4] ),
    .B(net31));
 sg13g2_o21ai_1 _1091_ (.B1(_0370_),
    .Y(_0021_),
    .A1(net31),
    .A2(_0369_));
 sg13g2_nor2b_1 _1092_ (.A(_0359_),
    .B_N(\add_output.bitseq[5] ),
    .Y(_0371_));
 sg13g2_a21oi_1 _1093_ (.A1(\add_output.bitseq[4] ),
    .A2(net28),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_nand2_1 _1094_ (.Y(_0373_),
    .A(\add_avg[5] ),
    .B(_0356_));
 sg13g2_o21ai_1 _1095_ (.B1(_0373_),
    .Y(_0022_),
    .A1(net31),
    .A2(_0372_));
 sg13g2_a22oi_1 _1096_ (.Y(_0374_),
    .B1(net28),
    .B2(\add_output.bitseq[5] ),
    .A2(_0355_),
    .A1(\add_avg[6] ));
 sg13g2_nand2_1 _1097_ (.Y(_0375_),
    .A(\add_output.bitseq[6] ),
    .B(_0362_));
 sg13g2_nand2_1 _1098_ (.Y(_0023_),
    .A(_0374_),
    .B(_0375_));
 sg13g2_a22oi_1 _1099_ (.Y(_0376_),
    .B1(net28),
    .B2(\add_output.bitseq[6] ),
    .A2(_0355_),
    .A1(\add_avg[7] ));
 sg13g2_nand2_1 _1100_ (.Y(_0377_),
    .A(\add_output.bitseq[7] ),
    .B(_0362_));
 sg13g2_nand2_1 _1101_ (.Y(_0024_),
    .A(_0376_),
    .B(_0377_));
 sg13g2_nor2b_1 _1102_ (.A(_0359_),
    .B_N(\add_output.bitseq[8] ),
    .Y(_0378_));
 sg13g2_a21oi_1 _1103_ (.A1(\add_output.bitseq[7] ),
    .A2(_0360_),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_nand2_1 _1104_ (.Y(_0380_),
    .A(\add_avg[8] ),
    .B(net31));
 sg13g2_o21ai_1 _1105_ (.B1(_0380_),
    .Y(_0025_),
    .A1(_0356_),
    .A2(_0379_));
 sg13g2_and2_1 _1106_ (.A(\add_output.bitseq[8] ),
    .B(net28),
    .X(_0026_));
 sg13g2_inv_1 _1107_ (.Y(_0381_),
    .A(\global_input.loop ));
 sg13g2_buf_1 _1108_ (.A(_0328_),
    .X(_0382_));
 sg13g2_buf_2 _1109_ (.A(net22),
    .X(_0383_));
 sg13g2_xor2_1 _1110_ (.B(_0319_),
    .A(\global_input.adjustment[0] ),
    .X(_0384_));
 sg13g2_xor2_1 _1111_ (.B(\add_up_counter.clk_counter[4] ),
    .A(\global_input.adjustment[4] ),
    .X(_0385_));
 sg13g2_xor2_1 _1112_ (.B(\add_up_counter.clk_counter[3] ),
    .A(\global_input.adjustment[3] ),
    .X(_0386_));
 sg13g2_xor2_1 _1113_ (.B(\add_up_counter.clk_counter[1] ),
    .A(\global_input.adjustment[1] ),
    .X(_0387_));
 sg13g2_nor4_1 _1114_ (.A(_0384_),
    .B(_0385_),
    .C(_0386_),
    .D(_0387_),
    .Y(_0388_));
 sg13g2_xnor2_1 _1115_ (.Y(_0389_),
    .A(\global_input.adjustment[2] ),
    .B(\add_up_counter.clk_counter[2] ));
 sg13g2_nand3_1 _1116_ (.B(_0388_),
    .C(_0389_),
    .A(_0381_),
    .Y(_0390_));
 sg13g2_buf_1 _1117_ (.A(_0390_),
    .X(_0391_));
 sg13g2_buf_1 _1118_ (.A(net27),
    .X(_0392_));
 sg13g2_o21ai_1 _1119_ (.B1(net26),
    .Y(_0027_),
    .A1(_0381_),
    .A2(net17));
 sg13g2_inv_1 _1120_ (.Y(_0049_),
    .A(net1));
 sg13g2_nand2_1 _1121_ (.Y(_0393_),
    .A(_0354_),
    .B(_0358_));
 sg13g2_nand2_1 _1122_ (.Y(_0394_),
    .A(_0353_),
    .B(_0055_));
 sg13g2_o21ai_1 _1123_ (.B1(_0394_),
    .Y(_0056_),
    .A1(_0353_),
    .A2(_0393_));
 sg13g2_nand2_1 _1124_ (.Y(_0395_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_xnor2_1 _1125_ (.Y(_0057_),
    .A(\add_output.counter[2] ),
    .B(_0395_));
 sg13g2_o21ai_1 _1126_ (.B1(_0354_),
    .Y(_0396_),
    .A1(_0353_),
    .A2(_0357_));
 sg13g2_nand2_1 _1127_ (.Y(_0397_),
    .A(_0354_),
    .B(\add_output.counter[2] ));
 sg13g2_o21ai_1 _1128_ (.B1(_0358_),
    .Y(_0398_),
    .A1(\add_output.counter[3] ),
    .A2(_0397_));
 sg13g2_a22oi_1 _1129_ (.Y(_0399_),
    .B1(_0398_),
    .B2(_0353_),
    .A2(_0396_),
    .A1(\add_output.counter[3] ));
 sg13g2_inv_1 _1130_ (.Y(_0058_),
    .A(_0399_));
 sg13g2_nand2_1 _1131_ (.Y(_0400_),
    .A(\add_avg[0] ),
    .B(net31));
 sg13g2_nand2b_1 _1132_ (.Y(_0401_),
    .B(\add_output.bitseq[0] ),
    .A_N(_0355_));
 sg13g2_a21oi_1 _1133_ (.A1(_0400_),
    .A2(_0401_),
    .Y(_0059_),
    .B1(net28));
 sg13g2_buf_8 _1134_ (.A(\add_up_counter.prob_counter[0] ),
    .X(_0402_));
 sg13g2_o21ai_1 _1135_ (.B1(\global_SN_gen.lfsr[3] ),
    .Y(_0403_),
    .A1(_0259_),
    .A2(_0260_));
 sg13g2_xnor2_1 _1136_ (.Y(_0404_),
    .A(\global_SN_gen.lfsr[19] ),
    .B(\global_SN_gen.Input_2[7] ));
 sg13g2_inv_1 _1137_ (.Y(_0405_),
    .A(\global_SN_gen.lfsr[18] ));
 sg13g2_xor2_1 _1138_ (.B(\global_SN_gen.Input_2[8] ),
    .A(\global_SN_gen.lfsr[20] ),
    .X(_0406_));
 sg13g2_a21oi_1 _1139_ (.A1(_0405_),
    .A2(\global_SN_gen.Input_2[6] ),
    .Y(_0407_),
    .B1(_0406_));
 sg13g2_nand2b_1 _1140_ (.Y(_0408_),
    .B(\global_SN_gen.lfsr[19] ),
    .A_N(\global_SN_gen.Input_2[7] ));
 sg13g2_nand2_1 _1141_ (.Y(_0409_),
    .A(\global_SN_gen.Input_2[8] ),
    .B(_0408_));
 sg13g2_nor2_1 _1142_ (.A(\global_SN_gen.Input_2[8] ),
    .B(_0408_),
    .Y(_0410_));
 sg13g2_a21o_1 _1143_ (.A2(_0409_),
    .A1(\global_SN_gen.lfsr[20] ),
    .B1(_0410_),
    .X(_0411_));
 sg13g2_a21oi_1 _1144_ (.A1(_0404_),
    .A2(_0407_),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_nor2_1 _1145_ (.A(_0405_),
    .B(\global_SN_gen.Input_2[6] ),
    .Y(_0413_));
 sg13g2_inv_1 _1146_ (.Y(_0414_),
    .A(\global_SN_gen.Input_2[1] ));
 sg13g2_nand2b_1 _1147_ (.Y(_0415_),
    .B(\global_SN_gen.Input_2[0] ),
    .A_N(\global_SN_gen.lfsr[12] ));
 sg13g2_o21ai_1 _1148_ (.B1(_0415_),
    .Y(_0416_),
    .A1(\global_SN_gen.lfsr[13] ),
    .A2(_0414_));
 sg13g2_inv_1 _1149_ (.Y(_0417_),
    .A(\global_SN_gen.Input_2[2] ));
 sg13g2_a22oi_1 _1150_ (.Y(_0418_),
    .B1(_0414_),
    .B2(\global_SN_gen.lfsr[13] ),
    .A2(_0417_),
    .A1(\global_SN_gen.lfsr[14] ));
 sg13g2_xnor2_1 _1151_ (.Y(_0419_),
    .A(\global_SN_gen.lfsr[15] ),
    .B(\global_SN_gen.Input_2[3] ));
 sg13g2_buf_2 _1152_ (.A(\global_SN_gen.lfsr[16] ),
    .X(_0420_));
 sg13g2_xnor2_1 _1153_ (.Y(_0421_),
    .A(_0420_),
    .B(\global_SN_gen.Input_2[4] ));
 sg13g2_nand2b_1 _1154_ (.Y(_0422_),
    .B(\global_SN_gen.Input_2[2] ),
    .A_N(\global_SN_gen.lfsr[14] ));
 sg13g2_xnor2_1 _1155_ (.Y(_0423_),
    .A(\global_SN_gen.lfsr[17] ),
    .B(\global_SN_gen.Input_2[5] ));
 sg13g2_nand4_1 _1156_ (.B(_0421_),
    .C(_0422_),
    .A(_0419_),
    .Y(_0424_),
    .D(_0423_));
 sg13g2_a21oi_1 _1157_ (.A1(_0416_),
    .A2(_0418_),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_nor2_1 _1158_ (.A(\global_SN_gen.Input_2[5] ),
    .B(\global_SN_gen.Input_2[4] ),
    .Y(_0426_));
 sg13g2_nor2b_1 _1159_ (.A(\global_SN_gen.Input_2[5] ),
    .B_N(_0420_),
    .Y(_0427_));
 sg13g2_nor2b_1 _1160_ (.A(\global_SN_gen.Input_2[3] ),
    .B_N(\global_SN_gen.lfsr[15] ),
    .Y(_0428_));
 sg13g2_o21ai_1 _1161_ (.B1(_0428_),
    .Y(_0429_),
    .A1(_0426_),
    .A2(_0427_));
 sg13g2_inv_1 _1162_ (.Y(_0430_),
    .A(\global_SN_gen.Input_2[4] ));
 sg13g2_a21oi_1 _1163_ (.A1(_0430_),
    .A2(_0427_),
    .Y(_0431_),
    .B1(\global_SN_gen.lfsr[17] ));
 sg13g2_o21ai_1 _1164_ (.B1(_0420_),
    .Y(_0432_),
    .A1(_0430_),
    .A2(_0428_));
 sg13g2_inv_1 _1165_ (.Y(_0433_),
    .A(\global_SN_gen.Input_2[5] ));
 sg13g2_a21oi_1 _1166_ (.A1(_0430_),
    .A2(_0428_),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_a22oi_1 _1167_ (.Y(_0435_),
    .B1(_0432_),
    .B2(_0434_),
    .A2(_0431_),
    .A1(_0429_));
 sg13g2_nor4_1 _1168_ (.A(_0411_),
    .B(_0413_),
    .C(_0425_),
    .D(_0435_),
    .Y(_0436_));
 sg13g2_inv_1 _1169_ (.Y(_0437_),
    .A(\global_SN_gen.lfsr[3] ));
 sg13g2_o21ai_1 _1170_ (.B1(_0437_),
    .Y(_0438_),
    .A1(_0412_),
    .A2(_0436_));
 sg13g2_inv_1 _1171_ (.Y(_0439_),
    .A(\add_up_counter.prob_counter[6] ));
 sg13g2_nand3_1 _1172_ (.B(_0402_),
    .C(\add_up_counter.prob_counter[2] ),
    .A(\add_up_counter.prob_counter[1] ),
    .Y(_0440_));
 sg13g2_buf_2 _1173_ (.A(\add_up_counter.prob_counter[3] ),
    .X(_0441_));
 sg13g2_nand3_1 _1174_ (.B(\add_up_counter.prob_counter[5] ),
    .C(\add_up_counter.prob_counter[4] ),
    .A(_0441_),
    .Y(_0442_));
 sg13g2_nor3_2 _1175_ (.A(_0439_),
    .B(_0440_),
    .C(_0442_),
    .Y(_0443_));
 sg13g2_and2_1 _1176_ (.A(\add_up_counter.prob_counter[9] ),
    .B(\add_up_counter.prob_counter[8] ),
    .X(_0444_));
 sg13g2_and4_1 _1177_ (.A(\add_up_counter.prob_counter[7] ),
    .B(\add_up_counter.prob_counter[10] ),
    .C(_0443_),
    .D(_0444_),
    .X(_0445_));
 sg13g2_buf_8 _1178_ (.A(_0445_),
    .X(_0446_));
 sg13g2_and2_1 _1179_ (.A(\add_up_counter.prob_counter[11] ),
    .B(\add_up_counter.prob_counter[12] ),
    .X(_0447_));
 sg13g2_nand4_1 _1180_ (.B(\add_up_counter.prob_counter[14] ),
    .C(_0446_),
    .A(\add_up_counter.prob_counter[13] ),
    .Y(_0448_),
    .D(_0447_));
 sg13g2_nand2_1 _1181_ (.Y(_0449_),
    .A(\add_up_counter.prob_counter[15] ),
    .B(\add_up_counter.prob_counter[16] ));
 sg13g2_nand2_2 _1182_ (.Y(_0450_),
    .A(\add_up_counter.clk_counter[17] ),
    .B(_0326_));
 sg13g2_o21ai_1 _1183_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_a21o_1 _1184_ (.A2(_0438_),
    .A1(_0403_),
    .B1(_0451_),
    .X(_0452_));
 sg13g2_buf_8 _1185_ (.A(_0452_),
    .X(_0453_));
 sg13g2_and3_1 _1186_ (.X(_0454_),
    .A(_0450_),
    .B(_0403_),
    .C(_0438_));
 sg13g2_buf_2 _1187_ (.A(_0454_),
    .X(_0455_));
 sg13g2_nand2_1 _1188_ (.Y(_0456_),
    .A(_0402_),
    .B(_0455_));
 sg13g2_o21ai_1 _1189_ (.B1(_0456_),
    .Y(_0069_),
    .A1(_0402_),
    .A2(_0453_));
 sg13g2_and2_1 _1190_ (.A(_0403_),
    .B(_0438_),
    .X(_0457_));
 sg13g2_buf_2 _1191_ (.A(_0457_),
    .X(_0458_));
 sg13g2_and3_1 _1192_ (.X(_0459_),
    .A(\add_up_counter.prob_counter[7] ),
    .B(_0443_),
    .C(_0444_));
 sg13g2_inv_1 _1193_ (.Y(_0460_),
    .A(_0459_));
 sg13g2_o21ai_1 _1194_ (.B1(\add_up_counter.prob_counter[10] ),
    .Y(_0461_),
    .A1(_0458_),
    .A2(_0460_));
 sg13g2_nand2_1 _1195_ (.Y(_0462_),
    .A(_0403_),
    .B(_0438_));
 sg13g2_nand3b_1 _1196_ (.B(net21),
    .C(_0459_),
    .Y(_0463_),
    .A_N(\add_up_counter.prob_counter[10] ));
 sg13g2_buf_1 _1197_ (.A(_0329_),
    .X(_0464_));
 sg13g2_a21oi_1 _1198_ (.A1(_0461_),
    .A2(_0463_),
    .Y(_0070_),
    .B1(net16));
 sg13g2_inv_1 _1199_ (.Y(_0465_),
    .A(_0446_));
 sg13g2_o21ai_1 _1200_ (.B1(\add_up_counter.prob_counter[11] ),
    .Y(_0466_),
    .A1(_0458_),
    .A2(_0465_));
 sg13g2_nand3b_1 _1201_ (.B(net21),
    .C(_0446_),
    .Y(_0467_),
    .A_N(\add_up_counter.prob_counter[11] ));
 sg13g2_a21oi_1 _1202_ (.A1(_0466_),
    .A2(_0467_),
    .Y(_0071_),
    .B1(net16));
 sg13g2_buf_8 _1203_ (.A(_0451_),
    .X(_0468_));
 sg13g2_nor2_1 _1204_ (.A(\add_up_counter.prob_counter[12] ),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_buf_1 _1205_ (.A(_0450_),
    .X(_0470_));
 sg13g2_and2_1 _1206_ (.A(\add_up_counter.prob_counter[12] ),
    .B(net25),
    .X(_0471_));
 sg13g2_nand3_1 _1207_ (.B(net21),
    .C(_0446_),
    .A(\add_up_counter.prob_counter[11] ),
    .Y(_0472_));
 sg13g2_mux2_1 _1208_ (.A0(_0469_),
    .A1(_0471_),
    .S(_0472_),
    .X(_0072_));
 sg13g2_nand2_1 _1209_ (.Y(_0473_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_o21ai_1 _1210_ (.B1(\add_up_counter.prob_counter[13] ),
    .Y(_0474_),
    .A1(_0458_),
    .A2(_0473_));
 sg13g2_or3_1 _1211_ (.A(\add_up_counter.prob_counter[13] ),
    .B(_0458_),
    .C(_0473_),
    .X(_0475_));
 sg13g2_a21oi_1 _1212_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0073_),
    .B1(net16));
 sg13g2_nand3_1 _1213_ (.B(_0446_),
    .C(_0447_),
    .A(\add_up_counter.prob_counter[13] ),
    .Y(_0476_));
 sg13g2_o21ai_1 _1214_ (.B1(\add_up_counter.prob_counter[14] ),
    .Y(_0477_),
    .A1(_0458_),
    .A2(_0476_));
 sg13g2_inv_1 _1215_ (.Y(_0478_),
    .A(\add_up_counter.prob_counter[14] ));
 sg13g2_nand3b_1 _1216_ (.B(net21),
    .C(_0478_),
    .Y(_0479_),
    .A_N(_0476_));
 sg13g2_a21oi_1 _1217_ (.A1(_0477_),
    .A2(_0479_),
    .Y(_0074_),
    .B1(net16));
 sg13g2_o21ai_1 _1218_ (.B1(\add_up_counter.prob_counter[15] ),
    .Y(_0480_),
    .A1(_0458_),
    .A2(_0448_));
 sg13g2_nor2_1 _1219_ (.A(_0478_),
    .B(_0476_),
    .Y(_0481_));
 sg13g2_nand3b_1 _1220_ (.B(net21),
    .C(_0481_),
    .Y(_0482_),
    .A_N(\add_up_counter.prob_counter[15] ));
 sg13g2_a21oi_1 _1221_ (.A1(_0480_),
    .A2(_0482_),
    .Y(_0075_),
    .B1(_0464_));
 sg13g2_nand2_1 _1222_ (.Y(_0483_),
    .A(\add_up_counter.prob_counter[15] ),
    .B(_0481_));
 sg13g2_o21ai_1 _1223_ (.B1(\add_up_counter.prob_counter[16] ),
    .Y(_0484_),
    .A1(_0458_),
    .A2(_0483_));
 sg13g2_inv_1 _1224_ (.Y(_0485_),
    .A(\add_up_counter.prob_counter[16] ));
 sg13g2_nand4_1 _1225_ (.B(_0485_),
    .C(_0462_),
    .A(\add_up_counter.prob_counter[15] ),
    .Y(_0486_),
    .D(_0481_));
 sg13g2_a21oi_1 _1226_ (.A1(_0484_),
    .A2(_0486_),
    .Y(_0076_),
    .B1(_0464_));
 sg13g2_nand2b_1 _1227_ (.Y(_0487_),
    .B(_0402_),
    .A_N(\add_up_counter.prob_counter[1] ));
 sg13g2_nor2_1 _1228_ (.A(_0402_),
    .B(net15),
    .Y(_0488_));
 sg13g2_o21ai_1 _1229_ (.B1(\add_up_counter.prob_counter[1] ),
    .Y(_0489_),
    .A1(_0455_),
    .A2(_0488_));
 sg13g2_o21ai_1 _1230_ (.B1(_0489_),
    .Y(_0077_),
    .A1(_0453_),
    .A2(_0487_));
 sg13g2_nand2_1 _1231_ (.Y(_0490_),
    .A(\add_up_counter.prob_counter[1] ),
    .B(_0402_));
 sg13g2_nand2_1 _1232_ (.Y(_0491_),
    .A(\add_up_counter.prob_counter[2] ),
    .B(_0490_));
 sg13g2_nor3_1 _1233_ (.A(\add_up_counter.prob_counter[2] ),
    .B(_0490_),
    .C(net15),
    .Y(_0492_));
 sg13g2_a22oi_1 _1234_ (.Y(_0493_),
    .B1(_0492_),
    .B2(net21),
    .A2(_0455_),
    .A1(\add_up_counter.prob_counter[2] ));
 sg13g2_o21ai_1 _1235_ (.B1(_0493_),
    .Y(_0078_),
    .A1(net15),
    .A2(_0491_));
 sg13g2_nor3_1 _1236_ (.A(_0441_),
    .B(_0440_),
    .C(_0453_),
    .Y(_0494_));
 sg13g2_and3_1 _1237_ (.X(_0495_),
    .A(\add_up_counter.prob_counter[1] ),
    .B(_0402_),
    .C(\add_up_counter.prob_counter[2] ));
 sg13g2_buf_1 _1238_ (.A(_0495_),
    .X(_0496_));
 sg13g2_nor2_1 _1239_ (.A(_0496_),
    .B(net15),
    .Y(_0497_));
 sg13g2_o21ai_1 _1240_ (.B1(_0441_),
    .Y(_0498_),
    .A1(_0455_),
    .A2(_0497_));
 sg13g2_nand2b_1 _1241_ (.Y(_0079_),
    .B(_0498_),
    .A_N(_0494_));
 sg13g2_nand3b_1 _1242_ (.B(_0496_),
    .C(_0441_),
    .Y(_0499_),
    .A_N(\add_up_counter.prob_counter[4] ));
 sg13g2_a21oi_1 _1243_ (.A1(_0441_),
    .A2(_0496_),
    .Y(_0500_),
    .B1(net15));
 sg13g2_o21ai_1 _1244_ (.B1(\add_up_counter.prob_counter[4] ),
    .Y(_0501_),
    .A1(_0455_),
    .A2(_0500_));
 sg13g2_o21ai_1 _1245_ (.B1(_0501_),
    .Y(_0080_),
    .A1(_0453_),
    .A2(_0499_));
 sg13g2_nand3_1 _1246_ (.B(\add_up_counter.prob_counter[4] ),
    .C(_0496_),
    .A(_0441_),
    .Y(_0502_));
 sg13g2_nor3_1 _1247_ (.A(\add_up_counter.prob_counter[5] ),
    .B(_0453_),
    .C(_0502_),
    .Y(_0503_));
 sg13g2_nor2b_1 _1248_ (.A(net15),
    .B_N(_0502_),
    .Y(_0504_));
 sg13g2_o21ai_1 _1249_ (.B1(\add_up_counter.prob_counter[5] ),
    .Y(_0505_),
    .A1(_0455_),
    .A2(_0504_));
 sg13g2_nand2b_1 _1250_ (.Y(_0081_),
    .B(_0505_),
    .A_N(_0503_));
 sg13g2_nor2_1 _1251_ (.A(_0440_),
    .B(_0442_),
    .Y(_0506_));
 sg13g2_nand2_1 _1252_ (.Y(_0507_),
    .A(_0439_),
    .B(_0506_));
 sg13g2_nor2_1 _1253_ (.A(_0506_),
    .B(net15),
    .Y(_0508_));
 sg13g2_o21ai_1 _1254_ (.B1(\add_up_counter.prob_counter[6] ),
    .Y(_0509_),
    .A1(_0455_),
    .A2(_0508_));
 sg13g2_o21ai_1 _1255_ (.B1(_0509_),
    .Y(_0082_),
    .A1(_0453_),
    .A2(_0507_));
 sg13g2_a21oi_1 _1256_ (.A1(net21),
    .A2(_0443_),
    .Y(_0510_),
    .B1(net23));
 sg13g2_nand2b_1 _1257_ (.Y(_0511_),
    .B(_0443_),
    .A_N(\add_up_counter.prob_counter[7] ));
 sg13g2_nor2_1 _1258_ (.A(_0453_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_a21o_1 _1259_ (.A2(_0510_),
    .A1(\add_up_counter.prob_counter[7] ),
    .B1(_0512_),
    .X(_0083_));
 sg13g2_and2_1 _1260_ (.A(\add_up_counter.prob_counter[8] ),
    .B(_0470_),
    .X(_0513_));
 sg13g2_nor2_1 _1261_ (.A(\add_up_counter.prob_counter[8] ),
    .B(_0468_),
    .Y(_0514_));
 sg13g2_and3_1 _1262_ (.X(_0515_),
    .A(\add_up_counter.prob_counter[7] ),
    .B(net21),
    .C(_0443_));
 sg13g2_mux2_1 _1263_ (.A0(_0513_),
    .A1(_0514_),
    .S(_0515_),
    .X(_0084_));
 sg13g2_nand3_1 _1264_ (.B(\add_up_counter.prob_counter[8] ),
    .C(_0443_),
    .A(\add_up_counter.prob_counter[7] ),
    .Y(_0516_));
 sg13g2_or2_1 _1265_ (.X(_0517_),
    .B(_0516_),
    .A(\add_up_counter.prob_counter[9] ));
 sg13g2_nor2b_1 _1266_ (.A(net15),
    .B_N(_0516_),
    .Y(_0518_));
 sg13g2_o21ai_1 _1267_ (.B1(\add_up_counter.prob_counter[9] ),
    .Y(_0519_),
    .A1(_0455_),
    .A2(_0518_));
 sg13g2_o21ai_1 _1268_ (.B1(_0519_),
    .Y(_0085_),
    .A1(_0453_),
    .A2(_0517_));
 sg13g2_buf_2 _1269_ (.A(\global_input.output_case[0] ),
    .X(_0520_));
 sg13g2_buf_1 _1270_ (.A(\global_input.output_case[2] ),
    .X(_0521_));
 sg13g2_buf_1 _1271_ (.A(\global_input.output_case[1] ),
    .X(_0522_));
 sg13g2_buf_1 _1272_ (.A(\global_input.output_case[3] ),
    .X(_0523_));
 sg13g2_o21ai_1 _1273_ (.B1(_0523_),
    .Y(_0524_),
    .A1(net37),
    .A2(net36));
 sg13g2_and4_1 _1274_ (.A(_0349_),
    .B(_0046_),
    .C(_0326_),
    .D(_0524_),
    .X(_0525_));
 sg13g2_buf_2 _1275_ (.A(_0525_),
    .X(_0526_));
 sg13g2_mux2_1 _1276_ (.A0(_0047_),
    .A1(_0520_),
    .S(_0526_),
    .X(_0086_));
 sg13g2_nand2_1 _1277_ (.Y(_0527_),
    .A(_0521_),
    .B(net36));
 sg13g2_o21ai_1 _1278_ (.B1(_0520_),
    .Y(_0528_),
    .A1(net37),
    .A2(net36));
 sg13g2_a21oi_1 _1279_ (.A1(_0527_),
    .A2(_0528_),
    .Y(_0529_),
    .B1(_0523_));
 sg13g2_mux2_1 _1280_ (.A0(\global_input.adjustment[1] ),
    .A1(_0529_),
    .S(_0526_),
    .X(_0087_));
 sg13g2_nand2b_1 _1281_ (.Y(_0530_),
    .B(_0520_),
    .A_N(\global_input.output_case[1] ));
 sg13g2_xnor2_1 _1282_ (.Y(_0531_),
    .A(net37),
    .B(_0523_));
 sg13g2_inv_1 _1283_ (.Y(_0532_),
    .A(_0523_));
 sg13g2_nor2_1 _1284_ (.A(net37),
    .B(_0520_),
    .Y(_0533_));
 sg13g2_nand3_1 _1285_ (.B(net36),
    .C(_0533_),
    .A(_0532_),
    .Y(_0534_));
 sg13g2_o21ai_1 _1286_ (.B1(_0534_),
    .Y(_0535_),
    .A1(_0530_),
    .A2(_0531_));
 sg13g2_mux2_1 _1287_ (.A0(\global_input.adjustment[2] ),
    .A1(_0535_),
    .S(_0526_),
    .X(_0088_));
 sg13g2_inv_1 _1288_ (.Y(_0536_),
    .A(_0048_));
 sg13g2_nor2_1 _1289_ (.A(_0532_),
    .B(_0522_),
    .Y(_0537_));
 sg13g2_nand2b_1 _1290_ (.Y(_0538_),
    .B(_0522_),
    .A_N(_0520_));
 sg13g2_nand3_1 _1291_ (.B(_0530_),
    .C(_0538_),
    .A(net37),
    .Y(_0539_));
 sg13g2_o21ai_1 _1292_ (.B1(_0539_),
    .Y(_0540_),
    .A1(net37),
    .A2(_0530_));
 sg13g2_a22oi_1 _1293_ (.Y(_0541_),
    .B1(_0540_),
    .B2(_0532_),
    .A2(_0537_),
    .A1(_0533_));
 sg13g2_nand2b_1 _1294_ (.Y(_0542_),
    .B(_0526_),
    .A_N(_0541_));
 sg13g2_o21ai_1 _1295_ (.B1(_0542_),
    .Y(_0089_),
    .A1(_0536_),
    .A2(_0526_));
 sg13g2_inv_1 _1296_ (.Y(_0543_),
    .A(\global_input.adjustment[4] ));
 sg13g2_o21ai_1 _1297_ (.B1(_0542_),
    .Y(_0090_),
    .A1(_0543_),
    .A2(_0526_));
 sg13g2_mux2_1 _1298_ (.A0(\global_input.output_bitcounter_1[0] ),
    .A1(\global_SN_gen.Input_1[0] ),
    .S(net26),
    .X(_0109_));
 sg13g2_mux2_1 _1299_ (.A0(\global_input.output_bitcounter_1[1] ),
    .A1(\global_SN_gen.Input_1[1] ),
    .S(net26),
    .X(_0110_));
 sg13g2_mux2_1 _1300_ (.A0(\global_input.output_bitcounter_1[2] ),
    .A1(\global_SN_gen.Input_1[2] ),
    .S(net26),
    .X(_0111_));
 sg13g2_mux2_1 _1301_ (.A0(\global_input.output_bitcounter_1[3] ),
    .A1(_0238_),
    .S(_0392_),
    .X(_0112_));
 sg13g2_mux2_1 _1302_ (.A0(\global_input.output_bitcounter_1[4] ),
    .A1(\global_SN_gen.Input_1[4] ),
    .S(_0392_),
    .X(_0113_));
 sg13g2_mux2_1 _1303_ (.A0(\global_input.output_bitcounter_1[5] ),
    .A1(\global_SN_gen.Input_1[5] ),
    .S(net26),
    .X(_0114_));
 sg13g2_mux2_1 _1304_ (.A0(\global_input.output_bitcounter_1[6] ),
    .A1(\global_SN_gen.Input_1[6] ),
    .S(net26),
    .X(_0115_));
 sg13g2_mux2_1 _1305_ (.A0(\global_input.output_bitcounter_1[7] ),
    .A1(\global_SN_gen.Input_1[7] ),
    .S(net26),
    .X(_0116_));
 sg13g2_mux2_1 _1306_ (.A0(\global_input.output_bitcounter_1[8] ),
    .A1(\global_SN_gen.Input_1[8] ),
    .S(net26),
    .X(_0117_));
 sg13g2_mux2_1 _1307_ (.A0(\global_input.output_bitcounter_2[0] ),
    .A1(\global_SN_gen.Input_2[0] ),
    .S(_0391_),
    .X(_0118_));
 sg13g2_mux2_1 _1308_ (.A0(\global_input.output_bitcounter_2[1] ),
    .A1(\global_SN_gen.Input_2[1] ),
    .S(_0391_),
    .X(_0119_));
 sg13g2_mux2_1 _1309_ (.A0(\global_input.output_bitcounter_2[2] ),
    .A1(\global_SN_gen.Input_2[2] ),
    .S(net27),
    .X(_0120_));
 sg13g2_mux2_1 _1310_ (.A0(\global_input.output_bitcounter_2[3] ),
    .A1(\global_SN_gen.Input_2[3] ),
    .S(net27),
    .X(_0121_));
 sg13g2_mux2_1 _1311_ (.A0(\global_input.output_bitcounter_2[4] ),
    .A1(\global_SN_gen.Input_2[4] ),
    .S(net27),
    .X(_0122_));
 sg13g2_mux2_1 _1312_ (.A0(\global_input.output_bitcounter_2[5] ),
    .A1(\global_SN_gen.Input_2[5] ),
    .S(net27),
    .X(_0123_));
 sg13g2_mux2_1 _1313_ (.A0(\global_input.output_bitcounter_2[6] ),
    .A1(\global_SN_gen.Input_2[6] ),
    .S(net27),
    .X(_0124_));
 sg13g2_mux2_1 _1314_ (.A0(\global_input.output_bitcounter_2[7] ),
    .A1(\global_SN_gen.Input_2[7] ),
    .S(net27),
    .X(_0125_));
 sg13g2_mux2_1 _1315_ (.A0(\global_input.output_bitcounter_2[8] ),
    .A1(\global_SN_gen.Input_2[8] ),
    .S(net27),
    .X(_0126_));
 sg13g2_buf_1 _1316_ (.A(\global_input.loop ),
    .X(_0544_));
 sg13g2_nand2_1 _1317_ (.Y(_0545_),
    .A(net35),
    .B(_0329_));
 sg13g2_xnor2_1 _1318_ (.Y(_0127_),
    .A(_0520_),
    .B(_0545_));
 sg13g2_inv_1 _1319_ (.Y(_0546_),
    .A(net37));
 sg13g2_a21oi_1 _1320_ (.A1(_0546_),
    .A2(_0523_),
    .Y(_0547_),
    .B1(net36));
 sg13g2_nand3_1 _1321_ (.B(_0520_),
    .C(net22),
    .A(\global_input.loop ),
    .Y(_0548_));
 sg13g2_mux2_1 _1322_ (.A0(_0547_),
    .A1(net36),
    .S(_0548_),
    .X(_0128_));
 sg13g2_nand4_1 _1323_ (.B(net36),
    .C(_0520_),
    .A(\global_input.loop ),
    .Y(_0549_),
    .D(_0328_));
 sg13g2_xnor2_1 _1324_ (.Y(_0129_),
    .A(net37),
    .B(_0549_));
 sg13g2_a21oi_1 _1325_ (.A1(_0546_),
    .A2(net36),
    .Y(_0550_),
    .B1(_0548_));
 sg13g2_nor2_1 _1326_ (.A(_0523_),
    .B(_0549_),
    .Y(_0551_));
 sg13g2_o21ai_1 _1327_ (.B1(_0521_),
    .Y(_0552_),
    .A1(_0537_),
    .A2(_0551_));
 sg13g2_o21ai_1 _1328_ (.B1(_0552_),
    .Y(_0130_),
    .A1(_0532_),
    .A2(_0550_));
 sg13g2_nand2_1 _1329_ (.Y(_0553_),
    .A(_0263_),
    .B(_0267_));
 sg13g2_nand2_1 _1330_ (.Y(_0554_),
    .A(_0262_),
    .B(_0131_));
 sg13g2_o21ai_1 _1331_ (.B1(_0554_),
    .Y(_0132_),
    .A1(_0262_),
    .A2(_0553_));
 sg13g2_nand2_1 _1332_ (.Y(_0555_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xnor2_1 _1333_ (.Y(_0133_),
    .A(\mul_output.counter[2] ),
    .B(_0555_));
 sg13g2_o21ai_1 _1334_ (.B1(_0263_),
    .Y(_0556_),
    .A1(_0262_),
    .A2(_0266_));
 sg13g2_nand2_1 _1335_ (.Y(_0557_),
    .A(_0263_),
    .B(\mul_output.counter[2] ));
 sg13g2_o21ai_1 _1336_ (.B1(_0267_),
    .Y(_0558_),
    .A1(\mul_output.counter[3] ),
    .A2(_0557_));
 sg13g2_a22oi_1 _1337_ (.Y(_0559_),
    .B1(_0558_),
    .B2(_0262_),
    .A2(_0556_),
    .A1(\mul_output.counter[3] ));
 sg13g2_inv_1 _1338_ (.Y(_0134_),
    .A(_0559_));
 sg13g2_nand2_1 _1339_ (.Y(_0560_),
    .A(\mul_avg[0] ),
    .B(net33));
 sg13g2_nand2b_1 _1340_ (.Y(_0561_),
    .B(\mul_output.bitseq[0] ),
    .A_N(_0264_));
 sg13g2_a21oi_1 _1341_ (.A1(_0560_),
    .A2(_0561_),
    .Y(_0135_),
    .B1(net30));
 sg13g2_and3_1 _1342_ (.X(_0562_),
    .A(\mul_up_counter.prob_counter[1] ),
    .B(\mul_up_counter.prob_counter[0] ),
    .C(\mul_up_counter.prob_counter[2] ));
 sg13g2_and4_1 _1343_ (.A(\mul_up_counter.prob_counter[3] ),
    .B(\mul_up_counter.prob_counter[5] ),
    .C(\mul_up_counter.prob_counter[4] ),
    .D(_0562_),
    .X(_0563_));
 sg13g2_buf_1 _1344_ (.A(_0563_),
    .X(_0564_));
 sg13g2_and3_1 _1345_ (.X(_0565_),
    .A(\mul_up_counter.prob_counter[7] ),
    .B(\mul_up_counter.prob_counter[6] ),
    .C(_0564_));
 sg13g2_and2_1 _1346_ (.A(\mul_up_counter.prob_counter[9] ),
    .B(\mul_up_counter.prob_counter[8] ),
    .X(_0566_));
 sg13g2_buf_1 _1347_ (.A(\mul_up_counter.prob_counter[11] ),
    .X(_0567_));
 sg13g2_and2_1 _1348_ (.A(_0567_),
    .B(\mul_up_counter.prob_counter[12] ),
    .X(_0568_));
 sg13g2_and4_1 _1349_ (.A(\mul_up_counter.prob_counter[10] ),
    .B(_0565_),
    .C(_0566_),
    .D(_0568_),
    .X(_0569_));
 sg13g2_and4_1 _1350_ (.A(\mul_up_counter.prob_counter[13] ),
    .B(\mul_up_counter.prob_counter[15] ),
    .C(\mul_up_counter.prob_counter[14] ),
    .D(_0569_),
    .X(_0570_));
 sg13g2_a21oi_1 _1351_ (.A1(\mul_up_counter.prob_counter[16] ),
    .A2(_0570_),
    .Y(_0571_),
    .B1(_0328_));
 sg13g2_nor2_1 _1352_ (.A(_0412_),
    .B(_0436_),
    .Y(_0572_));
 sg13g2_xnor2_1 _1353_ (.Y(_0573_),
    .A(_0261_),
    .B(_0572_));
 sg13g2_buf_1 _1354_ (.A(_0573_),
    .X(_0574_));
 sg13g2_buf_1 _1355_ (.A(net14),
    .X(_0575_));
 sg13g2_nand2_1 _1356_ (.Y(_0576_),
    .A(net20),
    .B(net10));
 sg13g2_buf_1 _1357_ (.A(net14),
    .X(_0577_));
 sg13g2_nand3b_1 _1358_ (.B(\mul_up_counter.prob_counter[0] ),
    .C(net25),
    .Y(_0578_),
    .A_N(net9));
 sg13g2_o21ai_1 _1359_ (.B1(_0578_),
    .Y(_0145_),
    .A1(\mul_up_counter.prob_counter[0] ),
    .A2(_0576_));
 sg13g2_buf_1 _1360_ (.A(net22),
    .X(_0579_));
 sg13g2_nor2_1 _1361_ (.A(\mul_up_counter.prob_counter[10] ),
    .B(net13),
    .Y(_0580_));
 sg13g2_inv_1 _1362_ (.Y(_0581_),
    .A(\mul_up_counter.prob_counter[10] ));
 sg13g2_nor2_1 _1363_ (.A(_0581_),
    .B(net23),
    .Y(_0582_));
 sg13g2_and2_1 _1364_ (.A(\mul_up_counter.prob_counter[8] ),
    .B(_0565_),
    .X(_0583_));
 sg13g2_nand3_1 _1365_ (.B(_0574_),
    .C(_0583_),
    .A(\mul_up_counter.prob_counter[9] ),
    .Y(_0584_));
 sg13g2_mux2_1 _1366_ (.A0(_0580_),
    .A1(_0582_),
    .S(_0584_),
    .X(_0146_));
 sg13g2_nand2_1 _1367_ (.Y(_0585_),
    .A(\mul_up_counter.prob_counter[6] ),
    .B(_0564_));
 sg13g2_nand4_1 _1368_ (.B(\mul_up_counter.prob_counter[9] ),
    .C(\mul_up_counter.prob_counter[8] ),
    .A(\mul_up_counter.prob_counter[7] ),
    .Y(_0586_),
    .D(\mul_up_counter.prob_counter[10] ));
 sg13g2_nor2_2 _1369_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_nand2_1 _1370_ (.Y(_0588_),
    .A(_0567_),
    .B(_0450_));
 sg13g2_a21oi_1 _1371_ (.A1(net10),
    .A2(_0587_),
    .Y(_0589_),
    .B1(_0588_));
 sg13g2_nor2_1 _1372_ (.A(_0567_),
    .B(net22),
    .Y(_0590_));
 sg13g2_nand3_1 _1373_ (.B(_0587_),
    .C(_0590_),
    .A(net10),
    .Y(_0591_));
 sg13g2_nand2b_1 _1374_ (.Y(_0147_),
    .B(_0591_),
    .A_N(_0589_));
 sg13g2_nor2_1 _1375_ (.A(\mul_up_counter.prob_counter[12] ),
    .B(net13),
    .Y(_0592_));
 sg13g2_and2_1 _1376_ (.A(\mul_up_counter.prob_counter[12] ),
    .B(net25),
    .X(_0593_));
 sg13g2_nand3_1 _1377_ (.B(net14),
    .C(_0587_),
    .A(_0567_),
    .Y(_0594_));
 sg13g2_mux2_1 _1378_ (.A0(_0592_),
    .A1(_0593_),
    .S(_0594_),
    .X(_0148_));
 sg13g2_nor2_1 _1379_ (.A(\mul_up_counter.prob_counter[13] ),
    .B(net13),
    .Y(_0595_));
 sg13g2_inv_1 _1380_ (.Y(_0596_),
    .A(\mul_up_counter.prob_counter[13] ));
 sg13g2_nor2_1 _1381_ (.A(_0596_),
    .B(net23),
    .Y(_0597_));
 sg13g2_nand4_1 _1382_ (.B(\mul_up_counter.prob_counter[12] ),
    .C(net14),
    .A(_0567_),
    .Y(_0598_),
    .D(_0587_));
 sg13g2_mux2_1 _1383_ (.A0(_0595_),
    .A1(_0597_),
    .S(_0598_),
    .X(_0149_));
 sg13g2_and4_1 _1384_ (.A(_0567_),
    .B(\mul_up_counter.prob_counter[13] ),
    .C(\mul_up_counter.prob_counter[12] ),
    .D(_0587_),
    .X(_0599_));
 sg13g2_buf_1 _1385_ (.A(_0599_),
    .X(_0600_));
 sg13g2_nand2_1 _1386_ (.Y(_0601_),
    .A(\mul_up_counter.prob_counter[14] ),
    .B(_0450_));
 sg13g2_a21oi_1 _1387_ (.A1(net10),
    .A2(_0600_),
    .Y(_0602_),
    .B1(_0601_));
 sg13g2_nor2_1 _1388_ (.A(\mul_up_counter.prob_counter[14] ),
    .B(net22),
    .Y(_0603_));
 sg13g2_nand3_1 _1389_ (.B(_0600_),
    .C(_0603_),
    .A(_0575_),
    .Y(_0604_));
 sg13g2_nand2b_1 _1390_ (.Y(_0150_),
    .B(_0604_),
    .A_N(_0602_));
 sg13g2_nor2_1 _1391_ (.A(\mul_up_counter.prob_counter[15] ),
    .B(net13),
    .Y(_0605_));
 sg13g2_and2_1 _1392_ (.A(\mul_up_counter.prob_counter[15] ),
    .B(net25),
    .X(_0606_));
 sg13g2_nand3_1 _1393_ (.B(net14),
    .C(_0600_),
    .A(\mul_up_counter.prob_counter[14] ),
    .Y(_0607_));
 sg13g2_mux2_1 _1394_ (.A0(_0605_),
    .A1(_0606_),
    .S(_0607_),
    .X(_0151_));
 sg13g2_nor2_1 _1395_ (.A(\mul_up_counter.prob_counter[16] ),
    .B(net13),
    .Y(_0608_));
 sg13g2_and2_1 _1396_ (.A(\mul_up_counter.prob_counter[16] ),
    .B(net25),
    .X(_0609_));
 sg13g2_nand4_1 _1397_ (.B(\mul_up_counter.prob_counter[14] ),
    .C(net14),
    .A(\mul_up_counter.prob_counter[15] ),
    .Y(_0610_),
    .D(_0600_));
 sg13g2_mux2_1 _1398_ (.A0(_0608_),
    .A1(_0609_),
    .S(_0610_),
    .X(_0152_));
 sg13g2_inv_1 _1399_ (.Y(_0611_),
    .A(\mul_up_counter.prob_counter[1] ));
 sg13g2_a21o_1 _1400_ (.A2(net9),
    .A1(\mul_up_counter.prob_counter[0] ),
    .B1(net23),
    .X(_0612_));
 sg13g2_nand4_1 _1401_ (.B(\mul_up_counter.prob_counter[0] ),
    .C(net20),
    .A(_0611_),
    .Y(_0613_),
    .D(net10));
 sg13g2_o21ai_1 _1402_ (.B1(_0613_),
    .Y(_0153_),
    .A1(_0611_),
    .A2(_0612_));
 sg13g2_and2_1 _1403_ (.A(\mul_up_counter.prob_counter[1] ),
    .B(\mul_up_counter.prob_counter[0] ),
    .X(_0614_));
 sg13g2_nand3_1 _1404_ (.B(net20),
    .C(net9),
    .A(_0614_),
    .Y(_0615_));
 sg13g2_nand2_1 _1405_ (.Y(_0616_),
    .A(\mul_up_counter.prob_counter[2] ),
    .B(_0450_));
 sg13g2_a21o_1 _1406_ (.A2(net9),
    .A1(_0614_),
    .B1(_0616_),
    .X(_0617_));
 sg13g2_o21ai_1 _1407_ (.B1(_0617_),
    .Y(_0154_),
    .A1(\mul_up_counter.prob_counter[2] ),
    .A2(_0615_));
 sg13g2_inv_1 _1408_ (.Y(_0618_),
    .A(\mul_up_counter.prob_counter[3] ));
 sg13g2_a21o_1 _1409_ (.A2(net9),
    .A1(_0562_),
    .B1(net23),
    .X(_0619_));
 sg13g2_nand4_1 _1410_ (.B(_0562_),
    .C(net20),
    .A(_0618_),
    .Y(_0620_),
    .D(net10));
 sg13g2_o21ai_1 _1411_ (.B1(_0620_),
    .Y(_0155_),
    .A1(_0618_),
    .A2(_0619_));
 sg13g2_inv_1 _1412_ (.Y(_0621_),
    .A(\mul_up_counter.prob_counter[4] ));
 sg13g2_and2_1 _1413_ (.A(\mul_up_counter.prob_counter[3] ),
    .B(_0562_),
    .X(_0622_));
 sg13g2_a21o_1 _1414_ (.A2(_0622_),
    .A1(net9),
    .B1(net23),
    .X(_0623_));
 sg13g2_nand4_1 _1415_ (.B(net20),
    .C(net10),
    .A(_0621_),
    .Y(_0624_),
    .D(_0622_));
 sg13g2_o21ai_1 _1416_ (.B1(_0624_),
    .Y(_0156_),
    .A1(_0621_),
    .A2(_0623_));
 sg13g2_inv_1 _1417_ (.Y(_0625_),
    .A(\mul_up_counter.prob_counter[5] ));
 sg13g2_and2_1 _1418_ (.A(\mul_up_counter.prob_counter[4] ),
    .B(_0622_),
    .X(_0626_));
 sg13g2_a21o_1 _1419_ (.A2(_0626_),
    .A1(net9),
    .B1(net22),
    .X(_0627_));
 sg13g2_nand4_1 _1420_ (.B(net20),
    .C(_0575_),
    .A(_0625_),
    .Y(_0628_),
    .D(_0626_));
 sg13g2_o21ai_1 _1421_ (.B1(_0628_),
    .Y(_0157_),
    .A1(_0625_),
    .A2(_0627_));
 sg13g2_inv_1 _1422_ (.Y(_0629_),
    .A(\mul_up_counter.prob_counter[6] ));
 sg13g2_a21o_1 _1423_ (.A2(_0577_),
    .A1(_0564_),
    .B1(net22),
    .X(_0630_));
 sg13g2_nand4_1 _1424_ (.B(_0564_),
    .C(_0571_),
    .A(_0629_),
    .Y(_0631_),
    .D(net10));
 sg13g2_o21ai_1 _1425_ (.B1(_0631_),
    .Y(_0158_),
    .A1(_0629_),
    .A2(_0630_));
 sg13g2_nor2_1 _1426_ (.A(\mul_up_counter.prob_counter[7] ),
    .B(net13),
    .Y(_0632_));
 sg13g2_and2_1 _1427_ (.A(\mul_up_counter.prob_counter[7] ),
    .B(net25),
    .X(_0633_));
 sg13g2_nand3_1 _1428_ (.B(_0564_),
    .C(net14),
    .A(\mul_up_counter.prob_counter[6] ),
    .Y(_0634_));
 sg13g2_mux2_1 _1429_ (.A0(_0632_),
    .A1(_0633_),
    .S(_0634_),
    .X(_0159_));
 sg13g2_inv_1 _1430_ (.Y(_0635_),
    .A(\mul_up_counter.prob_counter[8] ));
 sg13g2_a21o_1 _1431_ (.A2(_0574_),
    .A1(_0565_),
    .B1(_0382_),
    .X(_0636_));
 sg13g2_nand4_1 _1432_ (.B(_0565_),
    .C(net20),
    .A(_0635_),
    .Y(_0637_),
    .D(net9));
 sg13g2_o21ai_1 _1433_ (.B1(_0637_),
    .Y(_0160_),
    .A1(_0635_),
    .A2(_0636_));
 sg13g2_and3_1 _1434_ (.X(_0638_),
    .A(net20),
    .B(net14),
    .C(_0583_));
 sg13g2_a21oi_1 _1435_ (.A1(_0577_),
    .A2(_0583_),
    .Y(_0639_),
    .B1(net23));
 sg13g2_mux2_1 _1436_ (.A0(_0638_),
    .A1(_0639_),
    .S(\mul_up_counter.prob_counter[9] ),
    .X(_0161_));
 sg13g2_inv_1 _1437_ (.Y(_0162_),
    .A(_0290_));
 sg13g2_a21oi_1 _1438_ (.A1(_0294_),
    .A2(\smul_output.counter[3] ),
    .Y(_0640_),
    .B1(_0296_));
 sg13g2_a21o_1 _1439_ (.A2(_0291_),
    .A1(_0162_),
    .B1(_0640_),
    .X(_0163_));
 sg13g2_nand2_1 _1440_ (.Y(_0641_),
    .A(_0290_),
    .B(_0291_));
 sg13g2_xnor2_1 _1441_ (.Y(_0164_),
    .A(\smul_output.counter[2] ),
    .B(_0641_));
 sg13g2_o21ai_1 _1442_ (.B1(_0290_),
    .Y(_0642_),
    .A1(_0291_),
    .A2(_0294_));
 sg13g2_nand2_1 _1443_ (.Y(_0643_),
    .A(_0290_),
    .B(\smul_output.counter[2] ));
 sg13g2_o21ai_1 _1444_ (.B1(_0295_),
    .Y(_0644_),
    .A1(\smul_output.counter[3] ),
    .A2(_0643_));
 sg13g2_a22oi_1 _1445_ (.Y(_0645_),
    .B1(_0644_),
    .B2(_0291_),
    .A2(_0642_),
    .A1(\smul_output.counter[3] ));
 sg13g2_inv_1 _1446_ (.Y(_0165_),
    .A(_0645_));
 sg13g2_nand2_1 _1447_ (.Y(_0646_),
    .A(\smul_avg[0] ),
    .B(_0293_));
 sg13g2_nand2b_1 _1448_ (.Y(_0647_),
    .B(\smul_output.bitseq[0] ),
    .A_N(_0292_));
 sg13g2_a21oi_1 _1449_ (.A1(_0646_),
    .A2(_0647_),
    .Y(_0166_),
    .B1(_0298_));
 sg13g2_inv_1 _1450_ (.Y(_0648_),
    .A(\smul.SN_Bit_Q ));
 sg13g2_inv_1 _1451_ (.Y(_0649_),
    .A(\global_SN_gen.Input_1[7] ));
 sg13g2_nor2_1 _1452_ (.A(_0256_),
    .B(\global_SN_gen.lfsr[17] ),
    .Y(_0650_));
 sg13g2_nor2b_1 _1453_ (.A(\global_SN_gen.lfsr[18] ),
    .B_N(\global_SN_gen.Input_1[6] ),
    .Y(_0651_));
 sg13g2_nor2b_1 _1454_ (.A(\global_SN_gen.Input_1[5] ),
    .B_N(\global_SN_gen.lfsr[17] ),
    .Y(_0652_));
 sg13g2_nand2b_1 _1455_ (.Y(_0653_),
    .B(_0238_),
    .A_N(\global_SN_gen.lfsr[15] ));
 sg13g2_nor3_1 _1456_ (.A(_0420_),
    .B(_0652_),
    .C(_0653_),
    .Y(_0654_));
 sg13g2_a221oi_1 _1457_ (.B2(_0653_),
    .C1(_0245_),
    .B1(_0420_),
    .A1(_0256_),
    .Y(_0655_),
    .A2(\global_SN_gen.lfsr[17] ));
 sg13g2_nor4_1 _1458_ (.A(_0650_),
    .B(_0651_),
    .C(_0654_),
    .D(_0655_),
    .Y(_0656_));
 sg13g2_nand2b_1 _1459_ (.Y(_0657_),
    .B(\global_SN_gen.Input_1[0] ),
    .A_N(\global_SN_gen.lfsr[12] ));
 sg13g2_a21oi_1 _1460_ (.A1(_0233_),
    .A2(\global_SN_gen.lfsr[13] ),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_nand2b_1 _1461_ (.Y(_0659_),
    .B(\global_SN_gen.Input_1[2] ),
    .A_N(\global_SN_gen.lfsr[14] ));
 sg13g2_o21ai_1 _1462_ (.B1(_0659_),
    .Y(_0660_),
    .A1(_0233_),
    .A2(\global_SN_gen.lfsr[13] ));
 sg13g2_xor2_1 _1463_ (.B(\global_SN_gen.Input_1[4] ),
    .A(_0420_),
    .X(_0661_));
 sg13g2_nor2b_1 _1464_ (.A(\global_SN_gen.Input_1[2] ),
    .B_N(\global_SN_gen.lfsr[14] ),
    .Y(_0662_));
 sg13g2_xor2_1 _1465_ (.B(\global_SN_gen.lfsr[15] ),
    .A(_0238_),
    .X(_0663_));
 sg13g2_nor4_1 _1466_ (.A(_0652_),
    .B(_0661_),
    .C(_0662_),
    .D(_0663_),
    .Y(_0664_));
 sg13g2_o21ai_1 _1467_ (.B1(_0664_),
    .Y(_0665_),
    .A1(_0658_),
    .A2(_0660_));
 sg13g2_nand2_1 _1468_ (.Y(_0666_),
    .A(_0232_),
    .B(\global_SN_gen.lfsr[20] ));
 sg13g2_o21ai_1 _1469_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_0405_),
    .A2(\global_SN_gen.Input_1[6] ));
 sg13g2_a221oi_1 _1470_ (.B2(_0665_),
    .C1(_0667_),
    .B1(_0656_),
    .A1(\global_SN_gen.lfsr[19] ),
    .Y(_0668_),
    .A2(_0649_));
 sg13g2_nand3b_1 _1471_ (.B(\global_SN_gen.Input_1[7] ),
    .C(_0666_),
    .Y(_0669_),
    .A_N(\global_SN_gen.lfsr[19] ));
 sg13g2_o21ai_1 _1472_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0232_),
    .A2(\global_SN_gen.lfsr[20] ));
 sg13g2_or3_1 _1473_ (.A(_0648_),
    .B(_0668_),
    .C(_0670_),
    .X(_0671_));
 sg13g2_buf_1 _1474_ (.A(_0671_),
    .X(_0672_));
 sg13g2_o21ai_1 _1475_ (.B1(_0648_),
    .Y(_0673_),
    .A1(_0668_),
    .A2(_0670_));
 sg13g2_nand2_1 _1476_ (.Y(_0674_),
    .A(_0672_),
    .B(_0673_));
 sg13g2_buf_1 _1477_ (.A(_0674_),
    .X(_0675_));
 sg13g2_xor2_1 _1478_ (.B(net8),
    .A(\smul_up_counter.prob_counter[0] ),
    .X(_0676_));
 sg13g2_nor2_1 _1479_ (.A(net18),
    .B(_0676_),
    .Y(_0176_));
 sg13g2_buf_1 _1480_ (.A(_0672_),
    .X(_0677_));
 sg13g2_buf_1 _1481_ (.A(_0673_),
    .X(_0678_));
 sg13g2_and4_1 _1482_ (.A(\smul_up_counter.prob_counter[1] ),
    .B(\smul_up_counter.prob_counter[0] ),
    .C(\smul_up_counter.prob_counter[3] ),
    .D(\smul_up_counter.prob_counter[2] ),
    .X(_0679_));
 sg13g2_and4_1 _1483_ (.A(\smul_up_counter.prob_counter[5] ),
    .B(\smul_up_counter.prob_counter[4] ),
    .C(\smul_up_counter.prob_counter[6] ),
    .D(_0679_),
    .X(_0680_));
 sg13g2_and2_1 _1484_ (.A(\smul_up_counter.prob_counter[7] ),
    .B(_0680_),
    .X(_0681_));
 sg13g2_and3_1 _1485_ (.X(_0682_),
    .A(\smul_up_counter.prob_counter[9] ),
    .B(\smul_up_counter.prob_counter[8] ),
    .C(_0681_));
 sg13g2_and3_1 _1486_ (.X(_0683_),
    .A(net12),
    .B(net19),
    .C(_0682_));
 sg13g2_xnor2_1 _1487_ (.Y(_0684_),
    .A(\smul_up_counter.prob_counter[10] ),
    .B(_0683_));
 sg13g2_nor2_1 _1488_ (.A(net18),
    .B(_0684_),
    .Y(_0177_));
 sg13g2_nand4_1 _1489_ (.B(net12),
    .C(net19),
    .A(\smul_up_counter.prob_counter[10] ),
    .Y(_0685_),
    .D(_0682_));
 sg13g2_xor2_1 _1490_ (.B(_0685_),
    .A(\smul_up_counter.prob_counter[11] ),
    .X(_0686_));
 sg13g2_nor2_1 _1491_ (.A(net18),
    .B(_0686_),
    .Y(_0178_));
 sg13g2_buf_1 _1492_ (.A(_0450_),
    .X(_0687_));
 sg13g2_and3_1 _1493_ (.X(_0688_),
    .A(\smul_up_counter.prob_counter[11] ),
    .B(\smul_up_counter.prob_counter[10] ),
    .C(_0682_));
 sg13g2_buf_1 _1494_ (.A(_0688_),
    .X(_0689_));
 sg13g2_nand3_1 _1495_ (.B(net19),
    .C(_0689_),
    .A(net12),
    .Y(_0690_));
 sg13g2_xnor2_1 _1496_ (.Y(_0691_),
    .A(\smul_up_counter.prob_counter[12] ),
    .B(_0690_));
 sg13g2_and2_1 _1497_ (.A(net24),
    .B(_0691_),
    .X(_0179_));
 sg13g2_inv_1 _1498_ (.Y(_0692_),
    .A(\smul_up_counter.prob_counter[13] ));
 sg13g2_nand4_1 _1499_ (.B(net12),
    .C(_0678_),
    .A(\smul_up_counter.prob_counter[12] ),
    .Y(_0693_),
    .D(_0689_));
 sg13g2_xnor2_1 _1500_ (.Y(_0694_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_nor2_1 _1501_ (.A(net18),
    .B(_0694_),
    .Y(_0180_));
 sg13g2_and2_1 _1502_ (.A(\smul_up_counter.prob_counter[13] ),
    .B(\smul_up_counter.prob_counter[12] ),
    .X(_0193_));
 sg13g2_nand4_1 _1503_ (.B(net19),
    .C(_0689_),
    .A(net12),
    .Y(_0194_),
    .D(_0193_));
 sg13g2_xor2_1 _1504_ (.B(_0194_),
    .A(\smul_up_counter.prob_counter[14] ),
    .X(_0195_));
 sg13g2_nor2_1 _1505_ (.A(net18),
    .B(_0195_),
    .Y(_0181_));
 sg13g2_nand4_1 _1506_ (.B(\smul_up_counter.prob_counter[12] ),
    .C(\smul_up_counter.prob_counter[14] ),
    .A(\smul_up_counter.prob_counter[13] ),
    .Y(_0196_),
    .D(_0689_));
 sg13g2_o21ai_1 _1507_ (.B1(\smul_up_counter.prob_counter[15] ),
    .Y(_0197_),
    .A1(net8),
    .A2(_0196_));
 sg13g2_or3_1 _1508_ (.A(\smul_up_counter.prob_counter[15] ),
    .B(net8),
    .C(_0196_),
    .X(_0198_));
 sg13g2_a21oi_1 _1509_ (.A1(_0197_),
    .A2(_0198_),
    .Y(_0182_),
    .B1(net16));
 sg13g2_nand4_1 _1510_ (.B(\smul_up_counter.prob_counter[15] ),
    .C(_0689_),
    .A(\smul_up_counter.prob_counter[14] ),
    .Y(_0199_),
    .D(_0193_));
 sg13g2_o21ai_1 _1511_ (.B1(\smul_up_counter.prob_counter[16] ),
    .Y(_0200_),
    .A1(net8),
    .A2(_0199_));
 sg13g2_or3_1 _1512_ (.A(\smul_up_counter.prob_counter[16] ),
    .B(net8),
    .C(_0199_),
    .X(_0201_));
 sg13g2_a21oi_1 _1513_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0183_),
    .B1(net16));
 sg13g2_and3_1 _1514_ (.X(_0202_),
    .A(\smul_up_counter.prob_counter[0] ),
    .B(_0677_),
    .C(_0678_));
 sg13g2_xnor2_1 _1515_ (.Y(_0203_),
    .A(\smul_up_counter.prob_counter[1] ),
    .B(_0202_));
 sg13g2_nor2_1 _1516_ (.A(net18),
    .B(_0203_),
    .Y(_0184_));
 sg13g2_nand4_1 _1517_ (.B(\smul_up_counter.prob_counter[0] ),
    .C(_0672_),
    .A(\smul_up_counter.prob_counter[1] ),
    .Y(_0204_),
    .D(_0673_));
 sg13g2_nand2_1 _1518_ (.Y(_0205_),
    .A(\smul_up_counter.prob_counter[2] ),
    .B(_0204_));
 sg13g2_or2_1 _1519_ (.X(_0206_),
    .B(_0204_),
    .A(\smul_up_counter.prob_counter[2] ));
 sg13g2_a21oi_1 _1520_ (.A1(_0205_),
    .A2(_0206_),
    .Y(_0185_),
    .B1(net16));
 sg13g2_nand3_1 _1521_ (.B(\smul_up_counter.prob_counter[0] ),
    .C(\smul_up_counter.prob_counter[2] ),
    .A(\smul_up_counter.prob_counter[1] ),
    .Y(_0207_));
 sg13g2_nor2_1 _1522_ (.A(net8),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_nand2_1 _1523_ (.Y(_0209_),
    .A(\smul_up_counter.prob_counter[3] ),
    .B(_0470_));
 sg13g2_or4_1 _1524_ (.A(\smul_up_counter.prob_counter[3] ),
    .B(_0382_),
    .C(_0675_),
    .D(_0207_),
    .X(_0210_));
 sg13g2_o21ai_1 _1525_ (.B1(_0210_),
    .Y(_0186_),
    .A1(_0208_),
    .A2(_0209_));
 sg13g2_and3_1 _1526_ (.X(_0211_),
    .A(net12),
    .B(net19),
    .C(_0679_));
 sg13g2_xnor2_1 _1527_ (.Y(_0212_),
    .A(\smul_up_counter.prob_counter[4] ),
    .B(_0211_));
 sg13g2_nor2_1 _1528_ (.A(_0330_),
    .B(_0212_),
    .Y(_0187_));
 sg13g2_and4_1 _1529_ (.A(\smul_up_counter.prob_counter[4] ),
    .B(_0672_),
    .C(_0673_),
    .D(_0679_),
    .X(_0213_));
 sg13g2_xnor2_1 _1530_ (.Y(_0214_),
    .A(\smul_up_counter.prob_counter[5] ),
    .B(_0213_));
 sg13g2_nor2_1 _1531_ (.A(_0330_),
    .B(_0214_),
    .Y(_0188_));
 sg13g2_nand3_1 _1532_ (.B(\smul_up_counter.prob_counter[4] ),
    .C(_0679_),
    .A(\smul_up_counter.prob_counter[5] ),
    .Y(_0215_));
 sg13g2_o21ai_1 _1533_ (.B1(\smul_up_counter.prob_counter[6] ),
    .Y(_0216_),
    .A1(net8),
    .A2(_0215_));
 sg13g2_or3_1 _1534_ (.A(\smul_up_counter.prob_counter[6] ),
    .B(net8),
    .C(_0215_),
    .X(_0217_));
 sg13g2_a21oi_1 _1535_ (.A1(_0216_),
    .A2(_0217_),
    .Y(_0189_),
    .B1(net16));
 sg13g2_nand3_1 _1536_ (.B(net19),
    .C(_0680_),
    .A(_0677_),
    .Y(_0218_));
 sg13g2_nand2_1 _1537_ (.Y(_0219_),
    .A(\smul_up_counter.prob_counter[7] ),
    .B(_0218_));
 sg13g2_or2_1 _1538_ (.X(_0220_),
    .B(_0218_),
    .A(\smul_up_counter.prob_counter[7] ));
 sg13g2_a21oi_1 _1539_ (.A1(_0219_),
    .A2(_0220_),
    .Y(_0190_),
    .B1(net17));
 sg13g2_nand3_1 _1540_ (.B(net19),
    .C(_0681_),
    .A(net12),
    .Y(_0221_));
 sg13g2_xnor2_1 _1541_ (.Y(_0222_),
    .A(\smul_up_counter.prob_counter[8] ),
    .B(_0221_));
 sg13g2_and2_1 _1542_ (.A(net24),
    .B(_0222_),
    .X(_0191_));
 sg13g2_nand4_1 _1543_ (.B(net12),
    .C(net19),
    .A(\smul_up_counter.prob_counter[8] ),
    .Y(_0223_),
    .D(_0681_));
 sg13g2_xor2_1 _1544_ (.B(_0223_),
    .A(\smul_up_counter.prob_counter[9] ),
    .X(_0224_));
 sg13g2_nor2_1 _1545_ (.A(net18),
    .B(_0224_),
    .Y(_0192_));
 sg13g2_mux2_1 _1546_ (.A0(\add_avg[0] ),
    .A1(\add_up_counter.prob_counter[8] ),
    .S(net17),
    .X(_0060_));
 sg13g2_mux2_1 _1547_ (.A0(\add_avg[1] ),
    .A1(\add_up_counter.prob_counter[9] ),
    .S(net17),
    .X(_0061_));
 sg13g2_mux2_1 _1548_ (.A0(\add_avg[2] ),
    .A1(\add_up_counter.prob_counter[10] ),
    .S(net17),
    .X(_0062_));
 sg13g2_mux2_1 _1549_ (.A0(\add_avg[3] ),
    .A1(\add_up_counter.prob_counter[11] ),
    .S(net17),
    .X(_0063_));
 sg13g2_mux2_1 _1550_ (.A0(\add_avg[4] ),
    .A1(\add_up_counter.prob_counter[12] ),
    .S(net17),
    .X(_0064_));
 sg13g2_mux2_1 _1551_ (.A0(\add_avg[5] ),
    .A1(\add_up_counter.prob_counter[13] ),
    .S(_0383_),
    .X(_0065_));
 sg13g2_nand2_1 _1552_ (.Y(_0225_),
    .A(\add_avg[6] ),
    .B(net24));
 sg13g2_o21ai_1 _1553_ (.B1(_0225_),
    .Y(_0066_),
    .A1(_0478_),
    .A2(net24));
 sg13g2_mux2_1 _1554_ (.A0(\add_avg[7] ),
    .A1(\add_up_counter.prob_counter[15] ),
    .S(_0383_),
    .X(_0067_));
 sg13g2_nand2_1 _1555_ (.Y(_0226_),
    .A(\add_avg[8] ),
    .B(_0687_));
 sg13g2_o21ai_1 _1556_ (.B1(_0226_),
    .Y(_0068_),
    .A1(_0485_),
    .A2(_0687_));
 sg13g2_buf_1 _1557_ (.A(net35),
    .X(_0227_));
 sg13g2_mux2_1 _1558_ (.A0(\global_input.output_bitcounter_1[1] ),
    .A1(\global_input.output_bitcounter_1[0] ),
    .S(net34),
    .X(_0091_));
 sg13g2_mux2_1 _1559_ (.A0(\global_input.output_bitcounter_1[2] ),
    .A1(\global_input.output_bitcounter_1[1] ),
    .S(net34),
    .X(_0092_));
 sg13g2_mux2_1 _1560_ (.A0(\global_input.output_bitcounter_1[3] ),
    .A1(\global_input.output_bitcounter_1[2] ),
    .S(net34),
    .X(_0093_));
 sg13g2_mux2_1 _1561_ (.A0(\global_input.output_bitcounter_1[4] ),
    .A1(\global_input.output_bitcounter_1[3] ),
    .S(net34),
    .X(_0094_));
 sg13g2_mux2_1 _1562_ (.A0(\global_input.output_bitcounter_1[5] ),
    .A1(\global_input.output_bitcounter_1[4] ),
    .S(net34),
    .X(_0095_));
 sg13g2_mux2_1 _1563_ (.A0(\global_input.output_bitcounter_1[6] ),
    .A1(\global_input.output_bitcounter_1[5] ),
    .S(net34),
    .X(_0096_));
 sg13g2_mux2_1 _1564_ (.A0(\global_input.output_bitcounter_1[7] ),
    .A1(\global_input.output_bitcounter_1[6] ),
    .S(net34),
    .X(_0097_));
 sg13g2_mux2_1 _1565_ (.A0(\global_input.output_bitcounter_1[8] ),
    .A1(\global_input.output_bitcounter_1[7] ),
    .S(_0227_),
    .X(_0098_));
 sg13g2_mux2_1 _1566_ (.A0(net2),
    .A1(\global_input.output_bitcounter_1[8] ),
    .S(_0227_),
    .X(_0099_));
 sg13g2_mux2_1 _1567_ (.A0(\global_input.output_bitcounter_2[1] ),
    .A1(\global_input.output_bitcounter_2[0] ),
    .S(net34),
    .X(_0100_));
 sg13g2_mux2_1 _1568_ (.A0(\global_input.output_bitcounter_2[2] ),
    .A1(\global_input.output_bitcounter_2[1] ),
    .S(net35),
    .X(_0101_));
 sg13g2_mux2_1 _1569_ (.A0(\global_input.output_bitcounter_2[3] ),
    .A1(\global_input.output_bitcounter_2[2] ),
    .S(_0544_),
    .X(_0102_));
 sg13g2_mux2_1 _1570_ (.A0(\global_input.output_bitcounter_2[4] ),
    .A1(\global_input.output_bitcounter_2[3] ),
    .S(net35),
    .X(_0103_));
 sg13g2_mux2_1 _1571_ (.A0(\global_input.output_bitcounter_2[5] ),
    .A1(\global_input.output_bitcounter_2[4] ),
    .S(_0544_),
    .X(_0104_));
 sg13g2_mux2_1 _1572_ (.A0(\global_input.output_bitcounter_2[6] ),
    .A1(\global_input.output_bitcounter_2[5] ),
    .S(net35),
    .X(_0105_));
 sg13g2_mux2_1 _1573_ (.A0(\global_input.output_bitcounter_2[7] ),
    .A1(\global_input.output_bitcounter_2[6] ),
    .S(net35),
    .X(_0106_));
 sg13g2_mux2_1 _1574_ (.A0(\global_input.output_bitcounter_2[8] ),
    .A1(\global_input.output_bitcounter_2[7] ),
    .S(net35),
    .X(_0107_));
 sg13g2_mux2_1 _1575_ (.A0(net3),
    .A1(\global_input.output_bitcounter_2[8] ),
    .S(net35),
    .X(_0108_));
 sg13g2_mux2_1 _1576_ (.A0(\mul_avg[0] ),
    .A1(\mul_up_counter.prob_counter[8] ),
    .S(net17),
    .X(_0136_));
 sg13g2_buf_2 _1577_ (.A(net22),
    .X(_0228_));
 sg13g2_mux2_1 _1578_ (.A0(\mul_avg[1] ),
    .A1(\mul_up_counter.prob_counter[9] ),
    .S(net11),
    .X(_0137_));
 sg13g2_nand2_1 _1579_ (.Y(_0229_),
    .A(\mul_avg[2] ),
    .B(net24));
 sg13g2_o21ai_1 _1580_ (.B1(_0229_),
    .Y(_0138_),
    .A1(_0581_),
    .A2(net24));
 sg13g2_mux2_1 _1581_ (.A0(\mul_avg[3] ),
    .A1(_0567_),
    .S(net11),
    .X(_0139_));
 sg13g2_mux2_1 _1582_ (.A0(\mul_avg[4] ),
    .A1(\mul_up_counter.prob_counter[12] ),
    .S(net11),
    .X(_0140_));
 sg13g2_nand2_1 _1583_ (.Y(_0230_),
    .A(\mul_avg[5] ),
    .B(net25));
 sg13g2_o21ai_1 _1584_ (.B1(_0230_),
    .Y(_0141_),
    .A1(_0596_),
    .A2(net24));
 sg13g2_mux2_1 _1585_ (.A0(\mul_avg[6] ),
    .A1(\mul_up_counter.prob_counter[14] ),
    .S(net11),
    .X(_0142_));
 sg13g2_mux2_1 _1586_ (.A0(\mul_avg[7] ),
    .A1(\mul_up_counter.prob_counter[15] ),
    .S(_0228_),
    .X(_0143_));
 sg13g2_mux2_1 _1587_ (.A0(\mul_avg[8] ),
    .A1(\mul_up_counter.prob_counter[16] ),
    .S(_0228_),
    .X(_0144_));
 sg13g2_mux2_1 _1588_ (.A0(\smul_avg[0] ),
    .A1(\smul_up_counter.prob_counter[8] ),
    .S(net11),
    .X(_0167_));
 sg13g2_mux2_1 _1589_ (.A0(\smul_avg[1] ),
    .A1(\smul_up_counter.prob_counter[9] ),
    .S(net11),
    .X(_0168_));
 sg13g2_mux2_1 _1590_ (.A0(\smul_avg[2] ),
    .A1(\smul_up_counter.prob_counter[10] ),
    .S(net11),
    .X(_0169_));
 sg13g2_mux2_1 _1591_ (.A0(\smul_avg[3] ),
    .A1(\smul_up_counter.prob_counter[11] ),
    .S(net11),
    .X(_0170_));
 sg13g2_mux2_1 _1592_ (.A0(\smul_avg[4] ),
    .A1(\smul_up_counter.prob_counter[12] ),
    .S(net13),
    .X(_0171_));
 sg13g2_nand2_1 _1593_ (.Y(_0231_),
    .A(\smul_avg[5] ),
    .B(net25));
 sg13g2_o21ai_1 _1594_ (.B1(_0231_),
    .Y(_0172_),
    .A1(_0692_),
    .A2(net24));
 sg13g2_mux2_1 _1595_ (.A0(\smul_avg[6] ),
    .A1(\smul_up_counter.prob_counter[14] ),
    .S(net13),
    .X(_0173_));
 sg13g2_mux2_1 _1596_ (.A0(\smul_avg[7] ),
    .A1(\smul_up_counter.prob_counter[15] ),
    .S(_0579_),
    .X(_0174_));
 sg13g2_mux2_1 _1597_ (.A0(\smul_avg[8] ),
    .A1(\smul_up_counter.prob_counter[16] ),
    .S(_0579_),
    .X(_0175_));
 sg13g2_xnor2_1 _1598_ (.Y(_0050_),
    .A(\global_SN_gen.lfsr[30] ),
    .B(\global_SN_gen.lfsr[27] ));
 sg13g2_inv_1 _1599_ (.Y(_0051_),
    .A(\global_SN_gen.lfsr[9] ));
 sg13g2_inv_1 _1600_ (.Y(_0052_),
    .A(\global_SN_gen.lfsr[10] ));
 sg13g2_inv_1 _1601_ (.Y(_0053_),
    .A(\global_SN_gen.lfsr[0] ));
 sg13g2_inv_1 _1602_ (.Y(_0054_),
    .A(\global_SN_gen.lfsr[8] ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi \smul.delay_1_SN_Bit.Q$_DFF_P__95  (.L_HI(net95));
 sg13g2_buf_1 _1605_ (.A(net75),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1606_ (.A(net76),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1607_ (.A(net77),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1608_ (.A(net78),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1609_ (.A(net79),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1610_ (.A(net80),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1611_ (.A(net81),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1612_ (.A(net82),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1613_ (.A(net83),
    .X(uio_out[0]));
 sg13g2_buf_1 _1614_ (.A(net84),
    .X(uio_out[1]));
 sg13g2_buf_1 _1615_ (.A(net85),
    .X(uio_out[2]));
 sg13g2_buf_1 _1616_ (.A(net86),
    .X(uio_out[3]));
 sg13g2_buf_1 _1617_ (.A(net87),
    .X(uio_out[4]));
 sg13g2_buf_1 _1618_ (.A(net88),
    .X(uio_out[5]));
 sg13g2_buf_1 _1619_ (.A(net89),
    .X(uio_out[6]));
 sg13g2_buf_1 _1620_ (.A(net90),
    .X(uio_out[7]));
 sg13g2_buf_1 _1621_ (.A(mul_bit_out),
    .X(net4));
 sg13g2_buf_1 _1622_ (.A(add_bit_out),
    .X(net5));
 sg13g2_buf_1 _1623_ (.A(smul_bit_out),
    .X(net6));
 sg13g2_buf_1 _1624_ (.A(\add_up_counter.clk_counter[17] ),
    .X(net7));
 sg13g2_buf_1 _1625_ (.A(net91),
    .X(uo_out[4]));
 sg13g2_buf_1 _1626_ (.A(net92),
    .X(uo_out[5]));
 sg13g2_buf_1 _1627_ (.A(net93),
    .X(uo_out[6]));
 sg13g2_buf_1 _1628_ (.A(net94),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \add_output.bitseq[0]$_DFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net59),
    .D(_0018_),
    .Q_N(_0897_),
    .Q(\add_output.bitseq[0] ));
 sg13g2_dfrbp_1 \add_output.bitseq[1]$_DFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net59),
    .D(_0019_),
    .Q_N(_0896_),
    .Q(\add_output.bitseq[1] ));
 sg13g2_dfrbp_1 \add_output.bitseq[2]$_DFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net59),
    .D(_0020_),
    .Q_N(_0895_),
    .Q(\add_output.bitseq[2] ));
 sg13g2_dfrbp_1 \add_output.bitseq[3]$_DFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net60),
    .D(_0021_),
    .Q_N(_0894_),
    .Q(\add_output.bitseq[3] ));
 sg13g2_dfrbp_1 \add_output.bitseq[4]$_DFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net60),
    .D(_0022_),
    .Q_N(_0893_),
    .Q(\add_output.bitseq[4] ));
 sg13g2_dfrbp_1 \add_output.bitseq[5]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(_0023_),
    .Q_N(_0892_),
    .Q(\add_output.bitseq[5] ));
 sg13g2_dfrbp_1 \add_output.bitseq[6]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(_0024_),
    .Q_N(_0891_),
    .Q(\add_output.bitseq[6] ));
 sg13g2_dfrbp_1 \add_output.bitseq[7]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net62),
    .D(_0025_),
    .Q_N(_0890_),
    .Q(\add_output.bitseq[7] ));
 sg13g2_dfrbp_1 \add_output.bitseq[8]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(_0026_),
    .Q_N(_0889_),
    .Q(\add_output.bitseq[8] ));
 sg13g2_dfrbp_1 \add_output.counter[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net59),
    .D(_0055_),
    .Q_N(_0888_),
    .Q(\add_output.counter[0] ));
 sg13g2_dfrbp_1 \add_output.counter[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net59),
    .D(_0056_),
    .Q_N(_0887_),
    .Q(\add_output.counter[1] ));
 sg13g2_dfrbp_1 \add_output.counter[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net59),
    .D(_0057_),
    .Q_N(_0886_),
    .Q(\add_output.counter[2] ));
 sg13g2_dfrbp_1 \add_output.counter[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net59),
    .D(_0058_),
    .Q_N(_0885_),
    .Q(\add_output.counter[3] ));
 sg13g2_dfrbp_1 \add_output.output_bit$_DFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net64),
    .D(_0059_),
    .Q_N(_0884_),
    .Q(add_bit_out));
 sg13g2_dfrbp_1 \add_up_counter.average[0]$_DFFE_PP0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net58),
    .D(_0060_),
    .Q_N(_0883_),
    .Q(\add_avg[0] ));
 sg13g2_dfrbp_1 \add_up_counter.average[1]$_DFFE_PP0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net58),
    .D(_0061_),
    .Q_N(_0882_),
    .Q(\add_avg[1] ));
 sg13g2_dfrbp_1 \add_up_counter.average[2]$_DFFE_PP0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net58),
    .D(_0062_),
    .Q_N(_0881_),
    .Q(\add_avg[2] ));
 sg13g2_dfrbp_1 \add_up_counter.average[3]$_DFFE_PP0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net61),
    .D(_0063_),
    .Q_N(_0880_),
    .Q(\add_avg[3] ));
 sg13g2_dfrbp_1 \add_up_counter.average[4]$_DFFE_PP0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net61),
    .D(_0064_),
    .Q_N(_0879_),
    .Q(\add_avg[4] ));
 sg13g2_dfrbp_1 \add_up_counter.average[5]$_DFFE_PP0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net61),
    .D(_0065_),
    .Q_N(_0878_),
    .Q(\add_avg[5] ));
 sg13g2_dfrbp_1 \add_up_counter.average[6]$_DFFE_PP0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net57),
    .D(_0066_),
    .Q_N(_0877_),
    .Q(\add_avg[6] ));
 sg13g2_dfrbp_1 \add_up_counter.average[7]$_DFFE_PP0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net61),
    .D(_0067_),
    .Q_N(_0876_),
    .Q(\add_avg[7] ));
 sg13g2_dfrbp_1 \add_up_counter.average[8]$_DFFE_PP0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net57),
    .D(_0068_),
    .Q_N(_0875_),
    .Q(\add_avg[8] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net58),
    .D(_0069_),
    .Q_N(_0874_),
    .Q(\add_up_counter.prob_counter[0] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[10]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net56),
    .D(_0070_),
    .Q_N(_0873_),
    .Q(\add_up_counter.prob_counter[10] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[11]$_DFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net55),
    .D(_0071_),
    .Q_N(_0872_),
    .Q(\add_up_counter.prob_counter[11] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[12]$_DFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net61),
    .D(_0072_),
    .Q_N(_0871_),
    .Q(\add_up_counter.prob_counter[12] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[13]$_DFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net55),
    .D(_0073_),
    .Q_N(_0870_),
    .Q(\add_up_counter.prob_counter[13] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[14]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net55),
    .D(_0074_),
    .Q_N(_0869_),
    .Q(\add_up_counter.prob_counter[14] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[15]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net55),
    .D(_0075_),
    .Q_N(_0868_),
    .Q(\add_up_counter.prob_counter[15] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[16]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net55),
    .D(_0076_),
    .Q_N(_0867_),
    .Q(\add_up_counter.prob_counter[16] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net58),
    .D(_0077_),
    .Q_N(_0866_),
    .Q(\add_up_counter.prob_counter[1] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net58),
    .D(_0078_),
    .Q_N(_0865_),
    .Q(\add_up_counter.prob_counter[2] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net58),
    .D(_0079_),
    .Q_N(_0864_),
    .Q(\add_up_counter.prob_counter[3] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[4]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0080_),
    .Q_N(_0863_),
    .Q(\add_up_counter.prob_counter[4] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[5]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0081_),
    .Q_N(_0862_),
    .Q(\add_up_counter.prob_counter[5] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[6]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0082_),
    .Q_N(_0861_),
    .Q(\add_up_counter.prob_counter[6] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[7]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net56),
    .D(_0083_),
    .Q_N(_0860_),
    .Q(\add_up_counter.prob_counter[7] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[8]$_DFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net56),
    .D(_0084_),
    .Q_N(_0859_),
    .Q(\add_up_counter.prob_counter[8] ));
 sg13g2_dfrbp_1 \add_up_counter.prob_counter[9]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net58),
    .D(_0085_),
    .Q_N(_0858_),
    .Q(\add_up_counter.prob_counter[9] ));
 sg13g2_dfrbp_1 \clk_counter[0]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net53),
    .D(_0000_),
    .Q_N(_0857_),
    .Q(\add_up_counter.clk_counter[0] ));
 sg13g2_dfrbp_1 \clk_counter[10]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net48),
    .D(_0001_),
    .Q_N(_0856_),
    .Q(\add_up_counter.clk_counter[10] ));
 sg13g2_dfrbp_1 \clk_counter[11]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net48),
    .D(_0002_),
    .Q_N(_0855_),
    .Q(\add_up_counter.clk_counter[11] ));
 sg13g2_dfrbp_1 \clk_counter[12]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net48),
    .D(_0003_),
    .Q_N(_0854_),
    .Q(\add_up_counter.clk_counter[12] ));
 sg13g2_dfrbp_1 \clk_counter[13]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net49),
    .D(_0004_),
    .Q_N(_0853_),
    .Q(\add_up_counter.clk_counter[13] ));
 sg13g2_dfrbp_1 \clk_counter[14]$_DFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net49),
    .D(_0005_),
    .Q_N(_0852_),
    .Q(\add_up_counter.clk_counter[14] ));
 sg13g2_dfrbp_1 \clk_counter[15]$_DFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net49),
    .D(_0006_),
    .Q_N(_0851_),
    .Q(\add_up_counter.clk_counter[15] ));
 sg13g2_dfrbp_1 \clk_counter[16]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net49),
    .D(_0007_),
    .Q_N(_0850_),
    .Q(\add_up_counter.clk_counter[16] ));
 sg13g2_dfrbp_1 \clk_counter[17]$_DFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net52),
    .D(_0008_),
    .Q_N(_0849_),
    .Q(\add_up_counter.clk_counter[17] ));
 sg13g2_dfrbp_1 \clk_counter[1]$_DFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net52),
    .D(_0009_),
    .Q_N(_0848_),
    .Q(\add_up_counter.clk_counter[1] ));
 sg13g2_dfrbp_1 \clk_counter[2]$_DFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net52),
    .D(_0010_),
    .Q_N(_0847_),
    .Q(\add_up_counter.clk_counter[2] ));
 sg13g2_dfrbp_1 \clk_counter[3]$_DFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net51),
    .D(_0011_),
    .Q_N(_0846_),
    .Q(\add_up_counter.clk_counter[3] ));
 sg13g2_dfrbp_1 \clk_counter[4]$_DFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net51),
    .D(_0012_),
    .Q_N(_0845_),
    .Q(\add_up_counter.clk_counter[4] ));
 sg13g2_dfrbp_1 \clk_counter[5]$_DFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net51),
    .D(_0013_),
    .Q_N(_0844_),
    .Q(\add_up_counter.clk_counter[5] ));
 sg13g2_dfrbp_1 \clk_counter[6]$_DFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net51),
    .D(_0014_),
    .Q_N(_0843_),
    .Q(\add_up_counter.clk_counter[6] ));
 sg13g2_dfrbp_1 \clk_counter[7]$_DFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net49),
    .D(_0015_),
    .Q_N(_0842_),
    .Q(\add_up_counter.clk_counter[7] ));
 sg13g2_dfrbp_1 \clk_counter[8]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net49),
    .D(_0016_),
    .Q_N(_0841_),
    .Q(\add_up_counter.clk_counter[8] ));
 sg13g2_dfrbp_1 \clk_counter[9]$_DFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net48),
    .D(_0017_),
    .Q_N(_0840_),
    .Q(\add_up_counter.clk_counter[9] ));
 sg13g2_dfrbp_1 \global_input.adjustment[0]$_DFFE_PP1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net51),
    .D(_0086_),
    .Q_N(\global_input.adjustment[0] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 \global_input.adjustment[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net52),
    .D(_0087_),
    .Q_N(_0839_),
    .Q(\global_input.adjustment[1] ));
 sg13g2_dfrbp_1 \global_input.adjustment[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net52),
    .D(_0088_),
    .Q_N(_0838_),
    .Q(\global_input.adjustment[2] ));
 sg13g2_dfrbp_1 \global_input.adjustment[3]$_DFFE_PP1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net51),
    .D(_0089_),
    .Q_N(\global_input.adjustment[3] ),
    .Q(_0048_));
 sg13g2_dfrbp_1 \global_input.adjustment[4]$_DFFE_PP0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net51),
    .D(_0090_),
    .Q_N(_0837_),
    .Q(\global_input.adjustment[4] ));
 sg13g2_dfrbp_1 \global_input.loop$_DFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net52),
    .D(_0027_),
    .Q_N(_0046_),
    .Q(\global_input.loop ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[0]$_DFFE_PP0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net68),
    .D(_0091_),
    .Q_N(_0836_),
    .Q(\global_input.output_bitcounter_1[0] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[1]$_DFFE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net67),
    .D(_0092_),
    .Q_N(_0835_),
    .Q(\global_input.output_bitcounter_1[1] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[2]$_DFFE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net68),
    .D(_0093_),
    .Q_N(_0834_),
    .Q(\global_input.output_bitcounter_1[2] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[3]$_DFFE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net68),
    .D(_0094_),
    .Q_N(_0833_),
    .Q(\global_input.output_bitcounter_1[3] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[4]$_DFFE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net67),
    .D(_0095_),
    .Q_N(_0832_),
    .Q(\global_input.output_bitcounter_1[4] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[5]$_DFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net63),
    .D(_0096_),
    .Q_N(_0831_),
    .Q(\global_input.output_bitcounter_1[5] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[6]$_DFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net65),
    .D(_0097_),
    .Q_N(_0830_),
    .Q(\global_input.output_bitcounter_1[6] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[7]$_DFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0098_),
    .Q_N(_0829_),
    .Q(\global_input.output_bitcounter_1[7] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_1[8]$_DFFE_PP0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net69),
    .D(_0099_),
    .Q_N(_0828_),
    .Q(\global_input.output_bitcounter_1[8] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[0]$_DFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net71),
    .D(_0100_),
    .Q_N(_0827_),
    .Q(\global_input.output_bitcounter_2[0] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[1]$_DFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net71),
    .D(_0101_),
    .Q_N(_0826_),
    .Q(\global_input.output_bitcounter_2[1] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[2]$_DFFE_PP0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net69),
    .D(_0102_),
    .Q_N(_0825_),
    .Q(\global_input.output_bitcounter_2[2] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[3]$_DFFE_PP0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net70),
    .D(_0103_),
    .Q_N(_0824_),
    .Q(\global_input.output_bitcounter_2[3] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[4]$_DFFE_PP0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net70),
    .D(_0104_),
    .Q_N(_0823_),
    .Q(\global_input.output_bitcounter_2[4] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[5]$_DFFE_PP0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net65),
    .D(_0105_),
    .Q_N(_0822_),
    .Q(\global_input.output_bitcounter_2[5] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[6]$_DFFE_PP0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net65),
    .D(_0106_),
    .Q_N(_0821_),
    .Q(\global_input.output_bitcounter_2[6] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[7]$_DFFE_PP0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net64),
    .D(_0107_),
    .Q_N(_0820_),
    .Q(\global_input.output_bitcounter_2[7] ));
 sg13g2_dfrbp_1 \global_input.output_bitcounter_2[8]$_DFFE_PP0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net69),
    .D(_0108_),
    .Q_N(_0819_),
    .Q(\global_input.output_bitcounter_2[8] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net68),
    .D(_0109_),
    .Q_N(_0818_),
    .Q(\global_SN_gen.Input_1[0] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net68),
    .D(_0110_),
    .Q_N(_0817_),
    .Q(\global_SN_gen.Input_1[1] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net68),
    .D(_0111_),
    .Q_N(_0816_),
    .Q(\global_SN_gen.Input_1[2] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0112_),
    .Q_N(_0815_),
    .Q(\global_SN_gen.Input_1[3] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[4]$_DFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0113_),
    .Q_N(_0814_),
    .Q(\global_SN_gen.Input_1[4] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[5]$_DFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net66),
    .D(_0114_),
    .Q_N(_0813_),
    .Q(\global_SN_gen.Input_1[5] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[6]$_DFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net63),
    .D(_0115_),
    .Q_N(_0812_),
    .Q(\global_SN_gen.Input_1[6] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[7]$_DFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net63),
    .D(_0116_),
    .Q_N(_0811_),
    .Q(\global_SN_gen.Input_1[7] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_1[8]$_DFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0117_),
    .Q_N(_0810_),
    .Q(\global_SN_gen.Input_1[8] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0118_),
    .Q_N(_0809_),
    .Q(\global_SN_gen.Input_2[0] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net71),
    .D(_0119_),
    .Q_N(_0808_),
    .Q(\global_SN_gen.Input_2[1] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0120_),
    .Q_N(_0807_),
    .Q(\global_SN_gen.Input_2[2] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net70),
    .D(_0121_),
    .Q_N(_0806_),
    .Q(\global_SN_gen.Input_2[3] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[4]$_DFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net70),
    .D(_0122_),
    .Q_N(_0805_),
    .Q(\global_SN_gen.Input_2[4] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[5]$_DFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net65),
    .D(_0123_),
    .Q_N(_0804_),
    .Q(\global_SN_gen.Input_2[5] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[6]$_DFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net65),
    .D(_0124_),
    .Q_N(_0803_),
    .Q(\global_SN_gen.Input_2[6] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[7]$_DFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net64),
    .D(_0125_),
    .Q_N(_0802_),
    .Q(\global_SN_gen.Input_2[7] ));
 sg13g2_dfrbp_1 \global_input.output_bitseq_2[8]$_DFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net64),
    .D(_0126_),
    .Q_N(_0801_),
    .Q(\global_SN_gen.Input_2[8] ));
 sg13g2_dfrbp_1 \global_input.output_case[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net50),
    .D(_0127_),
    .Q_N(_0800_),
    .Q(\global_input.output_case[0] ));
 sg13g2_dfrbp_1 \global_input.output_case[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net53),
    .D(_0128_),
    .Q_N(_0799_),
    .Q(\global_input.output_case[1] ));
 sg13g2_dfrbp_1 \global_input.output_case[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net50),
    .D(_0129_),
    .Q_N(_0798_),
    .Q(\global_input.output_case[2] ));
 sg13g2_dfrbp_1 \global_input.output_case[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net53),
    .D(_0130_),
    .Q_N(_0797_),
    .Q(\global_input.output_case[3] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[0]$_DFF_PP1_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net68),
    .D(_0050_),
    .Q_N(\global_SN_gen.lfsr[0] ),
    .Q(_0899_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[10]$_DFF_PP1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net55),
    .D(_0051_),
    .Q_N(\global_SN_gen.lfsr[10] ),
    .Q(_0900_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[11]$_DFF_PP1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0052_),
    .Q_N(\global_SN_gen.lfsr[11] ),
    .Q(_0901_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[12]$_DFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(\global_SN_gen.lfsr[11] ),
    .Q_N(_0796_),
    .Q(\global_SN_gen.lfsr[12] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[13]$_DFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net70),
    .D(\global_SN_gen.lfsr[12] ),
    .Q_N(_0795_),
    .Q(\global_SN_gen.lfsr[13] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[14]$_DFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net70),
    .D(\global_SN_gen.lfsr[13] ),
    .Q_N(_0794_),
    .Q(\global_SN_gen.lfsr[14] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[15]$_DFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net70),
    .D(\global_SN_gen.lfsr[14] ),
    .Q_N(_0793_),
    .Q(\global_SN_gen.lfsr[15] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[16]$_DFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net64),
    .D(\global_SN_gen.lfsr[15] ),
    .Q_N(_0792_),
    .Q(\global_SN_gen.lfsr[16] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[17]$_DFF_PP1_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net70),
    .D(_0792_),
    .Q_N(\global_SN_gen.lfsr[17] ),
    .Q(_0902_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[18]$_DFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net65),
    .D(\global_SN_gen.lfsr[17] ),
    .Q_N(_0791_),
    .Q(\global_SN_gen.lfsr[18] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[19]$_DFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net64),
    .D(\global_SN_gen.lfsr[18] ),
    .Q_N(_0790_),
    .Q(\global_SN_gen.lfsr[19] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[1]$_DFF_PP1_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net67),
    .D(_0053_),
    .Q_N(\global_SN_gen.lfsr[1] ),
    .Q(_0903_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[20]$_DFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net64),
    .D(\global_SN_gen.lfsr[19] ),
    .Q_N(_0789_),
    .Q(\global_SN_gen.lfsr[20] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[21]$_DFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net55),
    .D(\global_SN_gen.lfsr[20] ),
    .Q_N(_0788_),
    .Q(\global_SN_gen.lfsr[21] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[22]$_DFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net57),
    .D(\global_SN_gen.lfsr[21] ),
    .Q_N(_0787_),
    .Q(\global_SN_gen.lfsr[22] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[23]$_DFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net55),
    .D(\global_SN_gen.lfsr[22] ),
    .Q_N(_0786_),
    .Q(\global_SN_gen.lfsr[23] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[24]$_DFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net61),
    .D(\global_SN_gen.lfsr[23] ),
    .Q_N(_0785_),
    .Q(\global_SN_gen.lfsr[24] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[25]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net61),
    .D(\global_SN_gen.lfsr[24] ),
    .Q_N(_0784_),
    .Q(\global_SN_gen.lfsr[25] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[26]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(\global_SN_gen.lfsr[25] ),
    .Q_N(_0783_),
    .Q(\global_SN_gen.lfsr[26] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[27]$_DFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net60),
    .D(\global_SN_gen.lfsr[26] ),
    .Q_N(_0782_),
    .Q(\global_SN_gen.lfsr[27] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[28]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net60),
    .D(\global_SN_gen.lfsr[27] ),
    .Q_N(_0781_),
    .Q(\global_SN_gen.lfsr[28] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[29]$_DFF_PP0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net62),
    .D(\global_SN_gen.lfsr[28] ),
    .Q_N(_0780_),
    .Q(\global_SN_gen.lfsr[29] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[2]$_DFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net67),
    .D(\global_SN_gen.lfsr[1] ),
    .Q_N(_0779_),
    .Q(\global_SN_gen.lfsr[2] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[30]$_DFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net62),
    .D(\global_SN_gen.lfsr[29] ),
    .Q_N(_0778_),
    .Q(\global_SN_gen.lfsr[30] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[3]$_DFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net63),
    .D(\global_SN_gen.lfsr[2] ),
    .Q_N(_0777_),
    .Q(\global_SN_gen.lfsr[3] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[4]$_DFF_PP1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0777_),
    .Q_N(\global_SN_gen.lfsr[4] ),
    .Q(_0904_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[5]$_DFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net63),
    .D(\global_SN_gen.lfsr[4] ),
    .Q_N(_0776_),
    .Q(\global_SN_gen.lfsr[5] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[6]$_DFF_PP1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net63),
    .D(_0776_),
    .Q_N(\global_SN_gen.lfsr[6] ),
    .Q(_0905_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[7]$_DFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net63),
    .D(\global_SN_gen.lfsr[6] ),
    .Q_N(_0775_),
    .Q(\global_SN_gen.lfsr[7] ));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[8]$_DFF_PP1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net63),
    .D(_0775_),
    .Q_N(\global_SN_gen.lfsr[8] ),
    .Q(_0906_));
 sg13g2_dfrbp_1 \global_lsfr.lfsr[9]$_DFF_PP1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net66),
    .D(_0054_),
    .Q_N(\global_SN_gen.lfsr[9] ),
    .Q(_0907_));
 sg13g2_dfrbp_1 \mul_output.bitseq[0]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net50),
    .D(_0028_),
    .Q_N(_0774_),
    .Q(\mul_output.bitseq[0] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[1]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net50),
    .D(_0029_),
    .Q_N(_0773_),
    .Q(\mul_output.bitseq[1] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[2]$_DFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net47),
    .D(_0030_),
    .Q_N(_0772_),
    .Q(\mul_output.bitseq[2] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[3]$_DFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net49),
    .D(_0031_),
    .Q_N(_0771_),
    .Q(\mul_output.bitseq[3] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[4]$_DFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net54),
    .D(_0032_),
    .Q_N(_0770_),
    .Q(\mul_output.bitseq[4] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[5]$_DFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net47),
    .D(_0033_),
    .Q_N(_0769_),
    .Q(\mul_output.bitseq[5] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[6]$_DFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0034_),
    .Q_N(_0768_),
    .Q(\mul_output.bitseq[6] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[7]$_DFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0035_),
    .Q_N(_0767_),
    .Q(\mul_output.bitseq[7] ));
 sg13g2_dfrbp_1 \mul_output.bitseq[8]$_DFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net46),
    .D(_0036_),
    .Q_N(_0766_),
    .Q(\mul_output.bitseq[8] ));
 sg13g2_dfrbp_1 \mul_output.counter[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net48),
    .D(_0131_),
    .Q_N(_0765_),
    .Q(\mul_output.counter[0] ));
 sg13g2_dfrbp_1 \mul_output.counter[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net48),
    .D(_0132_),
    .Q_N(_0764_),
    .Q(\mul_output.counter[1] ));
 sg13g2_dfrbp_1 \mul_output.counter[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net48),
    .D(_0133_),
    .Q_N(_0763_),
    .Q(\mul_output.counter[2] ));
 sg13g2_dfrbp_1 \mul_output.counter[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net48),
    .D(_0134_),
    .Q_N(_0762_),
    .Q(\mul_output.counter[3] ));
 sg13g2_dfrbp_1 \mul_output.output_bit$_DFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net64),
    .D(_0135_),
    .Q_N(_0761_),
    .Q(mul_bit_out));
 sg13g2_dfrbp_1 \mul_up_counter.average[0]$_DFFE_PP0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net50),
    .D(_0136_),
    .Q_N(_0760_),
    .Q(\mul_avg[0] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[1]$_DFFE_PP0N_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net50),
    .D(_0137_),
    .Q_N(_0759_),
    .Q(\mul_avg[1] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[2]$_DFFE_PP0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net50),
    .D(_0138_),
    .Q_N(_0758_),
    .Q(\mul_avg[2] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[3]$_DFFE_PP0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net47),
    .D(_0139_),
    .Q_N(_0757_),
    .Q(\mul_avg[3] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[4]$_DFFE_PP0N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net47),
    .D(_0140_),
    .Q_N(_0756_),
    .Q(\mul_avg[4] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[5]$_DFFE_PP0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net47),
    .D(_0141_),
    .Q_N(_0755_),
    .Q(\mul_avg[5] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[6]$_DFFE_PP0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0142_),
    .Q_N(_0754_),
    .Q(\mul_avg[6] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[7]$_DFFE_PP0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0143_),
    .Q_N(_0753_),
    .Q(\mul_avg[7] ));
 sg13g2_dfrbp_1 \mul_up_counter.average[8]$_DFFE_PP0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0144_),
    .Q_N(_0752_),
    .Q(\mul_avg[8] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net38),
    .D(_0145_),
    .Q_N(_0751_),
    .Q(\mul_up_counter.prob_counter[0] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[10]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net50),
    .D(_0146_),
    .Q_N(_0750_),
    .Q(\mul_up_counter.prob_counter[10] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[11]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net41),
    .D(_0147_),
    .Q_N(_0749_),
    .Q(\mul_up_counter.prob_counter[11] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[12]$_DFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net47),
    .D(_0148_),
    .Q_N(_0748_),
    .Q(\mul_up_counter.prob_counter[12] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[13]$_DFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net47),
    .D(_0149_),
    .Q_N(_0747_),
    .Q(\mul_up_counter.prob_counter[13] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[14]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net40),
    .D(_0150_),
    .Q_N(_0746_),
    .Q(\mul_up_counter.prob_counter[14] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[15]$_DFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0151_),
    .Q_N(_0745_),
    .Q(\mul_up_counter.prob_counter[15] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[16]$_DFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net46),
    .D(_0152_),
    .Q_N(_0744_),
    .Q(\mul_up_counter.prob_counter[16] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net38),
    .D(_0153_),
    .Q_N(_0743_),
    .Q(\mul_up_counter.prob_counter[1] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net40),
    .D(_0154_),
    .Q_N(_0742_),
    .Q(\mul_up_counter.prob_counter[2] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net40),
    .D(_0155_),
    .Q_N(_0741_),
    .Q(\mul_up_counter.prob_counter[3] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[4]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net40),
    .D(_0156_),
    .Q_N(_0740_),
    .Q(\mul_up_counter.prob_counter[4] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[5]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net40),
    .D(_0157_),
    .Q_N(_0739_),
    .Q(\mul_up_counter.prob_counter[5] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[6]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net40),
    .D(_0158_),
    .Q_N(_0738_),
    .Q(\mul_up_counter.prob_counter[6] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[7]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net40),
    .D(_0159_),
    .Q_N(_0737_),
    .Q(\mul_up_counter.prob_counter[7] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[8]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net44),
    .D(_0160_),
    .Q_N(_0736_),
    .Q(\mul_up_counter.prob_counter[8] ));
 sg13g2_dfrbp_1 \mul_up_counter.prob_counter[9]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net44),
    .D(_0161_),
    .Q_N(_0898_),
    .Q(\mul_up_counter.prob_counter[9] ));
 sg13g2_dfrbp_1 \smul.delay_1_SN_Bit.Q$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net95),
    .D(SN_Bit_1),
    .Q_N(_0735_),
    .Q(\smul.SN_Bit_Q ));
 sg13g2_dfrbp_1 \smul_output.bitseq[0]$_DFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net39),
    .D(_0037_),
    .Q_N(_0734_),
    .Q(\smul_output.bitseq[0] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[1]$_DFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net39),
    .D(_0038_),
    .Q_N(_0733_),
    .Q(\smul_output.bitseq[1] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[2]$_DFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net39),
    .D(_0039_),
    .Q_N(_0732_),
    .Q(\smul_output.bitseq[2] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[3]$_DFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net39),
    .D(_0040_),
    .Q_N(_0731_),
    .Q(\smul_output.bitseq[3] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[4]$_DFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net43),
    .D(_0041_),
    .Q_N(_0730_),
    .Q(\smul_output.bitseq[4] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[5]$_DFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net42),
    .D(_0042_),
    .Q_N(_0729_),
    .Q(\smul_output.bitseq[5] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[6]$_DFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net42),
    .D(_0043_),
    .Q_N(_0728_),
    .Q(\smul_output.bitseq[6] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[7]$_DFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net43),
    .D(_0044_),
    .Q_N(_0727_),
    .Q(\smul_output.bitseq[7] ));
 sg13g2_dfrbp_1 \smul_output.bitseq[8]$_DFF_PP0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net43),
    .D(_0045_),
    .Q_N(_0726_),
    .Q(\smul_output.bitseq[8] ));
 sg13g2_dfrbp_1 \smul_output.counter[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0162_),
    .Q_N(_0725_),
    .Q(\smul_output.counter[0] ));
 sg13g2_dfrbp_1 \smul_output.counter[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net56),
    .D(_0163_),
    .Q_N(_0724_),
    .Q(\smul_output.counter[1] ));
 sg13g2_dfrbp_1 \smul_output.counter[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net42),
    .D(_0164_),
    .Q_N(_0723_),
    .Q(\smul_output.counter[2] ));
 sg13g2_dfrbp_1 \smul_output.counter[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net42),
    .D(_0165_),
    .Q_N(_0722_),
    .Q(\smul_output.counter[3] ));
 sg13g2_dfrbp_1 \smul_output.output_bit$_DFFE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net51),
    .D(_0166_),
    .Q_N(_0721_),
    .Q(smul_bit_out));
 sg13g2_dfrbp_1 \smul_up_counter.average[0]$_DFFE_PP0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net38),
    .D(_0167_),
    .Q_N(_0720_),
    .Q(\smul_avg[0] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[1]$_DFFE_PP0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net39),
    .D(_0168_),
    .Q_N(_0719_),
    .Q(\smul_avg[1] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[2]$_DFFE_PP0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net38),
    .D(_0169_),
    .Q_N(_0718_),
    .Q(\smul_avg[2] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[3]$_DFFE_PP0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net38),
    .D(_0170_),
    .Q_N(_0717_),
    .Q(\smul_avg[3] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[4]$_DFFE_PP0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net38),
    .D(_0171_),
    .Q_N(_0716_),
    .Q(\smul_avg[4] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[5]$_DFFE_PP0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net43),
    .D(_0172_),
    .Q_N(_0715_),
    .Q(\smul_avg[5] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[6]$_DFFE_PP0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net43),
    .D(_0173_),
    .Q_N(_0714_),
    .Q(\smul_avg[6] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[7]$_DFFE_PP0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net42),
    .D(_0174_),
    .Q_N(_0713_),
    .Q(\smul_avg[7] ));
 sg13g2_dfrbp_1 \smul_up_counter.average[8]$_DFFE_PP0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net42),
    .D(_0175_),
    .Q_N(_0712_),
    .Q(\smul_avg[8] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net45),
    .D(_0176_),
    .Q_N(_0711_),
    .Q(\smul_up_counter.prob_counter[0] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[10]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net38),
    .D(_0177_),
    .Q_N(_0710_),
    .Q(\smul_up_counter.prob_counter[10] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[11]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net38),
    .D(_0178_),
    .Q_N(_0709_),
    .Q(\smul_up_counter.prob_counter[11] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[12]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net44),
    .D(_0179_),
    .Q_N(_0708_),
    .Q(\smul_up_counter.prob_counter[12] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[13]$_DFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net43),
    .D(_0180_),
    .Q_N(_0707_),
    .Q(\smul_up_counter.prob_counter[13] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[14]$_DFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net43),
    .D(_0181_),
    .Q_N(_0706_),
    .Q(\smul_up_counter.prob_counter[14] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[15]$_DFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net42),
    .D(_0182_),
    .Q_N(_0705_),
    .Q(\smul_up_counter.prob_counter[15] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[16]$_DFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net42),
    .D(_0183_),
    .Q_N(_0704_),
    .Q(\smul_up_counter.prob_counter[16] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net45),
    .D(_0184_),
    .Q_N(_0703_),
    .Q(\smul_up_counter.prob_counter[1] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[2]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net45),
    .D(_0185_),
    .Q_N(_0702_),
    .Q(\smul_up_counter.prob_counter[2] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[3]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net44),
    .D(_0186_),
    .Q_N(_0701_),
    .Q(\smul_up_counter.prob_counter[3] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[4]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net44),
    .D(_0187_),
    .Q_N(_0700_),
    .Q(\smul_up_counter.prob_counter[4] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[5]$_DFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net44),
    .D(_0188_),
    .Q_N(_0699_),
    .Q(\smul_up_counter.prob_counter[5] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[6]$_DFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net44),
    .D(_0189_),
    .Q_N(_0698_),
    .Q(\smul_up_counter.prob_counter[6] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[7]$_DFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net44),
    .D(_0190_),
    .Q_N(_0697_),
    .Q(\smul_up_counter.prob_counter[7] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[8]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net40),
    .D(_0191_),
    .Q_N(_0696_),
    .Q(\smul_up_counter.prob_counter[8] ));
 sg13g2_dfrbp_1 \smul_up_counter.prob_counter[9]$_DFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net41),
    .D(_0192_),
    .Q_N(_0695_),
    .Q(\smul_up_counter.prob_counter[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[0]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[1]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[2]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[3]));
 sg13g2_buf_2 fanout8 (.A(_0675_),
    .X(net8));
 sg13g2_buf_2 fanout9 (.A(_0577_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_0575_),
    .X(net10));
 sg13g2_buf_4 fanout11 (.X(net11),
    .A(_0228_));
 sg13g2_buf_2 fanout12 (.A(_0677_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0579_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0574_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0468_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0464_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0383_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0330_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0678_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0571_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0462_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0382_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0329_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0687_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0470_),
    .X(net25));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(_0392_));
 sg13g2_buf_2 fanout27 (.A(_0391_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0360_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0298_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0269_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0356_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0293_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0265_),
    .X(net33));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(_0227_));
 sg13g2_buf_2 fanout35 (.A(_0544_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0522_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0521_),
    .X(net37));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(net41));
 sg13g2_buf_2 fanout39 (.A(net41),
    .X(net39));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(net41));
 sg13g2_buf_2 fanout41 (.A(net74),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net43));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(net45));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(net45));
 sg13g2_buf_2 fanout45 (.A(net74),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(net47));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(net54));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(net49));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(net54));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(net53));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(net53));
 sg13g2_buf_2 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(net54),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net74),
    .X(net54));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(net57));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(net73));
 sg13g2_buf_2 fanout57 (.A(net73),
    .X(net57));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(net62));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(net62));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(net61));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net62));
 sg13g2_buf_2 fanout62 (.A(net73),
    .X(net62));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net66));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(net66));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(net73),
    .X(net66));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(net72));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(net72));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(net71));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(net72));
 sg13g2_buf_2 fanout71 (.A(net72),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(_0049_),
    .X(net74));
 sg13g2_tielo _1605__75 (.L_LO(net75));
 sg13g2_tielo _1606__76 (.L_LO(net76));
 sg13g2_tielo _1607__77 (.L_LO(net77));
 sg13g2_tielo _1608__78 (.L_LO(net78));
 sg13g2_tielo _1609__79 (.L_LO(net79));
 sg13g2_tielo _1610__80 (.L_LO(net80));
 sg13g2_tielo _1611__81 (.L_LO(net81));
 sg13g2_tielo _1612__82 (.L_LO(net82));
 sg13g2_tielo _1613__83 (.L_LO(net83));
 sg13g2_tielo _1614__84 (.L_LO(net84));
 sg13g2_tielo _1615__85 (.L_LO(net85));
 sg13g2_tielo _1616__86 (.L_LO(net86));
 sg13g2_tielo _1617__87 (.L_LO(net87));
 sg13g2_tielo _1618__88 (.L_LO(net88));
 sg13g2_tielo _1619__89 (.L_LO(net89));
 sg13g2_tielo _1620__90 (.L_LO(net90));
 sg13g2_tielo _1625__91 (.L_LO(net91));
 sg13g2_tielo _1626__92 (.L_LO(net92));
 sg13g2_tielo _1627__93 (.L_LO(net93));
 sg13g2_tielo _1628__94 (.L_LO(net94));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0166_));
 sg13g2_antennanp ANTENNA_2 (.A(_0166_));
 sg13g2_antennanp ANTENNA_3 (.A(_0166_));
 sg13g2_antennanp ANTENNA_4 (.A(_0166_));
 sg13g2_antennanp ANTENNA_5 (.A(_0166_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_4 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_4 FILLER_0_185 ();
 sg13g2_fill_2 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_4 FILLER_0_297 ();
 sg13g2_fill_2 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_fill_1 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_decap_8 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_100 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_fill_2 FILLER_1_189 ();
 sg13g2_fill_1 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_decap_8 FILLER_1_237 ();
 sg13g2_decap_8 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_decap_4 FILLER_1_265 ();
 sg13g2_fill_2 FILLER_1_269 ();
 sg13g2_decap_4 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_4 FILLER_2_70 ();
 sg13g2_fill_2 FILLER_2_90 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_decap_4 FILLER_2_124 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_fill_2 FILLER_2_187 ();
 sg13g2_fill_1 FILLER_2_189 ();
 sg13g2_fill_2 FILLER_2_208 ();
 sg13g2_fill_1 FILLER_2_210 ();
 sg13g2_fill_2 FILLER_2_219 ();
 sg13g2_fill_1 FILLER_2_221 ();
 sg13g2_decap_4 FILLER_2_248 ();
 sg13g2_fill_1 FILLER_2_252 ();
 sg13g2_fill_2 FILLER_2_279 ();
 sg13g2_fill_2 FILLER_2_317 ();
 sg13g2_fill_1 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_4 FILLER_3_63 ();
 sg13g2_fill_2 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_180 ();
 sg13g2_fill_1 FILLER_3_187 ();
 sg13g2_fill_2 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_3_201 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_4 FILLER_3_256 ();
 sg13g2_fill_1 FILLER_3_260 ();
 sg13g2_fill_2 FILLER_3_296 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_4 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_68 ();
 sg13g2_fill_2 FILLER_4_75 ();
 sg13g2_fill_1 FILLER_4_94 ();
 sg13g2_decap_4 FILLER_4_100 ();
 sg13g2_fill_2 FILLER_4_108 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_fill_2 FILLER_4_123 ();
 sg13g2_fill_1 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_131 ();
 sg13g2_fill_1 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_148 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_fill_1 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_fill_2 FILLER_4_199 ();
 sg13g2_fill_1 FILLER_4_201 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_4 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_fill_2 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_4 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_4 FILLER_4_370 ();
 sg13g2_fill_2 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_414 ();
 sg13g2_decap_8 FILLER_4_421 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_75 ();
 sg13g2_decap_4 FILLER_5_82 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_146 ();
 sg13g2_fill_2 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_164 ();
 sg13g2_decap_8 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_206 ();
 sg13g2_decap_8 FILLER_5_213 ();
 sg13g2_decap_8 FILLER_5_220 ();
 sg13g2_decap_8 FILLER_5_227 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_fill_2 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_fill_2 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_4 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_4 FILLER_5_369 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_4 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_32 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_decap_4 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_128 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_8 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_215 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_decap_4 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_fill_2 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_fill_1 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_fill_1 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_4 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_46 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_146 ();
 sg13g2_fill_2 FILLER_7_153 ();
 sg13g2_fill_2 FILLER_7_169 ();
 sg13g2_fill_1 FILLER_7_171 ();
 sg13g2_decap_4 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_228 ();
 sg13g2_fill_2 FILLER_7_235 ();
 sg13g2_fill_1 FILLER_7_237 ();
 sg13g2_fill_1 FILLER_7_264 ();
 sg13g2_fill_2 FILLER_7_272 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_1 FILLER_7_282 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_4 FILLER_7_380 ();
 sg13g2_decap_4 FILLER_7_397 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_decap_8 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_120 ();
 sg13g2_fill_2 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_fill_1 FILLER_8_251 ();
 sg13g2_fill_1 FILLER_8_265 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_fill_2 FILLER_8_316 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_40 ();
 sg13g2_decap_8 FILLER_9_47 ();
 sg13g2_decap_8 FILLER_9_54 ();
 sg13g2_decap_8 FILLER_9_61 ();
 sg13g2_decap_8 FILLER_9_68 ();
 sg13g2_fill_2 FILLER_9_75 ();
 sg13g2_decap_4 FILLER_9_84 ();
 sg13g2_fill_1 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_106 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_fill_2 FILLER_9_130 ();
 sg13g2_fill_1 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_171 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_191 ();
 sg13g2_decap_4 FILLER_9_198 ();
 sg13g2_fill_2 FILLER_9_202 ();
 sg13g2_fill_2 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_258 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_fill_2 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_4 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_1 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_4 FILLER_9_370 ();
 sg13g2_fill_1 FILLER_9_384 ();
 sg13g2_fill_2 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_16 ();
 sg13g2_decap_4 FILLER_10_64 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_4 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_fill_2 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_170 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_fill_2 FILLER_10_267 ();
 sg13g2_decap_4 FILLER_10_274 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_fill_1 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_fill_1 FILLER_10_378 ();
 sg13g2_fill_1 FILLER_10_388 ();
 sg13g2_fill_2 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_decap_8 FILLER_11_59 ();
 sg13g2_decap_8 FILLER_11_66 ();
 sg13g2_decap_4 FILLER_11_73 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_decap_4 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_135 ();
 sg13g2_decap_8 FILLER_11_142 ();
 sg13g2_decap_8 FILLER_11_149 ();
 sg13g2_decap_8 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_decap_8 FILLER_11_199 ();
 sg13g2_decap_8 FILLER_11_206 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_fill_2 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_4 FILLER_11_366 ();
 sg13g2_decap_4 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_45 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_decap_8 FILLER_12_61 ();
 sg13g2_decap_8 FILLER_12_68 ();
 sg13g2_decap_4 FILLER_12_75 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_151 ();
 sg13g2_fill_1 FILLER_12_153 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_4 FILLER_12_175 ();
 sg13g2_decap_4 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_201 ();
 sg13g2_decap_8 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_decap_4 FILLER_12_229 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_fill_2 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_16 ();
 sg13g2_decap_8 FILLER_13_59 ();
 sg13g2_decap_4 FILLER_13_66 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_143 ();
 sg13g2_fill_1 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_decap_4 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_239 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_4 FILLER_13_308 ();
 sg13g2_fill_2 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_4 FILLER_13_357 ();
 sg13g2_fill_1 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_decap_4 FILLER_13_372 ();
 sg13g2_fill_2 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_13_409 ();
 sg13g2_decap_8 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_58 ();
 sg13g2_decap_4 FILLER_14_65 ();
 sg13g2_fill_2 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_76 ();
 sg13g2_fill_2 FILLER_14_80 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_4 FILLER_14_130 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_393 ();
 sg13g2_fill_1 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_11 ();
 sg13g2_fill_1 FILLER_15_54 ();
 sg13g2_fill_1 FILLER_15_59 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_2 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_2 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_50 ();
 sg13g2_decap_8 FILLER_16_57 ();
 sg13g2_decap_8 FILLER_16_64 ();
 sg13g2_decap_4 FILLER_16_71 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_fill_2 FILLER_16_92 ();
 sg13g2_fill_2 FILLER_16_101 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_fill_2 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_4 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_18 ();
 sg13g2_fill_2 FILLER_17_43 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_4 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_71 ();
 sg13g2_decap_4 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_89 ();
 sg13g2_decap_4 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_114 ();
 sg13g2_decap_4 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_141 ();
 sg13g2_decap_8 FILLER_17_148 ();
 sg13g2_decap_8 FILLER_17_155 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_2 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_4 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_4 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_395 ();
 sg13g2_fill_1 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_424 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_decap_8 FILLER_18_155 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_4 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_decap_4 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_decap_4 FILLER_18_323 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_27 ();
 sg13g2_fill_1 FILLER_19_34 ();
 sg13g2_fill_1 FILLER_19_40 ();
 sg13g2_fill_1 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_2 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_178 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_decap_8 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_decap_4 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_decap_4 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_4 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_113 ();
 sg13g2_decap_4 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_decap_4 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_142 ();
 sg13g2_decap_8 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_4 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_fill_1 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_decap_4 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_4 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_45 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_232 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_290 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_412 ();
 sg13g2_decap_8 FILLER_22_419 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_45 ();
 sg13g2_decap_4 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_106 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_decap_4 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_decap_8 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_211 ();
 sg13g2_decap_4 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_258 ();
 sg13g2_decap_4 FILLER_23_265 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_4 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_330 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_157 ();
 sg13g2_decap_4 FILLER_24_164 ();
 sg13g2_fill_1 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_decap_4 FILLER_24_386 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_4 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_38 ();
 sg13g2_decap_8 FILLER_25_65 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_239 ();
 sg13g2_decap_4 FILLER_25_246 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_23 ();
 sg13g2_decap_4 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_58 ();
 sg13g2_decap_4 FILLER_26_66 ();
 sg13g2_decap_8 FILLER_26_75 ();
 sg13g2_fill_2 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_104 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_150 ();
 sg13g2_decap_4 FILLER_26_157 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_decap_4 FILLER_26_255 ();
 sg13g2_decap_4 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_311 ();
 sg13g2_decap_4 FILLER_26_318 ();
 sg13g2_decap_4 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_4 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_79 ();
 sg13g2_fill_2 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_143 ();
 sg13g2_decap_4 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_418 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_decap_4 FILLER_28_37 ();
 sg13g2_decap_4 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_decap_4 FILLER_28_142 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_decap_4 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_250 ();
 sg13g2_decap_4 FILLER_28_257 ();
 sg13g2_fill_2 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_4 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_fill_1 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_415 ();
 sg13g2_decap_8 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_33 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_54 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_fill_1 FILLER_29_69 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_4 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_fill_2 FILLER_29_381 ();
 sg13g2_fill_1 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_65 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_decap_8 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_decap_8 FILLER_30_93 ();
 sg13g2_decap_8 FILLER_30_100 ();
 sg13g2_decap_8 FILLER_30_107 ();
 sg13g2_decap_8 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_decap_4 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_9 ();
 sg13g2_decap_8 FILLER_31_66 ();
 sg13g2_decap_4 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_decap_8 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_4 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_2 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_61 ();
 sg13g2_decap_8 FILLER_32_68 ();
 sg13g2_decap_4 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_113 ();
 sg13g2_fill_1 FILLER_32_120 ();
 sg13g2_decap_8 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_206 ();
 sg13g2_decap_4 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_decap_4 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_286 ();
 sg13g2_decap_4 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_4 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_349 ();
 sg13g2_decap_4 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_decap_4 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_36 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_55 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_decap_4 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_decap_4 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_decap_4 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_52 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_decap_8 FILLER_34_106 ();
 sg13g2_decap_8 FILLER_34_113 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_269 ();
 sg13g2_decap_4 FILLER_34_276 ();
 sg13g2_fill_2 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_2 FILLER_35_104 ();
 sg13g2_fill_1 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_4 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_decap_4 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_decap_4 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_fill_1 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_416 ();
 sg13g2_decap_8 FILLER_35_423 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_16 ();
 sg13g2_decap_8 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_decap_8 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_decap_4 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_37_34 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_2 FILLER_37_58 ();
 sg13g2_decap_8 FILLER_37_68 ();
 sg13g2_fill_2 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_decap_4 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_decap_4 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_decap_4 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_267 ();
 sg13g2_decap_4 FILLER_37_274 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_4 FILLER_37_319 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_23 ();
 sg13g2_decap_8 FILLER_38_32 ();
 sg13g2_decap_4 FILLER_38_39 ();
 sg13g2_fill_2 FILLER_38_43 ();
 sg13g2_decap_8 FILLER_38_51 ();
 sg13g2_decap_8 FILLER_38_58 ();
 sg13g2_decap_8 FILLER_38_65 ();
 sg13g2_decap_8 FILLER_38_72 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_decap_4 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_4 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_379 ();
 sg13g2_decap_4 FILLER_38_388 ();
 sg13g2_fill_1 FILLER_38_392 ();
 sg13g2_fill_2 FILLER_38_415 ();
 sg13g2_fill_1 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
